//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 1 0 1 1 0 0 1 1 1 0 0 1 0 1 0 0 0 0 0 0 1 1 0 1 1 1 0 0 1 0 0 1 1 0 1 1 0 0 1 1 1 1 1 0 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:42 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  XNOR2_X1  g0001(.A(new_n201), .B(KEYINPUT64), .ZN(new_n202));
  INV_X1    g0002(.A(G77), .ZN(new_n203));
  AND2_X1   g0003(.A1(new_n202), .A2(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NOR2_X1   g0005(.A1(G58), .A2(G68), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  OR2_X1    g0007(.A1(new_n207), .A2(KEYINPUT65), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(KEYINPUT65), .ZN(new_n209));
  NAND3_X1  g0009(.A1(new_n208), .A2(G50), .A3(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  NOR3_X1   g0012(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G20), .ZN(new_n214));
  XOR2_X1   g0014(.A(KEYINPUT66), .B(G238), .Z(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  OR2_X1    g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G107), .A2(G264), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G58), .A2(G232), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G77), .A2(G244), .ZN(new_n220));
  NAND4_X1  g0020(.A1(new_n217), .A2(new_n218), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n221), .B1(G50), .B2(G226), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G116), .A2(G270), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G97), .A2(G257), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  AND2_X1   g0025(.A1(G87), .A2(G250), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n214), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT1), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n214), .A2(G13), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n229), .B(G250), .C1(G257), .C2(G264), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(KEYINPUT0), .ZN(new_n231));
  OR2_X1    g0031(.A1(new_n230), .A2(KEYINPUT0), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n213), .B(new_n228), .C1(new_n231), .C2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G250), .B(G257), .Z(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G68), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(KEYINPUT77), .ZN(new_n249));
  XOR2_X1   g0049(.A(KEYINPUT8), .B(G58), .Z(new_n250));
  INV_X1    g0050(.A(G1), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(G13), .A3(G20), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  AND2_X1   g0055(.A1(new_n255), .A2(new_n212), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n251), .A2(G20), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n254), .B1(new_n258), .B2(new_n250), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n262));
  OR2_X1    g0062(.A1(G223), .A2(G1698), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT3), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G33), .ZN(new_n265));
  INV_X1    g0065(.A(G226), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G1698), .ZN(new_n267));
  NAND4_X1  g0067(.A1(new_n262), .A2(new_n263), .A3(new_n265), .A4(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G87), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G41), .ZN(new_n271));
  OAI211_X1 g0071(.A(G1), .B(G13), .C1(new_n261), .C2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n251), .B1(G41), .B2(G45), .ZN(new_n275));
  AND3_X1   g0075(.A1(new_n272), .A2(G232), .A3(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G190), .ZN(new_n278));
  INV_X1    g0078(.A(G274), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n274), .A2(new_n277), .A3(new_n278), .A4(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n272), .B1(new_n268), .B2(new_n269), .ZN(new_n283));
  NOR3_X1   g0083(.A1(new_n283), .A2(new_n280), .A3(new_n276), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n282), .B1(new_n284), .B2(G200), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT74), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n286), .B1(new_n264), .B2(G33), .ZN(new_n287));
  OAI21_X1  g0087(.A(KEYINPUT75), .B1(new_n261), .B2(KEYINPUT3), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT75), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n289), .A2(new_n264), .A3(G33), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n261), .A2(KEYINPUT74), .A3(KEYINPUT3), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n287), .A2(new_n288), .A3(new_n290), .A4(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT7), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n293), .A2(G20), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n264), .A2(G33), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n211), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(new_n293), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n295), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G68), .ZN(new_n301));
  INV_X1    g0101(.A(G58), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n302), .A2(new_n216), .ZN(new_n303));
  OAI21_X1  g0103(.A(G20), .B1(new_n303), .B2(new_n206), .ZN(new_n304));
  NOR2_X1   g0104(.A1(G20), .A2(G33), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G159), .ZN(new_n306));
  AND2_X1   g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(KEYINPUT16), .B1(new_n301), .B2(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(KEYINPUT7), .A2(G20), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT73), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n311), .B1(new_n296), .B2(new_n297), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n262), .A2(new_n265), .A3(KEYINPUT73), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n310), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(G20), .B1(new_n262), .B2(new_n265), .ZN(new_n315));
  OAI21_X1  g0115(.A(G68), .B1(new_n315), .B2(new_n293), .ZN(new_n316));
  OAI211_X1 g0116(.A(KEYINPUT16), .B(new_n307), .C1(new_n314), .C2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n255), .A2(new_n212), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n260), .B(new_n285), .C1(new_n308), .C2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT17), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n304), .A2(new_n306), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n216), .B1(new_n298), .B2(KEYINPUT7), .ZN(new_n324));
  AND3_X1   g0124(.A1(new_n262), .A2(new_n265), .A3(KEYINPUT73), .ZN(new_n325));
  AOI21_X1  g0125(.A(KEYINPUT73), .B1(new_n262), .B2(new_n265), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n309), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n323), .B1(new_n324), .B2(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n256), .B1(new_n328), .B2(KEYINPUT16), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT16), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n216), .B1(new_n295), .B2(new_n299), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n330), .B1(new_n331), .B2(new_n323), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n259), .B1(new_n329), .B2(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(KEYINPUT17), .B1(new_n333), .B2(new_n285), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n249), .B1(new_n322), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT18), .ZN(new_n336));
  INV_X1    g0136(.A(G179), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n284), .A2(KEYINPUT76), .A3(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT76), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n274), .A2(new_n281), .A3(new_n277), .ZN(new_n340));
  INV_X1    g0140(.A(G169), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n340), .A2(G179), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n338), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n336), .B1(new_n344), .B2(new_n333), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n280), .B1(new_n270), .B2(new_n273), .ZN(new_n346));
  AND4_X1   g0146(.A1(KEYINPUT76), .A2(new_n346), .A3(new_n337), .A4(new_n277), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n284), .A2(new_n337), .ZN(new_n348));
  OAI21_X1  g0148(.A(KEYINPUT76), .B1(new_n284), .B2(G169), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n260), .B1(new_n308), .B2(new_n319), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n350), .A2(new_n351), .A3(KEYINPUT18), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n345), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n320), .A2(new_n321), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n333), .A2(KEYINPUT17), .A3(new_n285), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n354), .A2(new_n355), .A3(KEYINPUT77), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n335), .A2(new_n353), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT68), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n272), .A2(G238), .A3(new_n275), .ZN(new_n360));
  NOR2_X1   g0160(.A1(G226), .A2(G1698), .ZN(new_n361));
  INV_X1    g0161(.A(G232), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n361), .B1(new_n362), .B2(G1698), .ZN(new_n363));
  XNOR2_X1  g0163(.A(KEYINPUT3), .B(G33), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n363), .A2(new_n364), .B1(G33), .B2(G97), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n281), .B(new_n360), .C1(new_n365), .C2(new_n272), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(KEYINPUT13), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n262), .A2(new_n265), .ZN(new_n368));
  INV_X1    g0168(.A(G1698), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n266), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n362), .A2(G1698), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(G97), .ZN(new_n373));
  OAI22_X1  g0173(.A1(new_n368), .A2(new_n372), .B1(new_n261), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n280), .B1(new_n374), .B2(new_n273), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT13), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n375), .A2(new_n376), .A3(new_n360), .ZN(new_n377));
  AND2_X1   g0177(.A1(new_n367), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(G200), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n359), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n253), .A2(new_n216), .ZN(new_n381));
  XNOR2_X1  g0181(.A(new_n381), .B(KEYINPUT12), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT69), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n318), .B1(new_n251), .B2(G20), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n383), .B1(new_n384), .B2(G68), .ZN(new_n385));
  NOR3_X1   g0185(.A1(new_n258), .A2(KEYINPUT69), .A3(new_n216), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT11), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n305), .A2(G50), .B1(G20), .B2(new_n216), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n261), .A2(G20), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n388), .B1(new_n390), .B2(new_n203), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n387), .B1(new_n391), .B2(new_n318), .ZN(new_n392));
  AND3_X1   g0192(.A1(new_n391), .A2(new_n387), .A3(new_n318), .ZN(new_n393));
  OAI221_X1 g0193(.A(new_n382), .B1(new_n385), .B2(new_n386), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n394), .B1(new_n378), .B2(G190), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n367), .A2(new_n377), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n396), .A2(KEYINPUT68), .A3(G200), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n380), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(KEYINPUT70), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT70), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n380), .A2(new_n395), .A3(new_n400), .A4(new_n397), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n378), .A2(G179), .ZN(new_n403));
  OAI21_X1  g0203(.A(KEYINPUT71), .B1(new_n378), .B2(new_n341), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT72), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n341), .B1(new_n367), .B2(new_n377), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT71), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n404), .A2(new_n405), .A3(KEYINPUT14), .A4(new_n408), .ZN(new_n409));
  AND3_X1   g0209(.A1(new_n404), .A2(KEYINPUT14), .A3(new_n408), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT14), .ZN(new_n411));
  AOI21_X1  g0211(.A(KEYINPUT72), .B1(new_n406), .B2(new_n411), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n403), .B(new_n409), .C1(new_n410), .C2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n402), .B1(new_n413), .B2(new_n394), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n250), .A2(new_n389), .B1(G150), .B2(new_n305), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(new_n202), .B2(new_n211), .ZN(new_n416));
  INV_X1    g0216(.A(G50), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n416), .A2(new_n318), .B1(new_n417), .B2(new_n253), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n384), .A2(G50), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NOR2_X1   g0220(.A1(G222), .A2(G1698), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n369), .A2(G223), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n364), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n423), .B(new_n273), .C1(G77), .C2(new_n364), .ZN(new_n424));
  AND2_X1   g0224(.A1(new_n272), .A2(new_n275), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(G226), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n424), .A2(new_n281), .A3(new_n426), .ZN(new_n427));
  OR2_X1    g0227(.A1(new_n427), .A2(G179), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n341), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n420), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n425), .A2(G244), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n364), .A2(G232), .A3(new_n369), .ZN(new_n433));
  INV_X1    g0233(.A(G107), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n364), .A2(G1698), .ZN(new_n435));
  OAI221_X1 g0235(.A(new_n433), .B1(new_n434), .B2(new_n364), .C1(new_n435), .C2(new_n215), .ZN(new_n436));
  AOI211_X1 g0236(.A(new_n432), .B(new_n280), .C1(new_n436), .C2(new_n273), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(G190), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n250), .A2(new_n305), .B1(G20), .B2(G77), .ZN(new_n439));
  OR2_X1    g0239(.A1(KEYINPUT15), .A2(G87), .ZN(new_n440));
  NAND2_X1  g0240(.A1(KEYINPUT15), .A2(G87), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n439), .B1(new_n390), .B2(new_n442), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n443), .A2(new_n318), .B1(new_n203), .B2(new_n253), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n384), .A2(G77), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n438), .B(new_n447), .C1(new_n379), .C2(new_n437), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT9), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n420), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n427), .A2(G200), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n418), .A2(KEYINPUT9), .A3(new_n419), .ZN(new_n453));
  OR2_X1    g0253(.A1(new_n427), .A2(new_n278), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n451), .A2(new_n452), .A3(new_n453), .A4(new_n454), .ZN(new_n455));
  OR2_X1    g0255(.A1(new_n455), .A2(KEYINPUT10), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(KEYINPUT10), .ZN(new_n457));
  AOI211_X1 g0257(.A(new_n431), .B(new_n449), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n437), .A2(new_n337), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n459), .B(new_n446), .C1(G169), .C2(new_n437), .ZN(new_n460));
  AOI21_X1  g0260(.A(KEYINPUT67), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n457), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n455), .A2(KEYINPUT10), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n430), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT67), .ZN(new_n465));
  INV_X1    g0265(.A(new_n460), .ZN(new_n466));
  NOR4_X1   g0266(.A1(new_n464), .A2(new_n465), .A3(new_n466), .A4(new_n449), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n358), .B(new_n414), .C1(new_n461), .C2(new_n467), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n262), .A2(new_n265), .A3(G257), .A4(new_n369), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n262), .A2(new_n265), .A3(G264), .A4(G1698), .ZN(new_n470));
  INV_X1    g0270(.A(G303), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n469), .B(new_n470), .C1(new_n471), .C2(new_n364), .ZN(new_n472));
  XNOR2_X1  g0272(.A(KEYINPUT5), .B(G41), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n251), .A2(G45), .A3(G274), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT79), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT79), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n473), .A2(new_n475), .A3(new_n478), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n472), .A2(new_n273), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n473), .A2(new_n251), .A3(G45), .ZN(new_n481));
  AND2_X1   g0281(.A1(new_n481), .A2(new_n272), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G270), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(G116), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n255), .A2(new_n212), .B1(G20), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G283), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n488), .B(new_n211), .C1(G33), .C2(new_n373), .ZN(new_n489));
  AND3_X1   g0289(.A1(new_n487), .A2(KEYINPUT20), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(KEYINPUT20), .B1(new_n487), .B2(new_n489), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n252), .A2(G116), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n251), .A2(G33), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n252), .A2(new_n495), .A3(new_n212), .A4(new_n255), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n494), .B1(new_n486), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(KEYINPUT83), .B1(new_n492), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n487), .A2(new_n489), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT20), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n487), .A2(KEYINPUT20), .A3(new_n489), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n497), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT83), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n498), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n485), .A2(new_n507), .A3(G179), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n484), .A2(G200), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n480), .A2(new_n483), .A3(G190), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n509), .A2(new_n506), .A3(new_n498), .A4(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT21), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n341), .B1(new_n480), .B2(new_n483), .ZN(new_n513));
  AND3_X1   g0313(.A1(new_n507), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n512), .B1(new_n507), .B2(new_n513), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n508), .B(new_n511), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n262), .A2(new_n265), .A3(G244), .A4(new_n369), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT4), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n364), .A2(KEYINPUT4), .A3(G244), .A4(new_n369), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n364), .A2(G250), .A3(G1698), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n519), .A2(new_n520), .A3(new_n488), .A4(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n273), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n477), .A2(new_n479), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n482), .A2(G257), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G200), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n434), .B1(new_n295), .B2(new_n299), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n305), .A2(G77), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT6), .ZN(new_n530));
  NOR3_X1   g0330(.A1(new_n530), .A2(new_n373), .A3(G107), .ZN(new_n531));
  XNOR2_X1  g0331(.A(G97), .B(G107), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n531), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n529), .B1(new_n533), .B2(new_n211), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n318), .B1(new_n528), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n496), .A2(G97), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(G97), .B2(new_n253), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(KEYINPUT78), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT78), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n536), .B(new_n539), .C1(G97), .C2(new_n253), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n523), .A2(G190), .A3(new_n525), .A4(new_n524), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n527), .A2(new_n535), .A3(new_n541), .A4(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n526), .A2(new_n341), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n535), .A2(new_n541), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n523), .A2(new_n337), .A3(new_n525), .A4(new_n524), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n516), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n262), .A2(new_n265), .A3(G257), .A4(G1698), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n262), .A2(new_n265), .A3(G250), .A4(new_n369), .ZN(new_n551));
  NAND2_X1  g0351(.A1(G33), .A2(G294), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n273), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n481), .A2(G264), .A3(new_n272), .ZN(new_n555));
  AND3_X1   g0355(.A1(new_n554), .A2(KEYINPUT84), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(KEYINPUT84), .B1(new_n554), .B2(new_n555), .ZN(new_n557));
  OAI211_X1 g0357(.A(G179), .B(new_n524), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n554), .A2(new_n555), .ZN(new_n559));
  INV_X1    g0359(.A(new_n524), .ZN(new_n560));
  OAI21_X1  g0360(.A(G169), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n262), .A2(new_n265), .A3(new_n211), .A4(G87), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(KEYINPUT22), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT22), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n364), .A2(new_n565), .A3(new_n211), .A4(G87), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n389), .A2(G116), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n211), .A2(G107), .ZN(new_n569));
  XNOR2_X1  g0369(.A(new_n569), .B(KEYINPUT23), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n567), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT24), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n567), .A2(KEYINPUT24), .A3(new_n568), .A4(new_n570), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n573), .A2(new_n318), .A3(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(new_n496), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(G107), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n252), .A2(G107), .ZN(new_n578));
  XNOR2_X1  g0378(.A(new_n578), .B(KEYINPUT25), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n575), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n562), .A2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  NOR3_X1   g0382(.A1(new_n559), .A2(new_n560), .A3(G190), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n524), .B1(new_n556), .B2(new_n557), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n583), .B1(new_n584), .B2(new_n379), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n585), .A2(new_n580), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n211), .ZN(new_n589));
  INV_X1    g0389(.A(G87), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n590), .A2(new_n373), .A3(new_n434), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n262), .A2(new_n265), .A3(new_n211), .A4(G68), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n211), .A2(G33), .A3(G97), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT19), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n592), .A2(new_n593), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n318), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT80), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n252), .B1(new_n440), .B2(new_n441), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n598), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n589), .A2(new_n591), .B1(new_n594), .B2(new_n595), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n256), .B1(new_n603), .B2(new_n593), .ZN(new_n604));
  OAI21_X1  g0404(.A(KEYINPUT80), .B1(new_n604), .B2(new_n600), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n576), .A2(G87), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(G238), .A2(G1698), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n369), .A2(G244), .ZN(new_n610));
  NOR3_X1   g0410(.A1(new_n368), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n261), .A2(new_n486), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n273), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(G45), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n272), .B(G250), .C1(G1), .C2(new_n614), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n613), .A2(G190), .A3(new_n474), .A4(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n613), .A2(new_n474), .A3(new_n615), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(G200), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n608), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT82), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n496), .A2(new_n442), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(KEYINPUT81), .B1(new_n606), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT81), .ZN(new_n624));
  AOI211_X1 g0424(.A(new_n624), .B(new_n621), .C1(new_n602), .C2(new_n605), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n620), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n599), .B1(new_n598), .B2(new_n601), .ZN(new_n627));
  NOR3_X1   g0427(.A1(new_n604), .A2(KEYINPUT80), .A3(new_n600), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n622), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(new_n624), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n606), .A2(KEYINPUT81), .A3(new_n622), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n630), .A2(new_n631), .A3(KEYINPUT82), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n617), .A2(G169), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n633), .B1(new_n337), .B2(new_n617), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n626), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n549), .A2(new_n587), .A3(new_n619), .A4(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n468), .A2(new_n636), .ZN(G372));
  INV_X1    g0437(.A(new_n468), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n508), .B1(new_n514), .B2(new_n515), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT85), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  OAI211_X1 g0441(.A(KEYINPUT85), .B(new_n508), .C1(new_n514), .C2(new_n515), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n641), .A2(new_n581), .A3(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n634), .B1(new_n623), .B2(new_n625), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n619), .ZN(new_n645));
  NOR3_X1   g0445(.A1(new_n645), .A2(new_n586), .A3(new_n548), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n635), .A2(new_n619), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(KEYINPUT26), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT26), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n644), .A2(new_n651), .A3(new_n619), .A4(new_n648), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n647), .A2(new_n650), .A3(new_n644), .A4(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n638), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n335), .A2(new_n356), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n406), .B(KEYINPUT71), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n412), .B1(new_n656), .B2(KEYINPUT14), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n409), .A2(new_n403), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n394), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n466), .A2(new_n398), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n655), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n353), .ZN(new_n662));
  OAI22_X1  g0462(.A1(new_n661), .A2(new_n662), .B1(new_n462), .B2(new_n463), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n654), .A2(new_n430), .A3(new_n663), .ZN(G369));
  INV_X1    g0464(.A(G13), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n665), .A2(G20), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  OR3_X1    g0467(.A1(new_n667), .A2(KEYINPUT27), .A3(G1), .ZN(new_n668));
  OAI21_X1  g0468(.A(KEYINPUT27), .B1(new_n667), .B2(G1), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(G213), .A3(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(G343), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n507), .A2(new_n513), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(KEYINPUT21), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n507), .A2(new_n512), .A3(new_n513), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n672), .B1(new_n676), .B2(new_n508), .ZN(new_n677));
  INV_X1    g0477(.A(new_n672), .ZN(new_n678));
  AOI22_X1  g0478(.A1(new_n587), .A2(new_n677), .B1(new_n582), .B2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT88), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT86), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n516), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n676), .A2(KEYINPUT86), .A3(new_n508), .A4(new_n511), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n507), .A2(new_n672), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n684), .B1(new_n641), .B2(new_n642), .ZN(new_n686));
  OAI21_X1  g0486(.A(KEYINPUT87), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT87), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n641), .A2(new_n642), .ZN(new_n690));
  OAI211_X1 g0490(.A(new_n688), .B(new_n689), .C1(new_n690), .C2(new_n684), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n687), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(G330), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n580), .A2(new_n672), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n587), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(new_n581), .B2(new_n678), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n680), .B1(new_n693), .B2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NOR3_X1   g0499(.A1(new_n693), .A2(new_n680), .A3(new_n697), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n679), .B1(new_n699), .B2(new_n700), .ZN(G399));
  INV_X1    g0501(.A(new_n229), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(G41), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n591), .A2(G116), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n704), .A2(G1), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n210), .B2(new_n704), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT28), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n676), .A2(new_n581), .A3(new_n508), .ZN(new_n709));
  INV_X1    g0509(.A(new_n586), .ZN(new_n710));
  AND4_X1   g0510(.A1(new_n616), .A2(new_n618), .A3(new_n606), .A4(new_n607), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n630), .A2(new_n631), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n711), .B1(new_n712), .B2(new_n634), .ZN(new_n713));
  INV_X1    g0513(.A(new_n548), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n709), .A2(new_n710), .A3(new_n713), .A4(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n644), .A2(new_n619), .A3(new_n648), .ZN(new_n716));
  AOI22_X1  g0516(.A1(new_n716), .A2(KEYINPUT26), .B1(new_n712), .B2(new_n634), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n635), .A2(new_n651), .A3(new_n619), .A4(new_n648), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n715), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n719), .A2(KEYINPUT29), .A3(new_n678), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n652), .A2(new_n644), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n721), .B1(new_n643), .B2(new_n646), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n672), .B1(new_n722), .B2(new_n650), .ZN(new_n723));
  OAI211_X1 g0523(.A(KEYINPUT89), .B(new_n720), .C1(new_n723), .C2(KEYINPUT29), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n484), .A2(new_n617), .A3(new_n337), .ZN(new_n725));
  OR2_X1    g0525(.A1(new_n556), .A2(new_n557), .ZN(new_n726));
  INV_X1    g0526(.A(new_n526), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT30), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n725), .A2(new_n726), .A3(KEYINPUT30), .A4(new_n727), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n584), .A2(new_n337), .A3(new_n617), .A4(new_n526), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n730), .B(new_n731), .C1(new_n485), .C2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(new_n672), .ZN(new_n734));
  OAI211_X1 g0534(.A(new_n734), .B(KEYINPUT31), .C1(new_n636), .C2(new_n672), .ZN(new_n735));
  OR2_X1    g0535(.A1(new_n734), .A2(KEYINPUT31), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n735), .A2(G330), .A3(new_n736), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n720), .A2(KEYINPUT89), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n724), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(KEYINPUT90), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT90), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n724), .A2(new_n738), .A3(new_n741), .A4(new_n737), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n708), .B1(new_n743), .B2(G1), .ZN(G364));
  AOI21_X1  g0544(.A(new_n251), .B1(new_n666), .B2(G45), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n703), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n747), .B1(new_n692), .B2(G330), .ZN(new_n748));
  OR2_X1    g0548(.A1(new_n692), .A2(G330), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G13), .A2(G33), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(G20), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n688), .B(new_n752), .C1(new_n690), .C2(new_n684), .ZN(new_n753));
  INV_X1    g0553(.A(new_n747), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n212), .B1(G20), .B2(new_n341), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n211), .A2(G179), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G190), .A2(G200), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(G329), .ZN(new_n760));
  INV_X1    g0560(.A(G311), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n211), .A2(new_n337), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(new_n758), .ZN(new_n763));
  OAI221_X1 g0563(.A(new_n368), .B1(new_n759), .B2(new_n760), .C1(new_n761), .C2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n762), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n765), .A2(new_n278), .A3(G200), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(G322), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n757), .A2(G190), .A3(G200), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n767), .A2(new_n768), .B1(new_n769), .B2(new_n471), .ZN(new_n770));
  NOR3_X1   g0570(.A1(new_n765), .A2(new_n379), .A3(G190), .ZN(new_n771));
  XNOR2_X1  g0571(.A(KEYINPUT33), .B(G317), .ZN(new_n772));
  AOI211_X1 g0572(.A(new_n764), .B(new_n770), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  NOR3_X1   g0573(.A1(new_n278), .A2(G179), .A3(G200), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n211), .ZN(new_n775));
  INV_X1    g0575(.A(G294), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n762), .A2(G190), .A3(G200), .ZN(new_n777));
  INV_X1    g0577(.A(G326), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n775), .A2(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT92), .ZN(new_n780));
  INV_X1    g0580(.A(G283), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n757), .A2(new_n278), .A3(G200), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n773), .B(new_n780), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(G159), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n759), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(KEYINPUT32), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n785), .A2(new_n786), .B1(new_n434), .B2(new_n782), .ZN(new_n787));
  INV_X1    g0587(.A(new_n771), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n788), .A2(new_n216), .B1(new_n763), .B2(new_n203), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n787), .B(new_n789), .C1(G58), .C2(new_n766), .ZN(new_n790));
  INV_X1    g0590(.A(new_n777), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G50), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n368), .B1(new_n785), .B2(new_n786), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n769), .A2(new_n590), .ZN(new_n794));
  XOR2_X1   g0594(.A(new_n775), .B(KEYINPUT91), .Z(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n794), .B1(new_n796), .B2(G97), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n790), .A2(new_n792), .A3(new_n793), .A4(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n756), .B1(new_n783), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n752), .A2(new_n755), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n244), .A2(G45), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n325), .A2(new_n326), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(new_n702), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n801), .B(new_n803), .C1(G45), .C2(new_n210), .ZN(new_n804));
  INV_X1    g0604(.A(G355), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n364), .A2(new_n229), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n804), .B1(G116), .B2(new_n229), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n754), .B(new_n799), .C1(new_n800), .C2(new_n807), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n748), .A2(new_n749), .B1(new_n753), .B2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(G396));
  OAI21_X1  g0610(.A(new_n448), .B1(new_n447), .B2(new_n678), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(new_n460), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n460), .A2(new_n672), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n723), .B(new_n815), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(new_n737), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(new_n754), .ZN(new_n818));
  OR2_X1    g0618(.A1(new_n771), .A2(KEYINPUT93), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n771), .A2(KEYINPUT93), .ZN(new_n820));
  AND2_X1   g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n763), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n821), .A2(G283), .B1(G116), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n823), .A2(KEYINPUT94), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n364), .B(new_n824), .C1(G303), .C2(new_n791), .ZN(new_n825));
  INV_X1    g0625(.A(new_n769), .ZN(new_n826));
  INV_X1    g0626(.A(new_n759), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n826), .A2(G107), .B1(new_n827), .B2(G311), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n795), .A2(new_n373), .B1(new_n776), .B2(new_n767), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT95), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n782), .A2(new_n590), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(new_n823), .B2(KEYINPUT94), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n825), .A2(new_n828), .A3(new_n831), .A4(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n829), .A2(new_n830), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n766), .A2(G143), .B1(new_n791), .B2(G137), .ZN(new_n836));
  INV_X1    g0636(.A(G150), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n836), .B1(new_n837), .B2(new_n788), .C1(new_n784), .C2(new_n763), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT34), .ZN(new_n839));
  OR2_X1    g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n838), .A2(new_n839), .B1(G132), .B2(new_n827), .ZN(new_n841));
  INV_X1    g0641(.A(new_n782), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(G68), .ZN(new_n843));
  INV_X1    g0643(.A(new_n775), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n844), .A2(G58), .B1(new_n826), .B2(G50), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n840), .A2(new_n841), .A3(new_n843), .A4(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n802), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n834), .A2(new_n835), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(new_n755), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n754), .B1(new_n815), .B2(new_n750), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n755), .A2(new_n750), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n849), .B(new_n850), .C1(G77), .C2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n818), .A2(new_n853), .ZN(G384));
  INV_X1    g0654(.A(KEYINPUT35), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n211), .B(new_n212), .C1(new_n533), .C2(new_n855), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n856), .B(G116), .C1(new_n855), .C2(new_n533), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n857), .B(KEYINPUT36), .ZN(new_n858));
  OAI21_X1  g0658(.A(G77), .B1(new_n302), .B2(new_n216), .ZN(new_n859));
  OAI22_X1  g0659(.A1(new_n210), .A2(new_n859), .B1(G50), .B2(new_n216), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n860), .A2(G1), .A3(new_n665), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT97), .ZN(new_n862));
  INV_X1    g0662(.A(new_n317), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n307), .B1(new_n314), .B2(new_n316), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n256), .B1(new_n864), .B2(new_n330), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT96), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n863), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n318), .B1(new_n328), .B2(KEYINPUT16), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(KEYINPUT96), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n259), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n862), .B1(new_n870), .B2(new_n670), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n317), .B1(new_n868), .B2(KEYINPUT96), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n865), .A2(new_n866), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n260), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n670), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n874), .A2(KEYINPUT97), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n871), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n357), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT98), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n357), .A2(KEYINPUT98), .A3(new_n877), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n350), .A2(new_n351), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n351), .A2(new_n875), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT37), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n883), .A2(new_n884), .A3(new_n885), .A4(new_n320), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(KEYINPUT99), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n351), .B1(new_n350), .B2(new_n875), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT99), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n888), .A2(new_n889), .A3(new_n885), .A4(new_n320), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n320), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n892), .B1(new_n874), .B2(new_n350), .ZN(new_n893));
  AND3_X1   g0693(.A1(new_n893), .A2(new_n871), .A3(new_n876), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n891), .B1(new_n894), .B2(new_n885), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT38), .B1(new_n882), .B2(new_n895), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n357), .A2(KEYINPUT98), .A3(new_n877), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT98), .B1(new_n357), .B2(new_n877), .ZN(new_n898));
  OAI211_X1 g0698(.A(KEYINPUT38), .B(new_n895), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  OAI211_X1 g0700(.A(KEYINPUT100), .B(KEYINPUT39), .C1(new_n896), .C2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n902), .A2(new_n351), .A3(new_n875), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n887), .A2(new_n890), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n329), .A2(new_n332), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n344), .A2(new_n670), .B1(new_n905), .B2(new_n260), .ZN(new_n906));
  OAI21_X1  g0706(.A(KEYINPUT37), .B1(new_n906), .B2(new_n892), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT101), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI211_X1 g0709(.A(KEYINPUT101), .B(KEYINPUT37), .C1(new_n906), .C2(new_n892), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n903), .B1(new_n904), .B2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT38), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT39), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n899), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n916), .A2(KEYINPUT100), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n895), .B1(new_n897), .B2(new_n898), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n913), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n915), .B1(new_n919), .B2(new_n899), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n901), .B1(new_n917), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n413), .A2(new_n394), .A3(new_n678), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT102), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n919), .A2(new_n899), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n394), .A2(new_n672), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n659), .A2(new_n398), .A3(new_n927), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n394), .B(new_n672), .C1(new_n413), .C2(new_n402), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n815), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n653), .A2(new_n678), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n930), .B1(new_n932), .B2(new_n814), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n926), .A2(new_n933), .B1(new_n662), .B2(new_n670), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n924), .A2(new_n925), .A3(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(KEYINPUT39), .B1(new_n896), .B2(new_n900), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n916), .A2(KEYINPUT100), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n922), .B1(new_n938), .B2(new_n901), .ZN(new_n939));
  INV_X1    g0739(.A(new_n934), .ZN(new_n940));
  OAI21_X1  g0740(.A(KEYINPUT102), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n935), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n468), .B1(new_n724), .B2(new_n738), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n663), .A2(new_n430), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n942), .B(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n928), .A2(new_n929), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n947), .A2(new_n735), .A3(new_n736), .A4(new_n931), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n948), .B1(new_n919), .B2(new_n899), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n949), .A2(KEYINPUT40), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n735), .A2(new_n736), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n930), .A2(new_n815), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n899), .A2(new_n914), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n952), .A2(new_n953), .A3(KEYINPUT40), .A4(new_n951), .ZN(new_n954));
  NAND4_X1  g0754(.A1(new_n950), .A2(new_n638), .A3(new_n951), .A4(new_n954), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n954), .B(G330), .C1(new_n949), .C2(KEYINPUT40), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n468), .A2(new_n737), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n955), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n946), .A2(new_n959), .B1(new_n251), .B2(new_n666), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n960), .B(KEYINPUT103), .Z(new_n961));
  NAND2_X1  g0761(.A1(new_n946), .A2(new_n959), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n962), .B(KEYINPUT104), .Z(new_n963));
  OAI211_X1 g0763(.A(new_n858), .B(new_n861), .C1(new_n961), .C2(new_n963), .ZN(G367));
  INV_X1    g0764(.A(new_n803), .ZN(new_n965));
  OAI221_X1 g0765(.A(new_n800), .B1(new_n229), .B2(new_n442), .C1(new_n965), .C2(new_n240), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n766), .A2(G303), .B1(new_n791), .B2(G311), .ZN(new_n967));
  INV_X1    g0767(.A(new_n821), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n967), .B1(new_n968), .B2(new_n776), .ZN(new_n969));
  OAI21_X1  g0769(.A(KEYINPUT107), .B1(new_n769), .B2(new_n486), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n970), .A2(KEYINPUT46), .B1(new_n844), .B2(G107), .ZN(new_n971));
  AOI22_X1  g0771(.A1(G283), .A2(new_n822), .B1(new_n827), .B2(G317), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n971), .B(new_n972), .C1(KEYINPUT46), .C2(new_n970), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n782), .A2(new_n373), .ZN(new_n974));
  NOR4_X1   g0774(.A1(new_n969), .A2(new_n973), .A3(new_n802), .A4(new_n974), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT108), .Z(new_n976));
  OAI221_X1 g0776(.A(new_n364), .B1(new_n837), .B2(new_n767), .C1(new_n968), .C2(new_n784), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(G137), .B2(new_n827), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n822), .A2(G50), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n782), .A2(new_n203), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n769), .A2(new_n302), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n795), .A2(new_n216), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n982), .B(new_n983), .C1(G143), .C2(new_n791), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n978), .A2(new_n979), .A3(new_n981), .A4(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n976), .A2(new_n985), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n986), .B(KEYINPUT47), .Z(new_n987));
  OAI211_X1 g0787(.A(new_n747), .B(new_n966), .C1(new_n987), .C2(new_n756), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n713), .B1(new_n608), .B2(new_n678), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n608), .A2(new_n678), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n989), .B1(new_n644), .B2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n752), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n988), .A2(new_n993), .ZN(new_n994));
  AND2_X1   g0794(.A1(new_n740), .A2(new_n742), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n587), .A2(new_n677), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n696), .B2(new_n677), .ZN(new_n997));
  AND3_X1   g0797(.A1(new_n692), .A2(G330), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n997), .B1(new_n692), .B2(G330), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(KEYINPUT106), .B1(new_n743), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT106), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n1003), .B(new_n1000), .C1(new_n740), .C2(new_n742), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n700), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n545), .A2(new_n672), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n714), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(new_n547), .B2(new_n678), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n679), .A2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT45), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n679), .A2(new_n1009), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT44), .Z(new_n1013));
  OAI211_X1 g0813(.A(new_n1006), .B(new_n698), .C1(new_n1011), .C2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1013), .A2(new_n1011), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n699), .B2(new_n700), .ZN(new_n1016));
  AND2_X1   g0816(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n995), .B1(new_n1005), .B2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n703), .B(KEYINPUT41), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n745), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n996), .A2(new_n1008), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1022), .A2(KEYINPUT42), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(KEYINPUT42), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n547), .B1(new_n1008), .B2(new_n581), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n1023), .A2(new_n1024), .B1(new_n678), .B2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n991), .A2(KEYINPUT43), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT105), .ZN(new_n1029));
  AND2_X1   g0829(.A1(new_n991), .A2(KEYINPUT43), .ZN(new_n1030));
  NOR3_X1   g0830(.A1(new_n1026), .A2(new_n1027), .A3(new_n1030), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1006), .A2(new_n698), .A3(new_n1009), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1032), .B(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n994), .B1(new_n1021), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1036), .ZN(G387));
  NAND2_X1  g0837(.A1(new_n697), .A2(new_n752), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n250), .A2(new_n417), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT50), .Z(new_n1040));
  OAI21_X1  g0840(.A(new_n614), .B1(new_n216), .B2(new_n203), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n705), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT109), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1041), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1040), .B(new_n1044), .C1(new_n1043), .C2(new_n1042), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1045), .B(new_n803), .C1(new_n237), .C2(new_n614), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(G107), .B2(new_n229), .C1(new_n705), .C2(new_n806), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n754), .B1(new_n1047), .B2(new_n800), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n769), .A2(new_n203), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n795), .A2(new_n442), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1049), .B(new_n1050), .C1(G68), .C2(new_n822), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n802), .B1(new_n784), .B2(new_n777), .C1(new_n767), .C2(new_n417), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n974), .B(new_n1052), .C1(new_n250), .C2(new_n771), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1051), .B(new_n1053), .C1(new_n837), .C2(new_n759), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n766), .A2(G317), .B1(G303), .B2(new_n822), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1055), .B1(new_n768), .B2(new_n777), .C1(new_n968), .C2(new_n761), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT48), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1057), .B1(new_n781), .B2(new_n775), .C1(new_n776), .C2(new_n769), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT49), .Z(new_n1059));
  OAI221_X1 g0859(.A(new_n847), .B1(new_n486), .B2(new_n782), .C1(new_n778), .C2(new_n759), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT110), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1054), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  XOR2_X1   g0862(.A(new_n1062), .B(KEYINPUT111), .Z(new_n1063));
  OAI211_X1 g0863(.A(new_n1038), .B(new_n1048), .C1(new_n1063), .C2(new_n756), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n995), .A2(new_n1000), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n703), .B1(new_n743), .B2(new_n1001), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1064), .B1(new_n745), .B2(new_n1000), .C1(new_n1065), .C2(new_n1066), .ZN(G393));
  OAI21_X1  g0867(.A(new_n1003), .B1(new_n995), .B2(new_n1000), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n743), .A2(KEYINPUT106), .A3(new_n1001), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1068), .A2(new_n1017), .A3(new_n1069), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1070), .B(new_n703), .C1(new_n1017), .C2(new_n1065), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n800), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n229), .A2(new_n373), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1072), .B(new_n1073), .C1(new_n803), .C2(new_n247), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n250), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n968), .A2(new_n417), .B1(new_n1075), .B2(new_n763), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n795), .A2(new_n203), .ZN(new_n1077));
  NOR3_X1   g0877(.A1(new_n1076), .A2(new_n1077), .A3(new_n832), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n827), .A2(G143), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n826), .A2(G68), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n766), .A2(G159), .B1(new_n791), .B2(G150), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT51), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1082), .A2(new_n847), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n1078), .A2(new_n1079), .A3(new_n1080), .A4(new_n1083), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n844), .A2(G116), .B1(new_n822), .B2(G294), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n968), .B2(new_n471), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT114), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(G107), .B2(new_n842), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n827), .A2(G322), .ZN(new_n1089));
  INV_X1    g0889(.A(G317), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n767), .A2(new_n761), .B1(new_n777), .B2(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n364), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  OR2_X1    g0893(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1088), .A2(new_n1089), .A3(new_n1093), .A4(new_n1094), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n769), .A2(new_n781), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1084), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n754), .B(new_n1074), .C1(new_n1097), .C2(new_n755), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1009), .A2(new_n992), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT112), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n1017), .A2(new_n746), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1071), .A2(new_n1101), .ZN(G390));
  NAND3_X1  g0902(.A1(new_n719), .A2(new_n678), .A3(new_n812), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n814), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT115), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1103), .A2(KEYINPUT115), .A3(new_n814), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n947), .A2(KEYINPUT116), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT116), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n928), .A2(new_n929), .A3(new_n1110), .ZN(new_n1111));
  AND2_X1   g0911(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n953), .B(new_n922), .C1(new_n1108), .C2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT117), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n933), .B2(new_n923), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n813), .B1(new_n723), .B2(new_n931), .ZN(new_n1116));
  OAI211_X1 g0916(.A(KEYINPUT117), .B(new_n922), .C1(new_n1116), .C2(new_n930), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1113), .B1(new_n921), .B2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n735), .A2(G330), .A3(new_n736), .A4(new_n931), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1120), .A2(new_n930), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n938), .A2(new_n901), .A3(new_n1115), .A4(new_n1117), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n951), .A2(G330), .A3(new_n931), .A4(new_n947), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1123), .A2(new_n1113), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT118), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1116), .ZN(new_n1127));
  AND2_X1   g0927(.A1(new_n1120), .A2(new_n930), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1127), .B1(new_n1128), .B2(new_n1121), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1120), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1108), .A2(new_n1124), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  NOR3_X1   g0932(.A1(new_n943), .A2(new_n944), .A3(new_n958), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n1126), .B(new_n704), .C1(new_n1132), .C2(new_n1133), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1122), .B(new_n1125), .C1(new_n1134), .C2(new_n746), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(KEYINPUT118), .ZN(new_n1137));
  AND3_X1   g0937(.A1(new_n1123), .A2(new_n1113), .A3(new_n1124), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1124), .B1(new_n1123), .B2(new_n1113), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n703), .B(new_n1137), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n754), .B1(new_n1075), .B2(new_n851), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n821), .A2(G137), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n826), .A2(G150), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1142), .B1(KEYINPUT53), .B2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(KEYINPUT53), .B2(new_n1143), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n796), .A2(G159), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n766), .A2(G132), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(G128), .A2(new_n791), .B1(new_n842), .B2(G50), .ZN(new_n1148));
  XOR2_X1   g0948(.A(KEYINPUT54), .B(G143), .Z(new_n1149));
  AOI22_X1  g0949(.A1(new_n822), .A2(new_n1149), .B1(new_n827), .B2(G125), .ZN(new_n1150));
  AND3_X1   g0950(.A1(new_n1148), .A2(new_n364), .A3(new_n1150), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .A4(new_n1151), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n794), .B(new_n1077), .C1(G107), .C2(new_n821), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n843), .B1(new_n781), .B2(new_n777), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n763), .A2(new_n373), .B1(new_n759), .B2(new_n776), .ZN(new_n1155));
  NOR3_X1   g0955(.A1(new_n1154), .A2(new_n1155), .A3(new_n364), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1153), .B(new_n1156), .C1(new_n486), .C2(new_n767), .ZN(new_n1157));
  AND2_X1   g0957(.A1(new_n1152), .A2(new_n1157), .ZN(new_n1158));
  OAI221_X1 g0958(.A(new_n1141), .B1(new_n756), .B2(new_n1158), .C1(new_n921), .C2(new_n751), .ZN(new_n1159));
  AND3_X1   g0959(.A1(new_n1135), .A2(new_n1140), .A3(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(G378));
  NAND2_X1  g0961(.A1(new_n420), .A2(new_n875), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n464), .B(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1164));
  OR2_X1    g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT120), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1165), .A2(KEYINPUT120), .A3(new_n1166), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n957), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n956), .A2(new_n1166), .A3(new_n1165), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n925), .B1(new_n924), .B2(new_n934), .ZN(new_n1175));
  NOR3_X1   g0975(.A1(new_n939), .A2(KEYINPUT102), .A3(new_n940), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1174), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n935), .A2(new_n941), .A3(new_n1172), .A4(new_n1173), .ZN(new_n1178));
  AND2_X1   g0978(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1179));
  NOR3_X1   g0979(.A1(new_n1138), .A2(new_n1139), .A3(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1133), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1177), .B(new_n1178), .C1(new_n1180), .C2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT57), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n704), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1122), .A2(new_n1125), .A3(new_n1132), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n1133), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1186), .A2(KEYINPUT57), .A3(new_n1178), .A4(new_n1177), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1184), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1177), .A2(new_n746), .A3(new_n1178), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n842), .A2(G58), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1190), .B(KEYINPUT119), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n802), .B(new_n1191), .C1(G116), .C2(new_n791), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1049), .B1(G283), .B2(new_n827), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1193), .B1(new_n373), .B2(new_n788), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n767), .A2(new_n434), .ZN(new_n1195));
  NOR4_X1   g0995(.A1(new_n983), .A2(new_n1194), .A3(G41), .A4(new_n1195), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1192), .B(new_n1196), .C1(new_n442), .C2(new_n763), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT58), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n796), .A2(G150), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n766), .A2(G128), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n791), .A2(G125), .B1(new_n822), .B2(G137), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n771), .A2(G132), .B1(new_n826), .B2(new_n1149), .ZN(new_n1202));
  AND4_X1   g1002(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .A4(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT59), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n271), .B1(new_n782), .B2(new_n784), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(G124), .B2(new_n827), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1204), .A2(new_n261), .A3(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(G41), .B1(new_n802), .B2(G33), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1198), .B(new_n1207), .C1(G50), .C2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n754), .B1(new_n1209), .B2(new_n755), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1210), .B1(G50), .B2(new_n852), .C1(new_n1171), .C2(new_n751), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1189), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1188), .A2(new_n1213), .ZN(G375));
  NAND2_X1  g1014(.A1(new_n1112), .A2(new_n750), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n851), .A2(new_n216), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n364), .B1(new_n821), .B2(G116), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1217), .B1(new_n373), .B2(new_n769), .C1(new_n776), .C2(new_n777), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n980), .B(new_n1218), .C1(G283), .C2(new_n766), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n763), .A2(new_n434), .B1(new_n759), .B2(new_n471), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1050), .A2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n766), .A2(G137), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n796), .A2(G50), .B1(G159), .B2(new_n826), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n821), .A2(new_n1149), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n791), .A2(G132), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1223), .A2(new_n1224), .A3(new_n802), .A4(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(G128), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n763), .A2(new_n837), .B1(new_n759), .B2(new_n1227), .ZN(new_n1228));
  NOR3_X1   g1028(.A1(new_n1226), .A2(new_n1191), .A3(new_n1228), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n1219), .A2(new_n1221), .B1(new_n1222), .B2(new_n1229), .ZN(new_n1230));
  XOR2_X1   g1030(.A(new_n1230), .B(KEYINPUT121), .Z(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n755), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1215), .A2(new_n747), .A3(new_n1216), .A4(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1233), .B1(new_n1179), .B2(new_n745), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT122), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(new_n1234), .B(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1181), .A2(new_n1179), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1237), .A2(new_n1019), .A3(new_n1136), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1236), .A2(new_n1238), .ZN(G381));
  AOI21_X1  g1039(.A(new_n1212), .B1(new_n1184), .B2(new_n1187), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n1160), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(G384), .ZN(new_n1243));
  INV_X1    g1043(.A(G381), .ZN(new_n1244));
  NOR4_X1   g1044(.A1(G387), .A2(G396), .A3(G393), .A4(G390), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .A4(new_n1245), .ZN(G407));
  INV_X1    g1046(.A(G213), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1247), .A2(G343), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1241), .A2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1247), .B1(new_n1250), .B2(KEYINPUT123), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT123), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(new_n1241), .B2(new_n1249), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1251), .A2(G407), .A3(new_n1253), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(new_n1254), .B(KEYINPUT124), .ZN(G409));
  NAND4_X1  g1055(.A1(new_n1186), .A2(new_n1019), .A3(new_n1178), .A4(new_n1177), .ZN(new_n1256));
  AND2_X1   g1056(.A1(new_n1256), .A2(new_n1160), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1248), .B1(new_n1257), .B2(new_n1213), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1258), .B1(new_n1160), .B2(new_n1240), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT60), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1237), .A2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1181), .A2(new_n1179), .A3(KEYINPUT60), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1261), .A2(new_n703), .A3(new_n1136), .A4(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1236), .A2(G384), .A3(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(G384), .B1(new_n1236), .B2(new_n1263), .ZN(new_n1266));
  OAI211_X1 g1066(.A(G2897), .B(new_n1248), .C1(new_n1265), .C2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1266), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1248), .A2(G2897), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1268), .A2(new_n1264), .A3(new_n1269), .ZN(new_n1270));
  AND2_X1   g1070(.A1(new_n1267), .A2(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(KEYINPUT61), .B1(new_n1259), .B2(new_n1271), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1273));
  OAI211_X1 g1073(.A(new_n1258), .B(new_n1273), .C1(new_n1160), .C2(new_n1240), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(KEYINPUT62), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(G375), .A2(G378), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT62), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1276), .A2(new_n1277), .A3(new_n1273), .A4(new_n1258), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1272), .A2(new_n1275), .A3(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT126), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(G390), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1070), .A2(new_n743), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n1019), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1034), .B1(new_n1284), .B2(new_n745), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1282), .B1(new_n1285), .B2(new_n994), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1036), .A2(G390), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(G393), .B(G396), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1286), .A2(new_n1287), .A3(KEYINPUT125), .A4(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT125), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1291), .B1(new_n1036), .B2(G390), .ZN(new_n1292));
  AOI22_X1  g1092(.A1(new_n1292), .A2(new_n1288), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1290), .A2(new_n1293), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1272), .A2(new_n1275), .A3(new_n1278), .A4(KEYINPUT126), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1281), .A2(new_n1294), .A3(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT63), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1297), .B1(new_n1259), .B2(new_n1271), .ZN(new_n1298));
  MUX2_X1   g1098(.A(new_n1297), .B(new_n1298), .S(new_n1274), .Z(new_n1299));
  NOR2_X1   g1099(.A1(new_n1294), .A2(KEYINPUT61), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1296), .A2(new_n1301), .ZN(G405));
  NAND2_X1  g1102(.A1(new_n1276), .A2(new_n1241), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT127), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1304), .B1(new_n1290), .B2(new_n1293), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1292), .A2(new_n1288), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1308), .A2(KEYINPUT127), .A3(new_n1289), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1273), .ZN(new_n1310));
  AND3_X1   g1110(.A1(new_n1305), .A2(new_n1309), .A3(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1310), .B1(new_n1305), .B2(new_n1309), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1303), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1305), .A2(new_n1309), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(new_n1273), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1303), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1305), .A2(new_n1309), .A3(new_n1310), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1315), .A2(new_n1316), .A3(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1313), .A2(new_n1318), .ZN(G402));
endmodule


