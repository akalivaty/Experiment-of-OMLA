//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 1 1 0 0 1 1 0 0 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 0 1 1 0 1 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:02 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  INV_X1    g0014(.A(G97), .ZN(new_n215));
  INV_X1    g0015(.A(G257), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n211), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  OR2_X1    g0021(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n206), .A2(new_n207), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n211), .A2(G13), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n228), .B(G250), .C1(G257), .C2(G264), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT0), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n222), .A2(new_n227), .A3(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n221), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT2), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XOR2_X1   g0036(.A(G250), .B(G257), .Z(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT65), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(G1), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n249), .A2(G13), .A3(G20), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT66), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND4_X1  g0052(.A1(new_n249), .A2(KEYINPUT66), .A3(G13), .A4(G20), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NOR3_X1   g0054(.A1(new_n254), .A2(KEYINPUT12), .A3(G68), .ZN(new_n255));
  XOR2_X1   g0055(.A(new_n255), .B(KEYINPUT71), .Z(new_n256));
  OAI21_X1  g0056(.A(KEYINPUT12), .B1(new_n254), .B2(G68), .ZN(new_n257));
  XOR2_X1   g0057(.A(new_n257), .B(KEYINPUT72), .Z(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(new_n224), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n254), .B(new_n262), .C1(G1), .C2(new_n225), .ZN(new_n263));
  OR2_X1    g0063(.A1(new_n263), .A2(new_n203), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G20), .A2(G33), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  OAI22_X1  g0066(.A1(new_n266), .A2(new_n207), .B1(new_n225), .B2(G68), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n225), .A2(G33), .ZN(new_n268));
  INV_X1    g0068(.A(G77), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n261), .B1(new_n267), .B2(new_n270), .ZN(new_n271));
  XNOR2_X1  g0071(.A(KEYINPUT70), .B(KEYINPUT11), .ZN(new_n272));
  XNOR2_X1  g0072(.A(new_n271), .B(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n259), .A2(new_n264), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n224), .B1(G33), .B2(G41), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n249), .B1(G41), .B2(G45), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G238), .ZN(new_n279));
  INV_X1    g0079(.A(G274), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  OAI22_X1  g0082(.A1(new_n278), .A2(new_n279), .B1(KEYINPUT69), .B2(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n283), .B1(KEYINPUT69), .B2(new_n282), .ZN(new_n284));
  INV_X1    g0084(.A(G1698), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT3), .ZN(new_n286));
  INV_X1    g0086(.A(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(KEYINPUT3), .A2(G33), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n285), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G232), .ZN(new_n291));
  NAND2_X1  g0091(.A1(G33), .A2(G97), .ZN(new_n292));
  INV_X1    g0092(.A(G226), .ZN(new_n293));
  XNOR2_X1  g0093(.A(KEYINPUT3), .B(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n285), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n291), .B(new_n292), .C1(new_n293), .C2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n275), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n284), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(KEYINPUT13), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT13), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n284), .A2(new_n300), .A3(new_n297), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G169), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n303), .B1(KEYINPUT73), .B2(KEYINPUT14), .ZN(new_n304));
  NOR2_X1   g0104(.A1(KEYINPUT73), .A2(KEYINPUT14), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n302), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n299), .A2(G179), .A3(new_n301), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n305), .B1(new_n302), .B2(new_n304), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n274), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n290), .A2(G223), .ZN(new_n311));
  INV_X1    g0111(.A(G222), .ZN(new_n312));
  OAI221_X1 g0112(.A(new_n311), .B1(new_n269), .B2(new_n294), .C1(new_n312), .C2(new_n295), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(new_n275), .ZN(new_n314));
  INV_X1    g0114(.A(new_n278), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n281), .B1(new_n315), .B2(G226), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g0117(.A(KEYINPUT67), .B(G179), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n319), .B1(G169), .B2(new_n317), .ZN(new_n320));
  INV_X1    g0120(.A(new_n254), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n321), .A2(G50), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n322), .B1(G50), .B2(new_n263), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n208), .A2(G20), .ZN(new_n324));
  XNOR2_X1  g0124(.A(KEYINPUT8), .B(G58), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n268), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n326), .A2(new_n327), .B1(G150), .B2(new_n265), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n262), .B1(new_n324), .B2(new_n328), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n323), .A2(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n320), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(KEYINPUT9), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n317), .A2(G200), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT9), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n334), .B1(new_n323), .B2(new_n329), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n314), .A2(G190), .A3(new_n316), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n332), .A2(new_n333), .A3(new_n335), .A4(new_n336), .ZN(new_n337));
  OR2_X1    g0137(.A1(new_n337), .A2(KEYINPUT10), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(KEYINPUT10), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n331), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G200), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n302), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(G190), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n299), .A2(new_n343), .A3(new_n301), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n274), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  OR2_X1    g0146(.A1(new_n263), .A2(new_n269), .ZN(new_n347));
  XOR2_X1   g0147(.A(KEYINPUT15), .B(G87), .Z(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  OAI22_X1  g0149(.A1(new_n349), .A2(new_n268), .B1(new_n225), .B2(new_n269), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n325), .A2(new_n266), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n261), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n321), .A2(new_n269), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n347), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT68), .ZN(new_n355));
  OR2_X1    g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n354), .A2(new_n355), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n281), .B1(new_n315), .B2(G244), .ZN(new_n359));
  INV_X1    g0159(.A(G232), .ZN(new_n360));
  INV_X1    g0160(.A(G107), .ZN(new_n361));
  OAI22_X1  g0161(.A1(new_n295), .A2(new_n360), .B1(new_n361), .B2(new_n294), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n362), .B1(G238), .B2(new_n290), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n359), .B1(new_n363), .B2(new_n276), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(G169), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n365), .B1(new_n318), .B2(new_n364), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n358), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n364), .A2(new_n341), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n368), .B1(G190), .B2(new_n364), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n369), .A2(new_n357), .A3(new_n356), .ZN(new_n370));
  AND2_X1   g0170(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n310), .A2(new_n340), .A3(new_n346), .A4(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n290), .A2(KEYINPUT75), .A3(G226), .ZN(new_n373));
  AND2_X1   g0173(.A1(KEYINPUT3), .A2(G33), .ZN(new_n374));
  NOR2_X1   g0174(.A1(KEYINPUT3), .A2(G33), .ZN(new_n375));
  OAI211_X1 g0175(.A(G226), .B(G1698), .C1(new_n374), .C2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT75), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(G33), .A2(G87), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n294), .A2(G223), .A3(new_n285), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n373), .A2(new_n378), .A3(new_n379), .A4(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(new_n275), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n282), .B1(new_n278), .B2(new_n360), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n318), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n382), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n383), .B1(new_n381), .B2(new_n275), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n386), .B1(new_n387), .B2(new_n303), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n374), .A2(new_n375), .ZN(new_n389));
  AOI21_X1  g0189(.A(KEYINPUT7), .B1(new_n389), .B2(new_n225), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n288), .A2(KEYINPUT7), .A3(new_n225), .A4(new_n289), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(G68), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(G159), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n266), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(G58), .A2(G68), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n204), .A2(new_n205), .A3(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT74), .ZN(new_n400));
  AND3_X1   g0200(.A1(new_n399), .A2(new_n400), .A3(G20), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n400), .B1(new_n399), .B2(G20), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(KEYINPUT16), .B1(new_n397), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n288), .A2(new_n225), .A3(new_n289), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT7), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n391), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n395), .B1(new_n408), .B2(G68), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n399), .A2(G20), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT74), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n399), .A2(new_n400), .A3(G20), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT16), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n409), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n262), .B1(new_n404), .B2(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n321), .A2(new_n326), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n417), .B1(new_n326), .B2(new_n263), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n388), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT18), .ZN(new_n420));
  AND3_X1   g0220(.A1(new_n409), .A2(new_n413), .A3(new_n414), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n414), .B1(new_n409), .B2(new_n413), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n261), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n418), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n382), .A2(new_n384), .A3(new_n343), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(new_n387), .B2(G200), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n423), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT17), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n404), .A2(new_n415), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n418), .B1(new_n430), .B2(new_n261), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n431), .A2(KEYINPUT17), .A3(new_n426), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT18), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n433), .B(new_n388), .C1(new_n416), .C2(new_n418), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n420), .A2(new_n429), .A3(new_n432), .A4(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n372), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n249), .A2(G33), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n254), .A2(new_n262), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(G116), .ZN(new_n440));
  INV_X1    g0240(.A(G116), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n254), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n287), .A2(G97), .ZN(new_n444));
  NAND2_X1  g0244(.A1(G33), .A2(G283), .ZN(new_n445));
  AOI21_X1  g0245(.A(G20), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n225), .A2(new_n441), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n261), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT20), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n448), .A2(KEYINPUT83), .A3(new_n449), .ZN(new_n450));
  OAI211_X1 g0250(.A(KEYINPUT20), .B(new_n261), .C1(new_n446), .C2(new_n447), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(KEYINPUT83), .B1(new_n448), .B2(new_n449), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n443), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n249), .A2(G45), .ZN(new_n455));
  OR2_X1    g0255(.A1(KEYINPUT5), .A2(G41), .ZN(new_n456));
  NAND2_X1  g0256(.A1(KEYINPUT5), .A2(G41), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n455), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n458), .A2(new_n275), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n459), .A2(G270), .B1(G274), .B2(new_n458), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n294), .A2(G264), .A3(G1698), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n389), .A2(G303), .ZN(new_n462));
  OAI211_X1 g0262(.A(G257), .B(new_n285), .C1(new_n374), .C2(new_n375), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n275), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n460), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n466), .A2(KEYINPUT21), .A3(G169), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n460), .A2(new_n465), .A3(G179), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n303), .B1(new_n460), .B2(new_n465), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n454), .A2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT21), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n454), .A2(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n466), .A2(G190), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n474), .B1(new_n341), .B2(new_n466), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n473), .B1(new_n454), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n455), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G274), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n455), .A2(G250), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n275), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  OAI211_X1 g0281(.A(G244), .B(G1698), .C1(new_n374), .C2(new_n375), .ZN(new_n482));
  NAND2_X1  g0282(.A1(G33), .A2(G116), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT80), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n294), .A2(new_n485), .A3(G238), .A4(new_n285), .ZN(new_n486));
  OAI211_X1 g0286(.A(G238), .B(new_n285), .C1(new_n374), .C2(new_n375), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT80), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n484), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n318), .B(new_n481), .C1(new_n489), .C2(new_n276), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT81), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n488), .A2(new_n486), .ZN(new_n493));
  INV_X1    g0293(.A(new_n484), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n275), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n496), .A2(KEYINPUT81), .A3(new_n318), .A4(new_n481), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT77), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n439), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n254), .A2(KEYINPUT77), .A3(new_n262), .A4(new_n438), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n499), .A2(new_n348), .A3(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n254), .A2(new_n348), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT19), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n225), .B1(new_n292), .B2(new_n503), .ZN(new_n504));
  NOR4_X1   g0304(.A1(KEYINPUT82), .A2(G87), .A3(G97), .A4(G107), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT82), .ZN(new_n506));
  NOR2_X1   g0306(.A1(G87), .A2(G97), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n506), .B1(new_n507), .B2(new_n361), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n504), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n294), .A2(new_n225), .A3(G68), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n503), .B1(new_n292), .B2(G20), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n502), .B1(new_n512), .B2(new_n261), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n501), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n276), .B1(new_n493), .B2(new_n494), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n303), .B1(new_n515), .B2(new_n480), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n492), .A2(new_n497), .A3(new_n514), .A4(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(G200), .B1(new_n515), .B2(new_n480), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n499), .A2(G87), .A3(new_n500), .ZN(new_n519));
  OAI211_X1 g0319(.A(G190), .B(new_n481), .C1(new_n489), .C2(new_n276), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n518), .A2(new_n513), .A3(new_n519), .A4(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n476), .A2(new_n522), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n225), .B(G87), .C1(new_n374), .C2(new_n375), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT22), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT22), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n294), .A2(new_n526), .A3(new_n225), .A4(G87), .ZN(new_n527));
  AND2_X1   g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(KEYINPUT23), .B1(new_n225), .B2(G107), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT23), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n530), .A2(new_n361), .A3(G20), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n529), .B(new_n531), .C1(G20), .C2(new_n483), .ZN(new_n532));
  OAI211_X1 g0332(.A(KEYINPUT84), .B(KEYINPUT24), .C1(new_n528), .C2(new_n532), .ZN(new_n533));
  AOI211_X1 g0333(.A(KEYINPUT24), .B(new_n532), .C1(new_n525), .C2(new_n527), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT84), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n532), .B1(new_n525), .B2(new_n527), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT24), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n533), .A2(new_n535), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n261), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n321), .A2(new_n361), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT25), .ZN(new_n543));
  XNOR2_X1  g0343(.A(new_n542), .B(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n499), .A2(G107), .A3(new_n500), .ZN(new_n545));
  AND2_X1   g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n294), .A2(G257), .A3(G1698), .ZN(new_n548));
  NAND2_X1  g0348(.A1(G33), .A2(G294), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n548), .B(new_n549), .C1(new_n295), .C2(new_n214), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n275), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n458), .A2(G274), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n459), .A2(G264), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n554), .A2(G179), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n550), .A2(new_n275), .B1(G264), .B2(new_n459), .ZN(new_n556));
  AOI21_X1  g0356(.A(G169), .B1(new_n556), .B2(new_n552), .ZN(new_n557));
  NOR3_X1   g0357(.A1(new_n555), .A2(new_n557), .A3(KEYINPUT85), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT85), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n554), .A2(new_n303), .ZN(new_n560));
  INV_X1    g0360(.A(G179), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n556), .A2(new_n561), .A3(new_n552), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n559), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n547), .B1(new_n558), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n554), .A2(new_n341), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n556), .A2(new_n343), .A3(new_n552), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n541), .A2(new_n567), .A3(new_n546), .ZN(new_n568));
  AND2_X1   g0368(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n265), .A2(G77), .ZN(new_n570));
  OR2_X1    g0370(.A1(KEYINPUT76), .A2(KEYINPUT6), .ZN(new_n571));
  NAND2_X1  g0371(.A1(KEYINPUT76), .A2(KEYINPUT6), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n571), .B(new_n572), .C1(new_n215), .C2(G107), .ZN(new_n573));
  AND2_X1   g0373(.A1(new_n571), .A2(new_n572), .ZN(new_n574));
  XNOR2_X1  g0374(.A(G97), .B(G107), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n570), .B1(new_n576), .B2(new_n225), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n361), .B1(new_n407), .B2(new_n391), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n261), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n499), .A2(G97), .A3(new_n500), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n321), .A2(new_n215), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT79), .ZN(new_n583));
  INV_X1    g0383(.A(new_n445), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n584), .B1(new_n290), .B2(G250), .ZN(new_n585));
  OAI211_X1 g0385(.A(G244), .B(new_n285), .C1(new_n374), .C2(new_n375), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT78), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(KEYINPUT4), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n587), .A2(KEYINPUT4), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n585), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n589), .B1(new_n586), .B2(new_n588), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n275), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n459), .A2(G257), .B1(G274), .B2(new_n458), .ZN(new_n594));
  AND3_X1   g0394(.A1(new_n593), .A2(new_n385), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n303), .B1(new_n593), .B2(new_n594), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n582), .B(new_n583), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n593), .A2(new_n385), .A3(new_n594), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n456), .A2(new_n457), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n477), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n276), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n552), .B1(new_n602), .B2(new_n216), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n586), .A2(new_n588), .ZN(new_n604));
  INV_X1    g0404(.A(new_n589), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n606), .A2(new_n590), .A3(new_n585), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n603), .B1(new_n607), .B2(new_n275), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n599), .B1(new_n303), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n583), .B1(new_n609), .B2(new_n582), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n598), .A2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n582), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n608), .A2(new_n343), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n608), .A2(G200), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n612), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n523), .A2(new_n569), .A3(new_n611), .A4(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n437), .A2(new_n616), .ZN(G372));
  NAND2_X1  g0417(.A1(new_n423), .A2(new_n424), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n433), .B1(new_n618), .B2(new_n388), .ZN(new_n619));
  INV_X1    g0419(.A(new_n434), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n367), .ZN(new_n622));
  INV_X1    g0422(.A(new_n301), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n300), .B1(new_n284), .B2(new_n297), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n304), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n625), .B1(KEYINPUT73), .B2(KEYINPUT14), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n626), .A2(new_n306), .A3(new_n307), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n622), .B1(new_n627), .B2(new_n274), .ZN(new_n628));
  AOI21_X1  g0428(.A(KEYINPUT17), .B1(new_n431), .B2(new_n426), .ZN(new_n629));
  AND4_X1   g0429(.A1(KEYINPUT17), .A2(new_n423), .A3(new_n424), .A4(new_n426), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n346), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n621), .B1(new_n628), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n338), .A2(new_n339), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n331), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n514), .A2(new_n516), .A3(new_n490), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n609), .A2(new_n521), .A3(new_n636), .A4(new_n582), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n636), .B1(new_n637), .B2(KEYINPUT26), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n517), .B(new_n521), .C1(new_n598), .C2(new_n610), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n638), .B1(new_n639), .B2(KEYINPUT26), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n521), .A2(new_n636), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n555), .A2(new_n557), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n537), .A2(new_n538), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n534), .B1(new_n643), .B2(KEYINPUT84), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n262), .B1(new_n644), .B2(new_n539), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n499), .A2(new_n500), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n544), .B1(new_n646), .B2(new_n361), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n642), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n641), .B1(new_n648), .B2(new_n473), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n649), .A2(new_n611), .A3(new_n615), .A4(new_n568), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n640), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n635), .B1(new_n437), .B2(new_n652), .ZN(G369));
  NAND3_X1  g0453(.A1(new_n249), .A2(new_n225), .A3(G13), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n655), .A2(G213), .A3(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(G343), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n547), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n564), .A2(new_n568), .A3(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(KEYINPUT85), .B1(new_n555), .B2(new_n557), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n560), .A2(new_n559), .A3(new_n562), .ZN(new_n663));
  AOI22_X1  g0463(.A1(new_n662), .A2(new_n663), .B1(new_n541), .B2(new_n546), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n659), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n454), .A2(new_n659), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n476), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n473), .A2(new_n454), .A3(new_n659), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n669), .A2(G330), .A3(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n473), .A2(new_n659), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n674), .A2(new_n564), .A3(new_n568), .A4(new_n660), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n560), .A2(new_n562), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n676), .B1(new_n541), .B2(new_n546), .ZN(new_n677));
  INV_X1    g0477(.A(new_n659), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n673), .A2(new_n680), .ZN(G399));
  INV_X1    g0481(.A(new_n228), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(G41), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n223), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n683), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(G1), .ZN(new_n686));
  OR3_X1    g0486(.A1(new_n505), .A2(new_n508), .A3(G116), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n684), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT28), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n554), .A2(new_n318), .A3(new_n466), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n515), .A2(new_n480), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT30), .ZN(new_n693));
  INV_X1    g0493(.A(new_n468), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n694), .A2(new_n608), .A3(new_n691), .A4(new_n556), .ZN(new_n695));
  OAI22_X1  g0495(.A1(new_n692), .A2(new_n608), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n695), .A2(new_n693), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n659), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n698), .A2(KEYINPUT31), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n616), .B2(new_n659), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n698), .A2(KEYINPUT31), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(G330), .A3(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n641), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n469), .A2(new_n454), .ZN(new_n704));
  INV_X1    g0504(.A(new_n471), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n704), .B1(new_n705), .B2(KEYINPUT21), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n703), .B1(new_n664), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n582), .B1(new_n595), .B2(new_n596), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(KEYINPUT79), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n709), .A2(new_n568), .A3(new_n615), .A4(new_n597), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n636), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n712), .B1(new_n637), .B2(KEYINPUT26), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n639), .B2(KEYINPUT26), .ZN(new_n714));
  OAI211_X1 g0514(.A(KEYINPUT29), .B(new_n678), .C1(new_n711), .C2(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n659), .B1(new_n640), .B2(new_n650), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n715), .B1(KEYINPUT29), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n702), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n689), .B1(new_n719), .B2(G1), .ZN(G364));
  INV_X1    g0520(.A(new_n671), .ZN(new_n721));
  INV_X1    g0521(.A(G13), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(G20), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n686), .B1(G45), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(G330), .B1(new_n669), .B2(new_n670), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n669), .A2(new_n670), .ZN(new_n728));
  NOR2_X1   g0528(.A1(G13), .A2(G33), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(G20), .ZN(new_n731));
  AND2_X1   g0531(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n224), .B1(G20), .B2(new_n303), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n225), .A2(G190), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n385), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(new_n341), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR4_X1   g0538(.A1(new_n318), .A2(new_n225), .A3(new_n343), .A4(new_n341), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  OAI22_X1  g0540(.A1(new_n738), .A2(new_n203), .B1(new_n207), .B2(new_n740), .ZN(new_n741));
  NOR4_X1   g0541(.A1(new_n318), .A2(new_n225), .A3(new_n343), .A4(G200), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n741), .B1(G58), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G179), .A2(G200), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n735), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g0545(.A(KEYINPUT89), .B(KEYINPUT32), .ZN(new_n746));
  OR3_X1    g0546(.A1(new_n745), .A2(new_n746), .A3(new_n394), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n744), .A2(G190), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G20), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G97), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n746), .B1(new_n745), .B2(new_n394), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n747), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n341), .A2(G179), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n753), .A2(G20), .A3(G190), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G87), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n735), .A2(new_n753), .ZN(new_n757));
  OAI211_X1 g0557(.A(new_n756), .B(new_n294), .C1(new_n361), .C2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n736), .A2(G200), .ZN(new_n759));
  AOI211_X1 g0559(.A(new_n752), .B(new_n758), .C1(G77), .C2(new_n759), .ZN(new_n760));
  AOI22_X1  g0560(.A1(G322), .A2(new_n742), .B1(new_n739), .B2(G326), .ZN(new_n761));
  XNOR2_X1  g0561(.A(KEYINPUT33), .B(G317), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n737), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n759), .A2(G311), .ZN(new_n764));
  AND3_X1   g0564(.A1(new_n761), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n745), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n755), .A2(G303), .B1(new_n766), .B2(G329), .ZN(new_n767));
  INV_X1    g0567(.A(G283), .ZN(new_n768));
  OAI211_X1 g0568(.A(new_n767), .B(new_n389), .C1(new_n768), .C2(new_n757), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n769), .B1(G294), .B2(new_n749), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n743), .A2(new_n760), .B1(new_n765), .B2(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n734), .B1(new_n771), .B2(KEYINPUT90), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(KEYINPUT90), .B2(new_n771), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n682), .A2(new_n389), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n774), .A2(G355), .B1(new_n441), .B2(new_n682), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n389), .A2(new_n228), .ZN(new_n776));
  XOR2_X1   g0576(.A(new_n776), .B(KEYINPUT87), .Z(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n223), .A2(G45), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n779), .B1(new_n247), .B2(G45), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n775), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n731), .A2(new_n733), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n782), .B(KEYINPUT88), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  XOR2_X1   g0584(.A(new_n724), .B(KEYINPUT86), .Z(new_n785));
  NAND3_X1  g0585(.A1(new_n773), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n726), .A2(new_n727), .B1(new_n732), .B2(new_n786), .ZN(G396));
  AND3_X1   g0587(.A1(new_n358), .A2(new_n366), .A3(new_n678), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n358), .A2(new_n659), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(new_n370), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n788), .B1(new_n790), .B2(new_n367), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n716), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n641), .A2(new_n708), .ZN(new_n793));
  INV_X1    g0593(.A(KEYINPUT26), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n712), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n522), .B1(new_n709), .B2(new_n597), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n795), .B1(new_n796), .B2(new_n794), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n703), .B1(new_n706), .B2(new_n677), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n710), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n678), .B(new_n791), .C1(new_n797), .C2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(KEYINPUT95), .ZN(new_n801));
  INV_X1    g0601(.A(KEYINPUT95), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n651), .A2(new_n802), .A3(new_n678), .A4(new_n791), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n792), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n702), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OR2_X1    g0606(.A1(new_n806), .A2(KEYINPUT96), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(KEYINPUT96), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n724), .B1(new_n804), .B2(new_n805), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n807), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n733), .A2(new_n729), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n759), .ZN(new_n813));
  XNOR2_X1  g0613(.A(KEYINPUT91), .B(G283), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n441), .A2(new_n813), .B1(new_n738), .B2(new_n814), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n755), .A2(G107), .B1(new_n766), .B2(G311), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n757), .A2(new_n213), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(new_n294), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n816), .A2(new_n818), .A3(new_n750), .ZN(new_n819));
  INV_X1    g0619(.A(G294), .ZN(new_n820));
  INV_X1    g0620(.A(new_n742), .ZN(new_n821));
  INV_X1    g0621(.A(G303), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n820), .A2(new_n821), .B1(new_n740), .B2(new_n822), .ZN(new_n823));
  NOR3_X1   g0623(.A1(new_n815), .A2(new_n819), .A3(new_n823), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n754), .A2(new_n207), .B1(new_n757), .B2(new_n203), .ZN(new_n825));
  INV_X1    g0625(.A(G132), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n294), .B1(new_n745), .B2(new_n826), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT92), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n825), .B(new_n828), .C1(G58), .C2(new_n749), .ZN(new_n829));
  XOR2_X1   g0629(.A(new_n829), .B(KEYINPUT93), .Z(new_n830));
  AOI22_X1  g0630(.A1(new_n759), .A2(G159), .B1(G137), .B2(new_n739), .ZN(new_n831));
  INV_X1    g0631(.A(G143), .ZN(new_n832));
  INV_X1    g0632(.A(G150), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n831), .B1(new_n832), .B2(new_n821), .C1(new_n833), .C2(new_n738), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n834), .B(KEYINPUT34), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n824), .B1(new_n830), .B2(new_n835), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n785), .B1(G77), .B2(new_n812), .C1(new_n836), .C2(new_n734), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT94), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n730), .B2(new_n791), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n810), .A2(new_n839), .ZN(G384));
  NAND2_X1  g0640(.A1(G50), .A2(G77), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n399), .A2(new_n841), .B1(G50), .B2(new_n203), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n842), .A2(G1), .A3(new_n722), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT35), .ZN(new_n844));
  OR2_X1    g0644(.A1(new_n576), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n576), .A2(new_n844), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n845), .A2(G116), .A3(new_n226), .A4(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT36), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n843), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(new_n848), .B2(new_n847), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT38), .ZN(new_n851));
  XOR2_X1   g0651(.A(new_n657), .B(KEYINPUT98), .Z(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n416), .B2(new_n418), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(new_n621), .B2(new_n631), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT97), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n419), .A2(new_n855), .ZN(new_n856));
  OAI211_X1 g0656(.A(KEYINPUT97), .B(new_n388), .C1(new_n416), .C2(new_n418), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT37), .ZN(new_n859));
  AND3_X1   g0659(.A1(new_n853), .A2(new_n427), .A3(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n419), .A2(new_n853), .A3(new_n427), .ZN(new_n861));
  AOI22_X1  g0661(.A1(new_n858), .A2(new_n860), .B1(KEYINPUT37), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n851), .B1(new_n854), .B2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n657), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n864), .B1(new_n416), .B2(new_n418), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n419), .A2(new_n865), .A3(new_n427), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(KEYINPUT37), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT97), .B1(new_n618), .B2(new_n388), .ZN(new_n868));
  INV_X1    g0668(.A(new_n857), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n853), .A2(new_n427), .A3(new_n859), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n867), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n435), .A2(new_n618), .A3(new_n864), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n872), .A2(new_n873), .A3(KEYINPUT38), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n863), .A2(new_n874), .ZN(new_n875));
  OR2_X1    g0675(.A1(new_n875), .A2(KEYINPUT99), .ZN(new_n876));
  INV_X1    g0676(.A(new_n791), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n274), .A2(new_n659), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n310), .A2(new_n346), .A3(new_n878), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n274), .B(new_n659), .C1(new_n627), .C2(new_n345), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n877), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AND3_X1   g0681(.A1(new_n881), .A2(new_n700), .A3(new_n701), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n875), .A2(KEYINPUT99), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n876), .A2(new_n882), .A3(KEYINPUT40), .A4(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT40), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n881), .A2(new_n700), .A3(new_n701), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n865), .B1(new_n621), .B2(new_n631), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n858), .A2(new_n860), .B1(KEYINPUT37), .B2(new_n866), .ZN(new_n888));
  NOR3_X1   g0688(.A1(new_n887), .A2(new_n888), .A3(new_n851), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT38), .B1(new_n872), .B2(new_n873), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n885), .B1(new_n886), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n884), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n893), .B(KEYINPUT100), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n436), .A2(new_n700), .A3(new_n701), .ZN(new_n895));
  OR2_X1    g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n894), .A2(new_n895), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n896), .A2(G330), .A3(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n621), .A2(new_n852), .ZN(new_n899));
  OAI21_X1  g0699(.A(KEYINPUT39), .B1(new_n889), .B2(new_n890), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT39), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n863), .A2(new_n901), .A3(new_n874), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n627), .A2(new_n274), .A3(new_n678), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n899), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n788), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n800), .A2(KEYINPUT95), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n802), .B1(new_n716), .B2(new_n791), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n891), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n879), .A2(new_n880), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n906), .A2(new_n913), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n436), .B(new_n715), .C1(KEYINPUT29), .C2(new_n716), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n635), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n914), .B(new_n916), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n898), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(KEYINPUT101), .ZN(new_n919));
  OAI221_X1 g0719(.A(new_n919), .B1(new_n249), .B2(new_n723), .C1(new_n898), .C2(new_n917), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n918), .A2(KEYINPUT101), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n850), .B1(new_n920), .B2(new_n921), .ZN(G367));
  NAND2_X1  g0722(.A1(new_n582), .A2(new_n659), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n709), .A2(new_n597), .A3(new_n615), .A4(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n609), .A2(new_n582), .A3(new_n659), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n611), .B1(new_n926), .B2(new_n564), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n678), .ZN(new_n928));
  OAI21_X1  g0728(.A(KEYINPUT42), .B1(new_n926), .B2(new_n675), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n519), .A2(new_n513), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n659), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n641), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n636), .A2(new_n930), .A3(new_n659), .ZN(new_n933));
  AOI21_X1  g0733(.A(KEYINPUT43), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n675), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n924), .A2(new_n925), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT42), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n928), .A2(new_n929), .A3(new_n934), .A4(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(KEYINPUT102), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n938), .A2(new_n929), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT102), .ZN(new_n942));
  NAND4_X1  g0742(.A1(new_n941), .A2(new_n942), .A3(new_n934), .A4(new_n928), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT103), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n940), .A2(new_n943), .A3(KEYINPUT103), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n941), .A2(new_n928), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n932), .A2(new_n933), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT43), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n946), .A2(new_n947), .A3(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n673), .A2(new_n926), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n944), .A2(new_n945), .B1(new_n948), .B2(new_n950), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n956), .A2(new_n953), .A3(new_n947), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n683), .B(KEYINPUT41), .Z(new_n958));
  OAI22_X1  g0758(.A1(new_n680), .A2(new_n936), .B1(KEYINPUT104), .B2(KEYINPUT44), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n675), .A2(new_n679), .ZN(new_n960));
  NOR2_X1   g0760(.A1(KEYINPUT104), .A2(KEYINPUT44), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n960), .A2(new_n926), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(KEYINPUT104), .A2(KEYINPUT44), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(KEYINPUT45), .B1(new_n680), .B2(new_n936), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT45), .ZN(new_n967));
  NOR3_X1   g0767(.A1(new_n960), .A2(new_n967), .A3(new_n926), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n965), .A2(new_n970), .A3(new_n673), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n675), .B1(new_n666), .B2(new_n674), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n721), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n671), .B(new_n675), .C1(new_n666), .C2(new_n674), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n702), .A2(new_n717), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(KEYINPUT105), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n959), .A2(new_n962), .B1(KEYINPUT104), .B2(KEYINPUT44), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n672), .B1(new_n978), .B2(new_n969), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT105), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n702), .A2(new_n717), .A3(new_n975), .A4(new_n980), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n971), .A2(new_n977), .A3(new_n979), .A4(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n958), .B1(new_n982), .B2(new_n719), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n723), .A2(G45), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(G1), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n955), .B(new_n957), .C1(new_n983), .C2(new_n985), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n755), .A2(G58), .B1(new_n766), .B2(G137), .ZN(new_n987));
  INV_X1    g0787(.A(new_n749), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n987), .B1(new_n203), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n294), .B1(new_n757), .B2(new_n269), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n740), .A2(new_n832), .B1(KEYINPUT106), .B2(new_n990), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n989), .B(new_n991), .C1(KEYINPUT106), .C2(new_n990), .ZN(new_n992));
  AOI22_X1  g0792(.A1(G50), .A2(new_n759), .B1(new_n737), .B2(G159), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n992), .B(new_n993), .C1(new_n833), .C2(new_n821), .ZN(new_n994));
  INV_X1    g0794(.A(G317), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n389), .B1(new_n745), .B2(new_n995), .C1(new_n215), .C2(new_n757), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n755), .A2(KEYINPUT46), .A3(G116), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT46), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n754), .B2(new_n441), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n997), .B(new_n999), .C1(new_n361), .C2(new_n988), .ZN(new_n1000));
  AOI211_X1 g0800(.A(new_n996), .B(new_n1000), .C1(G294), .C2(new_n737), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n814), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n759), .A2(new_n1002), .B1(G311), .B2(new_n739), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n1001), .B(new_n1003), .C1(new_n822), .C2(new_n821), .ZN(new_n1004));
  AND2_X1   g0804(.A1(new_n994), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n734), .B1(new_n1005), .B2(KEYINPUT47), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(KEYINPUT47), .B2(new_n1005), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n782), .B1(new_n228), .B2(new_n349), .C1(new_n778), .C2(new_n239), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1007), .A2(new_n785), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(new_n731), .B2(new_n949), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n986), .A2(new_n1011), .ZN(G387));
  NAND2_X1  g0812(.A1(new_n326), .A2(new_n207), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT50), .ZN(new_n1014));
  INV_X1    g0814(.A(G45), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n203), .B2(new_n269), .ZN(new_n1016));
  NOR3_X1   g0816(.A1(new_n1014), .A2(new_n687), .A3(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n777), .B1(new_n236), .B2(new_n1015), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n687), .A2(new_n774), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1017), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n228), .A2(G107), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n783), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(new_n785), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n755), .A2(G294), .B1(new_n1002), .B2(new_n749), .ZN(new_n1024));
  XOR2_X1   g0824(.A(KEYINPUT108), .B(G322), .Z(new_n1025));
  AOI22_X1  g0825(.A1(new_n737), .A2(G311), .B1(new_n739), .B2(new_n1025), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1026), .B1(new_n822), .B2(new_n813), .C1(new_n995), .C2(new_n821), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT48), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1024), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(new_n1028), .B2(new_n1027), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(KEYINPUT109), .B(KEYINPUT49), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n389), .B1(new_n757), .B2(new_n441), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(G326), .B2(new_n766), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1032), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n813), .A2(new_n203), .B1(new_n207), .B2(new_n821), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(new_n326), .B2(new_n737), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n739), .A2(G159), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT107), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n988), .A2(new_n349), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n294), .B1(new_n757), .B2(new_n215), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n754), .A2(new_n269), .B1(new_n745), .B2(new_n833), .ZN(new_n1043));
  NOR3_X1   g0843(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1038), .A2(new_n1040), .A3(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n734), .B1(new_n1036), .B2(new_n1045), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n1023), .B(new_n1046), .C1(new_n667), .C2(new_n731), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(new_n975), .B2(new_n985), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n975), .ZN(new_n1049));
  AND3_X1   g0849(.A1(new_n718), .A2(new_n1049), .A3(KEYINPUT111), .ZN(new_n1050));
  AOI21_X1  g0850(.A(KEYINPUT111), .B1(new_n718), .B2(new_n1049), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n685), .B1(new_n977), .B2(new_n981), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT110), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1052), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1048), .B1(new_n1055), .B2(new_n1056), .ZN(G393));
  NAND3_X1  g0857(.A1(new_n971), .A2(new_n979), .A3(new_n985), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n244), .A2(new_n778), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n782), .B1(new_n215), .B2(new_n228), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n785), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n755), .A2(new_n1002), .B1(new_n766), .B2(new_n1025), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1062), .B(new_n389), .C1(new_n361), .C2(new_n757), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT113), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n737), .A2(G303), .B1(G116), .B2(new_n749), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1064), .B(new_n1065), .C1(new_n820), .C2(new_n813), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(G311), .A2(new_n742), .B1(new_n739), .B2(G317), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT52), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(G150), .A2(new_n739), .B1(new_n742), .B2(G159), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT51), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G50), .A2(new_n737), .B1(new_n759), .B2(new_n326), .ZN(new_n1071));
  OR2_X1    g0871(.A1(new_n1071), .A2(KEYINPUT112), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1071), .A2(KEYINPUT112), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n988), .A2(new_n269), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n754), .A2(new_n203), .B1(new_n745), .B2(new_n832), .ZN(new_n1075));
  NOR4_X1   g0875(.A1(new_n1074), .A2(new_n1075), .A3(new_n389), .A4(new_n817), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1072), .A2(new_n1073), .A3(new_n1076), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n1066), .A2(new_n1068), .B1(new_n1070), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1061), .B1(new_n1078), .B2(new_n733), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n731), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1079), .B1(new_n936), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1058), .A2(new_n1081), .ZN(new_n1082));
  AND2_X1   g0882(.A1(new_n982), .A2(new_n683), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n971), .A2(new_n979), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n977), .A2(new_n981), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1082), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(G390));
  AOI21_X1  g0888(.A(new_n788), .B1(new_n801), .B2(new_n803), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n912), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n904), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  AND3_X1   g0891(.A1(new_n863), .A2(new_n901), .A3(new_n874), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n851), .B1(new_n887), .B2(new_n888), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n901), .B1(new_n1093), .B2(new_n874), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1091), .A2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n678), .B1(new_n711), .B2(new_n714), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n790), .A2(new_n367), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n907), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n912), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n876), .A2(new_n883), .A3(new_n1101), .A4(new_n904), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1096), .A2(new_n1102), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n881), .A2(new_n700), .A3(G330), .A4(new_n701), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1096), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n700), .A2(G330), .A3(new_n701), .A4(new_n791), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n1090), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n1104), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n1089), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n436), .A2(new_n700), .A3(G330), .A4(new_n701), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n915), .A2(new_n1113), .A3(new_n635), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1110), .A2(new_n1100), .A3(new_n1104), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1112), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n685), .B1(new_n1108), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1117), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1106), .A2(new_n1119), .A3(new_n1107), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n985), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1108), .A2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n903), .A2(new_n730), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(G116), .A2(new_n742), .B1(new_n739), .B2(G283), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n1125), .B1(new_n738), .B2(new_n361), .C1(new_n215), .C2(new_n813), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1074), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n757), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(G68), .A2(new_n1128), .B1(new_n766), .B2(G294), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1127), .A2(new_n389), .A3(new_n756), .A4(new_n1129), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n737), .A2(G137), .B1(G132), .B2(new_n742), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n757), .A2(new_n207), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n389), .B(new_n1132), .C1(G125), .C2(new_n766), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1131), .B(new_n1133), .C1(new_n394), .C2(new_n988), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n754), .A2(new_n833), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1135), .B(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n739), .A2(G128), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(KEYINPUT54), .B(G143), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1137), .B(new_n1138), .C1(new_n813), .C2(new_n1139), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n1126), .A2(new_n1130), .B1(new_n1134), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n733), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1142), .B(new_n785), .C1(new_n326), .C2(new_n812), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1124), .A2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1123), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1121), .A2(new_n1145), .ZN(G378));
  AND3_X1   g0946(.A1(new_n884), .A2(G330), .A3(new_n892), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n330), .A2(new_n657), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(new_n340), .B(new_n1148), .ZN(new_n1149));
  XOR2_X1   g0949(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1150));
  XNOR2_X1  g0950(.A(new_n1149), .B(new_n1150), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n906), .A2(new_n913), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1151), .B1(new_n906), .B2(new_n913), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1147), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1151), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n1095), .A2(new_n904), .B1(new_n621), .B2(new_n852), .ZN(new_n1156));
  NOR3_X1   g0956(.A1(new_n1089), .A2(new_n891), .A3(new_n1090), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1155), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n884), .A2(G330), .A3(new_n892), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n906), .A2(new_n913), .A3(new_n1151), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1154), .A2(new_n1161), .ZN(new_n1162));
  AND3_X1   g0962(.A1(new_n1096), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1104), .B1(new_n1096), .B2(new_n1102), .ZN(new_n1164));
  NOR3_X1   g0964(.A1(new_n1163), .A2(new_n1164), .A3(new_n1117), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1162), .B(KEYINPUT57), .C1(new_n1165), .C2(new_n1114), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(KEYINPUT116), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1162), .B1(new_n1165), .B2(new_n1114), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT57), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1120), .A2(new_n1115), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT116), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1171), .A2(new_n1172), .A3(KEYINPUT57), .A4(new_n1162), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1167), .A2(new_n1170), .A3(new_n683), .A4(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n724), .B1(G50), .B2(new_n812), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1155), .A2(new_n730), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n988), .A2(new_n833), .B1(new_n1139), .B2(new_n754), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n759), .A2(G137), .B1(G128), .B2(new_n742), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n826), .B2(new_n738), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n1177), .B(new_n1179), .C1(G125), .C2(new_n739), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT59), .ZN(new_n1181));
  OR2_X1    g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(G33), .A2(G41), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n757), .B2(new_n394), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(G124), .B2(new_n766), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1182), .A2(new_n1183), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(G41), .ZN(new_n1188));
  AOI211_X1 g0988(.A(G50), .B(new_n1184), .C1(new_n389), .C2(new_n1188), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1188), .B(new_n389), .C1(new_n745), .C2(new_n768), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n754), .A2(new_n269), .B1(new_n757), .B2(new_n202), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n1190), .B(new_n1191), .C1(G68), .C2(new_n749), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n759), .A2(new_n348), .B1(G116), .B2(new_n739), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n737), .A2(G97), .B1(G107), .B2(new_n742), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT58), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1189), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1187), .B(new_n1197), .C1(new_n1196), .C2(new_n1195), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n1175), .B(new_n1176), .C1(new_n733), .C2(new_n1198), .ZN(new_n1199));
  OR2_X1    g0999(.A1(new_n1199), .A2(KEYINPUT115), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(KEYINPUT115), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1200), .A2(new_n1201), .B1(new_n985), .B2(new_n1162), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1174), .A2(new_n1202), .ZN(G375));
  NAND3_X1  g1003(.A1(new_n1112), .A2(new_n985), .A3(new_n1116), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n785), .B1(G68), .B2(new_n812), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n755), .A2(G159), .B1(new_n766), .B2(G128), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1206), .B1(new_n207), .B2(new_n988), .C1(new_n738), .C2(new_n1139), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n389), .B1(new_n1128), .B2(G58), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n813), .A2(new_n833), .B1(new_n1209), .B2(KEYINPUT118), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1207), .A2(new_n1210), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n1209), .A2(KEYINPUT118), .B1(G137), .B2(new_n742), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1211), .B(new_n1212), .C1(new_n826), .C2(new_n740), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n759), .A2(G107), .B1(G294), .B2(new_n739), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n441), .B2(new_n738), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1215), .B(KEYINPUT117), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n755), .A2(G97), .B1(new_n766), .B2(G303), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1217), .B(new_n389), .C1(new_n269), .C2(new_n757), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1218), .A2(new_n1041), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1219), .B1(new_n768), .B2(new_n821), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1213), .B1(new_n1216), .B2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1205), .B1(new_n1221), .B2(new_n733), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n912), .B2(new_n730), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1204), .A2(new_n1223), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1119), .A2(new_n958), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1112), .A2(new_n1116), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(new_n1114), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1224), .B1(new_n1225), .B2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(G381));
  INV_X1    g1029(.A(G378), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1174), .A2(new_n1230), .A3(new_n1202), .ZN(new_n1231));
  INV_X1    g1031(.A(G396), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1232), .B(new_n1048), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1233));
  INV_X1    g1033(.A(G384), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1228), .A2(new_n1234), .A3(new_n1087), .ZN(new_n1235));
  OR4_X1    g1035(.A1(G387), .A2(new_n1231), .A3(new_n1233), .A4(new_n1235), .ZN(G407));
  OAI211_X1 g1036(.A(G407), .B(G213), .C1(G343), .C2(new_n1231), .ZN(G409));
  NAND2_X1  g1037(.A1(G393), .A2(G396), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n1238), .A2(KEYINPUT123), .A3(new_n1233), .ZN(new_n1239));
  AOI21_X1  g1039(.A(KEYINPUT123), .B1(new_n1238), .B2(new_n1233), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(G387), .A2(new_n1087), .ZN(new_n1242));
  OR2_X1    g1042(.A1(new_n983), .A2(new_n985), .ZN(new_n1243));
  AND2_X1   g1043(.A1(new_n955), .A2(new_n957), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1010), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1245), .A2(G390), .ZN(new_n1246));
  OR3_X1    g1046(.A1(new_n1241), .A2(new_n1242), .A3(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1245), .A2(KEYINPUT124), .A3(G390), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT124), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(G387), .B2(new_n1087), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1248), .B1(new_n1250), .B2(new_n1242), .ZN(new_n1251));
  AND3_X1   g1051(.A1(new_n1251), .A2(new_n1241), .A3(KEYINPUT125), .ZN(new_n1252));
  AOI21_X1  g1052(.A(KEYINPUT125), .B1(new_n1251), .B2(new_n1241), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1247), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1254), .A2(KEYINPUT127), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT127), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1251), .A2(new_n1241), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT125), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1251), .A2(new_n1241), .A3(KEYINPUT125), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1256), .B1(new_n1261), .B2(new_n1247), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1255), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT61), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n658), .A2(G213), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1174), .A2(G378), .A3(new_n1202), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1199), .B1(new_n1162), .B2(new_n985), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1268), .B1(new_n1168), .B2(new_n958), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1230), .A2(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1266), .B1(new_n1267), .B2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1266), .A2(G2897), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT60), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1226), .A2(new_n1274), .A3(new_n1114), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1274), .B1(new_n1226), .B2(new_n1114), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n683), .B(new_n1117), .C1(new_n1276), .C2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1224), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1278), .A2(G384), .A3(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(G384), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1280), .B1(new_n1281), .B2(KEYINPUT119), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1117), .A2(new_n683), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1277), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1283), .B1(new_n1284), .B2(new_n1275), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1234), .B1(new_n1285), .B2(new_n1224), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT119), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1273), .B1(new_n1282), .B2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1281), .A2(KEYINPUT119), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1290), .A2(new_n1291), .A3(new_n1280), .A4(new_n1272), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1289), .A2(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1264), .B1(new_n1271), .B2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(KEYINPUT126), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT126), .ZN(new_n1296));
  OAI211_X1 g1096(.A(new_n1296), .B(new_n1264), .C1(new_n1271), .C2(new_n1293), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1282), .A2(new_n1288), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1271), .A2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(KEYINPUT62), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1295), .A2(new_n1297), .A3(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT120), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1299), .A2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1271), .A2(KEYINPUT120), .A3(new_n1298), .ZN(new_n1304));
  AOI21_X1  g1104(.A(KEYINPUT62), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1263), .B1(new_n1301), .B2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1271), .A2(KEYINPUT121), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1293), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1271), .A2(KEYINPUT121), .ZN(new_n1310));
  OAI21_X1  g1110(.A(KEYINPUT122), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT63), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1303), .A2(new_n1312), .A3(new_n1304), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1293), .B1(new_n1271), .B2(KEYINPUT121), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT122), .ZN(new_n1315));
  OAI211_X1 g1115(.A(new_n1314), .B(new_n1315), .C1(KEYINPUT121), .C2(new_n1271), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1271), .A2(KEYINPUT63), .A3(new_n1298), .ZN(new_n1317));
  AND3_X1   g1117(.A1(new_n1317), .A2(new_n1264), .A3(new_n1254), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1311), .A2(new_n1313), .A3(new_n1316), .A4(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1306), .A2(new_n1319), .ZN(G405));
  INV_X1    g1120(.A(new_n1298), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1254), .A2(KEYINPUT127), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1261), .A2(new_n1256), .A3(new_n1247), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(G375), .A2(G378), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(new_n1231), .ZN(new_n1325));
  AND3_X1   g1125(.A1(new_n1322), .A2(new_n1323), .A3(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1325), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1321), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1325), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1329), .B1(new_n1255), .B2(new_n1262), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1322), .A2(new_n1323), .A3(new_n1325), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1330), .A2(new_n1298), .A3(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1328), .A2(new_n1332), .ZN(G402));
endmodule


