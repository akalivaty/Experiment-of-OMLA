//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 0 0 1 0 1 0 0 1 0 1 0 1 0 0 1 1 0 0 0 1 1 0 1 1 0 0 1 1 0 1 1 0 0 0 1 1 1 0 1 0 1 0 1 0 0 1 0 1 0 0 1 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:17 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n548, new_n549, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n558, new_n559, new_n560, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n569, new_n570, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n583, new_n584, new_n585, new_n588, new_n590, new_n591,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT66), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  XOR2_X1   g031(.A(G325), .B(KEYINPUT67), .Z(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(KEYINPUT68), .B1(new_n462), .B2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n464), .A2(new_n465), .A3(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n468));
  NAND4_X1  g043(.A1(new_n463), .A2(new_n466), .A3(new_n467), .A4(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G137), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n465), .A2(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(new_n468), .A3(G125), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n467), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AND3_X1   g050(.A1(new_n467), .A2(G101), .A3(G2104), .ZN(new_n476));
  NOR3_X1   g051(.A1(new_n471), .A2(new_n475), .A3(new_n476), .ZN(G160));
  INV_X1    g052(.A(G136), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n467), .A2(G112), .ZN(new_n479));
  OAI21_X1  g054(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n480));
  OAI22_X1  g055(.A1(new_n469), .A2(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AND2_X1   g056(.A1(new_n466), .A2(new_n468), .ZN(new_n482));
  NAND4_X1  g057(.A1(new_n482), .A2(KEYINPUT69), .A3(G2105), .A4(new_n463), .ZN(new_n483));
  NAND4_X1  g058(.A1(new_n463), .A2(new_n466), .A3(G2105), .A4(new_n468), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT69), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n481), .B1(new_n487), .B2(G124), .ZN(G162));
  NAND2_X1  g063(.A1(KEYINPUT4), .A2(G138), .ZN(new_n489));
  OR2_X1    g064(.A1(new_n469), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n472), .A2(new_n468), .A3(G138), .A4(new_n467), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  AND2_X1   g067(.A1(KEYINPUT71), .A2(G114), .ZN(new_n493));
  NOR2_X1   g068(.A1(KEYINPUT71), .A2(G114), .ZN(new_n494));
  OAI21_X1  g069(.A(G2105), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  AOI22_X1  g072(.A1(new_n491), .A2(new_n492), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  AND2_X1   g073(.A1(G126), .A2(G2105), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n463), .A2(new_n466), .A3(new_n468), .A4(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n501));
  AND2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n500), .A2(new_n501), .ZN(new_n503));
  OAI211_X1 g078(.A(new_n490), .B(new_n498), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  OR2_X1    g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G50), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n507), .A2(new_n508), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT5), .B(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n510), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OR2_X1    g093(.A1(new_n515), .A2(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  NAND3_X1  g095(.A1(new_n512), .A2(G63), .A3(G651), .ZN(new_n521));
  XOR2_X1   g096(.A(new_n521), .B(KEYINPUT72), .Z(new_n522));
  AOI21_X1  g097(.A(new_n522), .B1(G51), .B2(new_n509), .ZN(new_n523));
  INV_X1    g098(.A(new_n513), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n524), .A2(G89), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT73), .B(KEYINPUT7), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n526), .B(new_n527), .ZN(new_n528));
  OAI21_X1  g103(.A(KEYINPUT74), .B1(new_n525), .B2(new_n528), .ZN(new_n529));
  OR3_X1    g104(.A1(new_n525), .A2(KEYINPUT74), .A3(new_n528), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n523), .A2(new_n529), .A3(new_n530), .ZN(G286));
  INV_X1    g106(.A(G286), .ZN(G168));
  NAND2_X1  g107(.A1(new_n509), .A2(G52), .ZN(new_n533));
  INV_X1    g108(.A(G90), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n533), .B1(new_n513), .B2(new_n534), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n536), .A2(new_n517), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n535), .A2(new_n537), .ZN(G171));
  XOR2_X1   g113(.A(KEYINPUT75), .B(G81), .Z(new_n539));
  NAND2_X1  g114(.A1(new_n524), .A2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(G43), .ZN(new_n541));
  INV_X1    g116(.A(new_n509), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  OAI221_X1 g118(.A(new_n540), .B1(new_n541), .B2(new_n542), .C1(new_n517), .C2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  NAND4_X1  g121(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND4_X1  g124(.A1(G319), .A2(G483), .A3(G661), .A4(new_n549), .ZN(G188));
  INV_X1    g125(.A(KEYINPUT76), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n509), .A2(new_n551), .A3(G53), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT9), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n524), .A2(G91), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n512), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n555));
  OAI211_X1 g130(.A(new_n553), .B(new_n554), .C1(new_n517), .C2(new_n555), .ZN(G299));
  INV_X1    g131(.A(G171), .ZN(G301));
  NAND2_X1  g132(.A1(new_n509), .A2(G49), .ZN(new_n558));
  OAI21_X1  g133(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n559));
  INV_X1    g134(.A(G87), .ZN(new_n560));
  OAI211_X1 g135(.A(new_n558), .B(new_n559), .C1(new_n560), .C2(new_n513), .ZN(G288));
  NAND2_X1  g136(.A1(new_n509), .A2(G48), .ZN(new_n562));
  INV_X1    g137(.A(G86), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n513), .B2(new_n563), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n512), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n565), .A2(new_n517), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(G305));
  AOI22_X1  g143(.A1(new_n524), .A2(G85), .B1(G47), .B2(new_n509), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n517), .B2(new_n570), .ZN(G290));
  NAND2_X1  g146(.A1(G301), .A2(G868), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n524), .A2(G92), .ZN(new_n573));
  XOR2_X1   g148(.A(new_n573), .B(KEYINPUT10), .Z(new_n574));
  NAND2_X1  g149(.A1(new_n512), .A2(G66), .ZN(new_n575));
  INV_X1    g150(.A(G79), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n576), .B2(new_n506), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n577), .A2(G651), .B1(G54), .B2(new_n509), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n572), .B1(new_n580), .B2(G868), .ZN(G284));
  XNOR2_X1  g156(.A(G284), .B(KEYINPUT77), .ZN(G321));
  INV_X1    g157(.A(G868), .ZN(new_n583));
  NOR2_X1   g158(.A1(G286), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g159(.A(G299), .B(KEYINPUT78), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n584), .B1(new_n583), .B2(new_n585), .ZN(G297));
  AOI21_X1  g161(.A(new_n584), .B1(new_n583), .B2(new_n585), .ZN(G280));
  INV_X1    g162(.A(G559), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n580), .B1(new_n588), .B2(G860), .ZN(G148));
  NAND2_X1  g164(.A1(new_n580), .A2(new_n588), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT79), .ZN(new_n591));
  MUX2_X1   g166(.A(new_n544), .B(new_n591), .S(G868), .Z(G323));
  XNOR2_X1  g167(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g168(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n594));
  INV_X1    g169(.A(G111), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n594), .B1(new_n595), .B2(G2105), .ZN(new_n596));
  INV_X1    g171(.A(new_n469), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n596), .B1(new_n597), .B2(G135), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n599), .B1(new_n487), .B2(G123), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  OR2_X1    g176(.A1(new_n601), .A2(G2096), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(G2096), .ZN(new_n603));
  XNOR2_X1  g178(.A(KEYINPUT80), .B(G2100), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT13), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n467), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n606));
  XOR2_X1   g181(.A(new_n606), .B(KEYINPUT12), .Z(new_n607));
  XNOR2_X1  g182(.A(new_n605), .B(new_n607), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n602), .A2(new_n603), .A3(new_n608), .ZN(G156));
  XOR2_X1   g184(.A(G2451), .B(G2454), .Z(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT16), .ZN(new_n611));
  XNOR2_X1  g186(.A(G1341), .B(G1348), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT81), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n611), .B(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT14), .ZN(new_n615));
  XNOR2_X1  g190(.A(G2427), .B(G2438), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(G2430), .ZN(new_n617));
  XNOR2_X1  g192(.A(KEYINPUT15), .B(G2435), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n615), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(new_n618), .B2(new_n617), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n614), .B(new_n620), .Z(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(G2443), .B(G2446), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(G14), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n625), .B1(new_n624), .B2(new_n622), .ZN(G401));
  XNOR2_X1  g201(.A(G2072), .B(G2078), .ZN(new_n627));
  INV_X1    g202(.A(KEYINPUT82), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT17), .Z(new_n630));
  XNOR2_X1  g205(.A(G2067), .B(G2678), .ZN(new_n631));
  INV_X1    g206(.A(new_n631), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2084), .B(G2090), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(new_n629), .B2(new_n631), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT83), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n632), .A2(new_n634), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n629), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT18), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n631), .A2(new_n634), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n640), .B1(new_n630), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n637), .A2(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(G2100), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT84), .B(G2096), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n643), .B(G2100), .ZN(new_n648));
  INV_X1    g223(.A(new_n646), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n647), .A2(new_n650), .ZN(G227));
  XOR2_X1   g226(.A(G1971), .B(G1976), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT19), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1956), .B(G2474), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1961), .B(G1966), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AND2_X1   g231(.A1(new_n654), .A2(new_n655), .ZN(new_n657));
  NOR3_X1   g232(.A1(new_n653), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n653), .A2(new_n656), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT20), .Z(new_n660));
  AOI211_X1 g235(.A(new_n658), .B(new_n660), .C1(new_n653), .C2(new_n657), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1991), .B(G1996), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1981), .B(G1986), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(G229));
  INV_X1    g243(.A(G16), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(G22), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n670), .B1(G166), .B2(new_n669), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(G1971), .Z(new_n672));
  NOR2_X1   g247(.A1(G16), .A2(G23), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT86), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n674), .B1(G288), .B2(new_n669), .ZN(new_n675));
  XOR2_X1   g250(.A(KEYINPUT33), .B(G1976), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  NOR2_X1   g252(.A1(G6), .A2(G16), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n678), .B1(new_n567), .B2(G16), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT32), .B(G1981), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n672), .A2(new_n677), .A3(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT34), .Z(new_n683));
  NOR2_X1   g258(.A1(G25), .A2(G29), .ZN(new_n684));
  OAI21_X1  g259(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n685));
  INV_X1    g260(.A(G107), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n685), .B1(new_n686), .B2(G2105), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT85), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n688), .B1(G131), .B2(new_n597), .ZN(new_n689));
  INV_X1    g264(.A(G119), .ZN(new_n690));
  INV_X1    g265(.A(new_n487), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n689), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n684), .B1(new_n693), .B2(G29), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT35), .B(G1991), .Z(new_n696));
  OR2_X1    g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n695), .A2(new_n696), .ZN(new_n698));
  MUX2_X1   g273(.A(G24), .B(G290), .S(G16), .Z(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(G1986), .Z(new_n700));
  NAND4_X1  g275(.A1(new_n683), .A2(new_n697), .A3(new_n698), .A4(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT36), .ZN(new_n702));
  INV_X1    g277(.A(KEYINPUT90), .ZN(new_n703));
  INV_X1    g278(.A(G129), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(new_n483), .B2(new_n486), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n467), .A2(G105), .A3(G2104), .ZN(new_n707));
  OR2_X1    g282(.A1(KEYINPUT89), .A2(KEYINPUT26), .ZN(new_n708));
  NAND3_X1  g283(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n709));
  NAND2_X1  g284(.A1(KEYINPUT89), .A2(KEYINPUT26), .ZN(new_n710));
  AND3_X1   g285(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n709), .B1(new_n708), .B2(new_n710), .ZN(new_n712));
  INV_X1    g287(.A(G141), .ZN(new_n713));
  OAI221_X1 g288(.A(new_n707), .B1(new_n711), .B2(new_n712), .C1(new_n713), .C2(new_n469), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n703), .B1(new_n706), .B2(new_n715), .ZN(new_n716));
  NOR3_X1   g291(.A1(new_n705), .A2(new_n714), .A3(KEYINPUT90), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G29), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G29), .B2(G32), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT27), .B(G1996), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT91), .Z(new_n723));
  INV_X1    g298(.A(G29), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G33), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n597), .A2(G139), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT25), .Z(new_n728));
  AND2_X1   g303(.A1(new_n472), .A2(new_n468), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n729), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n726), .B(new_n728), .C1(new_n467), .C2(new_n730), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT87), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n725), .B1(new_n732), .B2(new_n724), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT88), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(G2072), .ZN(new_n735));
  INV_X1    g310(.A(G2084), .ZN(new_n736));
  INV_X1    g311(.A(G34), .ZN(new_n737));
  AOI21_X1  g312(.A(G29), .B1(new_n737), .B2(KEYINPUT24), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(KEYINPUT24), .B2(new_n737), .ZN(new_n739));
  INV_X1    g314(.A(G160), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n739), .B1(new_n740), .B2(new_n724), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n723), .B(new_n735), .C1(new_n736), .C2(new_n741), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n742), .A2(KEYINPUT92), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(KEYINPUT92), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n669), .A2(G21), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G168), .B2(new_n669), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G1966), .ZN(new_n747));
  AOI21_X1  g322(.A(KEYINPUT23), .B1(new_n669), .B2(G20), .ZN(new_n748));
  AND3_X1   g323(.A1(new_n669), .A2(KEYINPUT23), .A3(G20), .ZN(new_n749));
  AOI211_X1 g324(.A(new_n748), .B(new_n749), .C1(G299), .C2(G16), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT93), .B(G1956), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n751), .A2(new_n752), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n741), .A2(new_n736), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n753), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(G4), .A2(G16), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n580), .B2(G16), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G1348), .ZN(new_n759));
  INV_X1    g334(.A(G28), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n760), .A2(KEYINPUT30), .ZN(new_n761));
  AOI21_X1  g336(.A(G29), .B1(new_n760), .B2(KEYINPUT30), .ZN(new_n762));
  OR2_X1    g337(.A1(KEYINPUT31), .A2(G11), .ZN(new_n763));
  NAND2_X1  g338(.A1(KEYINPUT31), .A2(G11), .ZN(new_n764));
  AOI22_X1  g339(.A1(new_n761), .A2(new_n762), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n545), .A2(G16), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G16), .B2(G19), .ZN(new_n767));
  INV_X1    g342(.A(G1341), .ZN(new_n768));
  OAI221_X1 g343(.A(new_n765), .B1(new_n724), .B2(new_n601), .C1(new_n767), .C2(new_n768), .ZN(new_n769));
  OR4_X1    g344(.A1(new_n747), .A2(new_n756), .A3(new_n759), .A4(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n720), .A2(new_n721), .ZN(new_n771));
  INV_X1    g346(.A(G2090), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n724), .A2(G35), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G162), .B2(new_n724), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT29), .Z(new_n775));
  AOI21_X1  g350(.A(new_n771), .B1(new_n772), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n772), .B2(new_n775), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n724), .A2(G26), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT28), .ZN(new_n779));
  INV_X1    g354(.A(G128), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n483), .B2(new_n486), .ZN(new_n781));
  INV_X1    g356(.A(G140), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n467), .A2(G116), .ZN(new_n783));
  OAI21_X1  g358(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n784));
  OAI22_X1  g359(.A1(new_n469), .A2(new_n782), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n779), .B1(new_n786), .B2(new_n724), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G2067), .ZN(new_n788));
  NOR2_X1   g363(.A1(G164), .A2(new_n724), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G27), .B2(new_n724), .ZN(new_n790));
  INV_X1    g365(.A(G2078), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n767), .A2(new_n768), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n790), .A2(new_n791), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n669), .A2(G5), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G171), .B2(new_n669), .ZN(new_n796));
  INV_X1    g371(.A(G1961), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n792), .A2(new_n793), .A3(new_n794), .A4(new_n798), .ZN(new_n799));
  NOR4_X1   g374(.A1(new_n770), .A2(new_n777), .A3(new_n788), .A4(new_n799), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n702), .A2(new_n743), .A3(new_n744), .A4(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(G311));
  XOR2_X1   g377(.A(new_n801), .B(KEYINPUT94), .Z(G150));
  NAND2_X1  g378(.A1(new_n580), .A2(G559), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT38), .ZN(new_n805));
  AOI22_X1  g380(.A1(new_n524), .A2(G93), .B1(G55), .B2(new_n509), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n806), .B1(new_n517), .B2(new_n807), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n544), .B(new_n808), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n805), .B(new_n809), .Z(new_n810));
  AND2_X1   g385(.A1(new_n810), .A2(KEYINPUT39), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n810), .A2(KEYINPUT39), .ZN(new_n812));
  NOR3_X1   g387(.A1(new_n811), .A2(new_n812), .A3(G860), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n808), .A2(G860), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT95), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT37), .Z(new_n816));
  NOR2_X1   g391(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT96), .Z(G145));
  XNOR2_X1  g393(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT99), .B(G37), .Z(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT97), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n487), .A2(G128), .ZN(new_n824));
  INV_X1    g399(.A(new_n785), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n823), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NOR3_X1   g401(.A1(new_n781), .A2(KEYINPUT97), .A3(new_n785), .ZN(new_n827));
  NOR3_X1   g402(.A1(new_n826), .A2(new_n827), .A3(new_n504), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n824), .A2(new_n823), .A3(new_n825), .ZN(new_n829));
  OAI21_X1  g404(.A(KEYINPUT97), .B1(new_n781), .B2(new_n785), .ZN(new_n830));
  AOI21_X1  g405(.A(G164), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OAI22_X1  g406(.A1(new_n828), .A2(new_n831), .B1(new_n716), .B2(new_n717), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n504), .B1(new_n826), .B2(new_n827), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n829), .A2(new_n830), .A3(G164), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n718), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n832), .A2(new_n732), .A3(new_n835), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n705), .A2(new_n714), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(new_n828), .B2(new_n831), .ZN(new_n838));
  INV_X1    g413(.A(new_n837), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n833), .A2(new_n839), .A3(new_n834), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n838), .A2(new_n840), .A3(new_n731), .ZN(new_n841));
  AND3_X1   g416(.A1(new_n836), .A2(new_n841), .A3(new_n692), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n692), .B1(new_n836), .B2(new_n841), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n607), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n836), .A2(new_n841), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(new_n693), .ZN(new_n846));
  INV_X1    g421(.A(new_n607), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n836), .A2(new_n841), .A3(new_n692), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  OR2_X1    g424(.A1(G106), .A2(G2105), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n850), .B(G2104), .C1(G118), .C2(new_n467), .ZN(new_n851));
  INV_X1    g426(.A(G142), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n851), .B1(new_n469), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n853), .B1(new_n487), .B2(G130), .ZN(new_n854));
  AND3_X1   g429(.A1(new_n844), .A2(new_n849), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n854), .B1(new_n844), .B2(new_n849), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n600), .B(G160), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(G162), .Z(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n822), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT100), .ZN(new_n862));
  INV_X1    g437(.A(new_n854), .ZN(new_n863));
  NOR3_X1   g438(.A1(new_n842), .A2(new_n843), .A3(new_n607), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n847), .B1(new_n846), .B2(new_n848), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n844), .A2(new_n849), .A3(new_n854), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(KEYINPUT98), .B1(new_n868), .B2(new_n859), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT98), .ZN(new_n870));
  AOI211_X1 g445(.A(new_n870), .B(new_n860), .C1(new_n866), .C2(new_n867), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n861), .B(new_n862), .C1(new_n869), .C2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n859), .B1(new_n855), .B2(new_n856), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(new_n870), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n868), .A2(KEYINPUT98), .A3(new_n859), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n862), .B1(new_n877), .B2(new_n861), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n820), .B1(new_n873), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n861), .B1(new_n869), .B2(new_n871), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(KEYINPUT100), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n881), .A2(new_n872), .A3(new_n819), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n879), .A2(new_n882), .ZN(G395));
  NAND2_X1  g458(.A1(new_n808), .A2(new_n583), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n591), .B(new_n809), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n579), .B(G299), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n886), .B(KEYINPUT41), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n887), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  XOR2_X1   g464(.A(G303), .B(KEYINPUT102), .Z(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(G290), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n567), .B(G288), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n891), .B(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(KEYINPUT42), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n889), .B(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n884), .B1(new_n895), .B2(new_n583), .ZN(G295));
  OAI21_X1  g471(.A(new_n884), .B1(new_n895), .B2(new_n583), .ZN(G331));
  INV_X1    g472(.A(KEYINPUT44), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n809), .B(G301), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(G286), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(new_n888), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n901), .B1(new_n886), .B2(new_n900), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n893), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n903), .B1(KEYINPUT103), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(G37), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT103), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n902), .A2(new_n907), .A3(new_n893), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n905), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n909), .A2(KEYINPUT43), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n822), .B1(new_n902), .B2(new_n893), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n911), .B1(new_n893), .B2(new_n902), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n912), .A2(KEYINPUT43), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n898), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n898), .B1(new_n912), .B2(KEYINPUT43), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT104), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT43), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n905), .A2(new_n917), .A3(new_n906), .A4(new_n908), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n915), .A2(new_n916), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n916), .B1(new_n915), .B2(new_n918), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n914), .B1(new_n919), .B2(new_n920), .ZN(G397));
  INV_X1    g496(.A(KEYINPUT126), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n786), .B(G2067), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n924), .B1(G1996), .B2(new_n839), .ZN(new_n925));
  INV_X1    g500(.A(G1996), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n718), .A2(new_n926), .ZN(new_n927));
  OR2_X1    g502(.A1(new_n693), .A2(new_n696), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n693), .A2(new_n696), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n925), .A2(new_n927), .A3(new_n928), .A4(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(G290), .A2(G1986), .ZN(new_n931));
  AND2_X1   g506(.A1(G290), .A2(G1986), .ZN(new_n932));
  OR3_X1    g507(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n491), .A2(new_n492), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n495), .A2(new_n497), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n469), .A2(new_n489), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n500), .B(new_n501), .ZN(new_n939));
  AOI21_X1  g514(.A(G1384), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(G160), .A2(G40), .ZN(new_n941));
  NOR3_X1   g516(.A1(new_n940), .A2(new_n941), .A3(KEYINPUT45), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n933), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(G8), .ZN(new_n945));
  INV_X1    g520(.A(G1966), .ZN(new_n946));
  INV_X1    g521(.A(G40), .ZN(new_n947));
  NOR4_X1   g522(.A1(new_n471), .A2(new_n475), .A3(new_n947), .A4(new_n476), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n948), .B1(new_n940), .B2(KEYINPUT45), .ZN(new_n949));
  INV_X1    g524(.A(G1384), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n504), .A2(KEYINPUT45), .A3(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  OAI211_X1 g527(.A(KEYINPUT110), .B(new_n946), .C1(new_n949), .C2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT50), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n940), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n502), .A2(new_n503), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n934), .B(new_n935), .C1(new_n469), .C2(new_n489), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n950), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT50), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n955), .A2(new_n959), .A3(new_n736), .A4(new_n948), .ZN(new_n960));
  AND2_X1   g535(.A1(new_n953), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT45), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n941), .B1(new_n958), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n951), .ZN(new_n964));
  AOI21_X1  g539(.A(KEYINPUT110), .B1(new_n964), .B2(new_n946), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n945), .B1(new_n961), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(G168), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(G303), .A2(G8), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n970), .B(KEYINPUT55), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(KEYINPUT105), .B(G1971), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n973), .B1(new_n963), .B2(new_n951), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n955), .A2(new_n959), .A3(new_n948), .ZN(new_n975));
  OAI22_X1  g550(.A1(new_n974), .A2(KEYINPUT106), .B1(G2090), .B2(new_n975), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n974), .A2(KEYINPUT106), .ZN(new_n977));
  OAI211_X1 g552(.A(G8), .B(new_n972), .C1(new_n976), .C2(new_n977), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n958), .A2(new_n941), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n979), .A2(new_n945), .ZN(new_n980));
  INV_X1    g555(.A(G1976), .ZN(new_n981));
  OR2_X1    g556(.A1(G288), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(KEYINPUT52), .B1(G288), .B2(new_n981), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n980), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT49), .ZN(new_n985));
  XOR2_X1   g560(.A(KEYINPUT107), .B(G1981), .Z(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n567), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(G1981), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n567), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n985), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n988), .B(KEYINPUT49), .C1(new_n990), .C2(new_n567), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n980), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n940), .A2(new_n948), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n995), .A2(G8), .A3(new_n982), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT52), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n984), .A2(new_n994), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT63), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(G8), .B1(new_n976), .B2(new_n977), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n971), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n969), .A2(new_n978), .A3(new_n1000), .A4(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT109), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n998), .A2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n984), .A2(new_n994), .A3(KEYINPUT109), .A4(new_n997), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n975), .A2(G2090), .ZN(new_n1007));
  OAI21_X1  g582(.A(G8), .B1(new_n1007), .B2(new_n974), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(new_n971), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n978), .A2(new_n1005), .A3(new_n1006), .A4(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n999), .B1(new_n1010), .B2(new_n968), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1003), .A2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g587(.A1(G288), .A2(G1976), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n989), .B1(new_n994), .B2(new_n1013), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n1014), .A2(KEYINPUT108), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n980), .B1(new_n1014), .B2(KEYINPUT108), .ZN(new_n1016));
  OR2_X1    g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n1012), .B(new_n1017), .C1(new_n978), .C2(new_n998), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT122), .ZN(new_n1019));
  NOR2_X1   g594(.A1(G168), .A2(new_n945), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1021), .B1(new_n961), .B2(new_n966), .ZN(new_n1022));
  XOR2_X1   g597(.A(KEYINPUT118), .B(KEYINPUT51), .Z(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n953), .A2(new_n960), .ZN(new_n1025));
  OAI21_X1  g600(.A(G8), .B1(new_n1025), .B2(new_n965), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1024), .B1(new_n1026), .B2(new_n1021), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT119), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1020), .A2(KEYINPUT51), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1028), .B1(new_n1026), .B2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1026), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1022), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT62), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1019), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1027), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(KEYINPUT119), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1036), .A2(new_n1038), .A3(new_n1032), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1022), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1041), .A2(KEYINPUT122), .A3(KEYINPUT62), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1035), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1010), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n963), .A2(KEYINPUT53), .A3(new_n791), .A4(new_n951), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT120), .ZN(new_n1046));
  OR2_X1    g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n963), .A2(new_n791), .A3(new_n951), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n1049));
  AOI22_X1  g624(.A1(new_n1048), .A2(new_n1049), .B1(new_n975), .B2(new_n797), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1048), .A2(new_n1046), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1047), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  AND2_X1   g627(.A1(new_n1052), .A2(G171), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1044), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1054), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1018), .B1(new_n1043), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(G1348), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n975), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(G2067), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n948), .A2(new_n504), .A3(new_n950), .A4(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g635(.A(new_n1060), .B(KEYINPUT112), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1062), .A2(new_n579), .ZN(new_n1063));
  XOR2_X1   g638(.A(G299), .B(KEYINPUT57), .Z(new_n1064));
  XNOR2_X1  g639(.A(KEYINPUT56), .B(G2072), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n963), .A2(new_n951), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT111), .ZN(new_n1067));
  INV_X1    g642(.A(G1956), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n975), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT111), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n963), .A2(new_n1070), .A3(new_n951), .A4(new_n1065), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1064), .A2(new_n1067), .A3(new_n1069), .A4(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1063), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1067), .A2(new_n1069), .A3(new_n1071), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1064), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  AND2_X1   g651(.A1(new_n1073), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT60), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT115), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1078), .B1(new_n580), .B2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1080), .A2(new_n1061), .A3(new_n1058), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT60), .B1(new_n1058), .B2(new_n1061), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n580), .A2(new_n1079), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1081), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1083), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1062), .A2(new_n1080), .A3(new_n1085), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1084), .A2(new_n1086), .A3(KEYINPUT116), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT116), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT61), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1090), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1091));
  XNOR2_X1  g666(.A(KEYINPUT58), .B(G1341), .ZN(new_n1092));
  OAI22_X1  g667(.A1(new_n964), .A2(G1996), .B1(new_n979), .B2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n544), .A2(KEYINPUT113), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(KEYINPUT59), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1093), .A2(new_n1097), .A3(new_n1094), .ZN(new_n1098));
  AOI22_X1  g673(.A1(new_n1091), .A2(new_n1072), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT114), .ZN(new_n1100));
  AND3_X1   g675(.A1(new_n1076), .A2(new_n1100), .A3(new_n1072), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1090), .B1(new_n1076), .B2(new_n1100), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1099), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1077), .B1(new_n1089), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT117), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1077), .B(KEYINPUT117), .C1(new_n1089), .C2(new_n1103), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT54), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1050), .A2(new_n1045), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1109), .A2(G171), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1108), .B1(new_n1053), .B2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1108), .B1(new_n1109), .B2(G171), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1047), .A2(new_n1050), .A3(G301), .A4(new_n1051), .ZN(new_n1113));
  AND3_X1   g688(.A1(new_n1112), .A2(KEYINPUT121), .A3(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(KEYINPUT121), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1111), .B(new_n1044), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1116), .A2(new_n1033), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1106), .A2(new_n1107), .A3(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n944), .B1(new_n1056), .B2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n942), .B1(new_n924), .B2(new_n839), .ZN(new_n1120));
  XNOR2_X1  g695(.A(new_n1120), .B(KEYINPUT125), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n942), .A2(new_n926), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT46), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  XOR2_X1   g699(.A(new_n1124), .B(KEYINPUT124), .Z(new_n1125));
  NAND2_X1  g700(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1126));
  XOR2_X1   g701(.A(new_n1126), .B(KEYINPUT123), .Z(new_n1127));
  NAND3_X1  g702(.A1(new_n1121), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT47), .ZN(new_n1129));
  OR2_X1    g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n786), .A2(new_n1059), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n925), .A2(new_n927), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1131), .B1(new_n1132), .B2(new_n929), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n930), .A2(new_n942), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n942), .A2(new_n931), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n1135), .B(KEYINPUT48), .ZN(new_n1136));
  AOI22_X1  g711(.A1(new_n942), .A2(new_n1133), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1138));
  AND3_X1   g713(.A1(new_n1130), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n922), .B1(new_n1119), .B2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(KEYINPUT122), .B1(new_n1041), .B2(KEYINPUT62), .ZN(new_n1142));
  AOI211_X1 g717(.A(new_n1019), .B(new_n1034), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1055), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1018), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1118), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(new_n943), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1147), .A2(KEYINPUT126), .A3(new_n1139), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1141), .A2(new_n1148), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g724(.A1(G401), .A2(new_n460), .ZN(new_n1151));
  NAND3_X1  g725(.A1(new_n647), .A2(new_n650), .A3(new_n1151), .ZN(new_n1152));
  AND2_X1   g726(.A1(new_n1152), .A2(KEYINPUT127), .ZN(new_n1153));
  NOR2_X1   g727(.A1(new_n1152), .A2(KEYINPUT127), .ZN(new_n1154));
  NOR3_X1   g728(.A1(G229), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  OAI21_X1  g729(.A(new_n1155), .B1(new_n910), .B2(new_n913), .ZN(new_n1156));
  AOI21_X1  g730(.A(new_n1156), .B1(new_n881), .B2(new_n872), .ZN(G308));
  OAI221_X1 g731(.A(new_n1155), .B1(new_n910), .B2(new_n913), .C1(new_n873), .C2(new_n878), .ZN(G225));
endmodule


