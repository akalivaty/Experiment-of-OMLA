//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 1 0 1 0 1 0 1 0 1 1 1 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 0 0 0 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:54 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  NOR2_X1   g001(.A1(G237), .A2(G953), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G210), .ZN(new_n189));
  INV_X1    g003(.A(G101), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n192));
  XOR2_X1   g006(.A(new_n191), .B(new_n192), .Z(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT1), .B1(new_n194), .B2(G146), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n194), .A2(G146), .ZN(new_n196));
  INV_X1    g010(.A(G146), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(G143), .ZN(new_n198));
  OAI211_X1 g012(.A(G128), .B(new_n195), .C1(new_n196), .C2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(G143), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n194), .A2(G146), .ZN(new_n201));
  INV_X1    g015(.A(G128), .ZN(new_n202));
  OAI211_X1 g016(.A(new_n200), .B(new_n201), .C1(KEYINPUT1), .C2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G134), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(G137), .ZN(new_n205));
  INV_X1    g019(.A(G137), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n206), .A2(G134), .ZN(new_n207));
  OAI21_X1  g021(.A(G131), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n199), .A2(new_n203), .A3(new_n208), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n206), .B(G134), .C1(KEYINPUT64), .C2(KEYINPUT11), .ZN(new_n210));
  AOI22_X1  g024(.A1(new_n204), .A2(G137), .B1(KEYINPUT64), .B2(KEYINPUT11), .ZN(new_n211));
  AND2_X1   g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G131), .ZN(new_n213));
  NOR2_X1   g027(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n214), .B1(new_n204), .B2(G137), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n212), .A2(KEYINPUT65), .A3(new_n213), .A4(new_n215), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n215), .A2(new_n210), .A3(new_n211), .A4(new_n213), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT65), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n209), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n215), .A2(new_n210), .A3(new_n211), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G131), .ZN(new_n222));
  AND2_X1   g036(.A1(new_n217), .A2(new_n218), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n217), .A2(new_n218), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n200), .A2(new_n201), .A3(KEYINPUT0), .A4(G128), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n196), .A2(new_n198), .ZN(new_n227));
  XNOR2_X1  g041(.A(KEYINPUT0), .B(G128), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n226), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n220), .B1(new_n225), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g045(.A(G116), .B(G119), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT67), .B1(new_n232), .B2(KEYINPUT66), .ZN(new_n233));
  INV_X1    g047(.A(G119), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G116), .ZN(new_n235));
  INV_X1    g049(.A(G116), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G119), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT66), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT67), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  XOR2_X1   g055(.A(KEYINPUT2), .B(G113), .Z(new_n242));
  AND3_X1   g056(.A1(new_n233), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n242), .B1(new_n233), .B2(new_n241), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n231), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  AND2_X1   g062(.A1(new_n199), .A2(new_n203), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n249), .B(new_n208), .C1(new_n223), .C2(new_n224), .ZN(new_n250));
  AOI22_X1  g064(.A1(new_n216), .A2(new_n219), .B1(G131), .B2(new_n221), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n250), .B1(new_n251), .B2(new_n229), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n253), .B1(new_n243), .B2(new_n244), .ZN(new_n254));
  INV_X1    g068(.A(new_n242), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n240), .B1(new_n238), .B2(new_n239), .ZN(new_n256));
  AOI211_X1 g070(.A(KEYINPUT66), .B(KEYINPUT67), .C1(new_n235), .C2(new_n237), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n233), .A2(new_n241), .A3(new_n242), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n258), .A2(KEYINPUT68), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n254), .A2(new_n260), .ZN(new_n261));
  NOR3_X1   g075(.A1(new_n252), .A2(new_n261), .A3(KEYINPUT69), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n263));
  NOR3_X1   g077(.A1(new_n243), .A2(new_n244), .A3(new_n253), .ZN(new_n264));
  AOI21_X1  g078(.A(KEYINPUT68), .B1(new_n258), .B2(new_n259), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n263), .B1(new_n266), .B2(new_n231), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n248), .B1(new_n262), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT28), .ZN(new_n269));
  AOI21_X1  g083(.A(KEYINPUT28), .B1(new_n266), .B2(new_n231), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n193), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT30), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n216), .A2(new_n219), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n229), .B1(new_n274), .B2(new_n222), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n273), .B1(new_n275), .B2(new_n220), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n250), .B(KEYINPUT30), .C1(new_n251), .C2(new_n229), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n276), .A2(new_n245), .A3(new_n277), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n193), .B(new_n278), .C1(new_n262), .C2(new_n267), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT31), .ZN(new_n280));
  OAI21_X1  g094(.A(KEYINPUT69), .B1(new_n252), .B2(new_n261), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n266), .A2(new_n263), .A3(new_n231), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT31), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n283), .A2(new_n284), .A3(new_n193), .A4(new_n278), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n280), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n187), .B1(new_n272), .B2(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT32), .B1(new_n287), .B2(KEYINPUT70), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT70), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT32), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n270), .B1(new_n268), .B2(KEYINPUT28), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n280), .B(new_n285), .C1(new_n291), .C2(new_n193), .ZN(new_n292));
  AOI211_X1 g106(.A(new_n289), .B(new_n290), .C1(new_n292), .C2(new_n187), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT71), .ZN(new_n294));
  INV_X1    g108(.A(G472), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n193), .A2(KEYINPUT29), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  AOI22_X1  g111(.A1(new_n281), .A2(new_n282), .B1(new_n261), .B2(new_n252), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT28), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n271), .B(new_n297), .C1(new_n298), .C2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G902), .ZN(new_n301));
  AND2_X1   g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n278), .B1(new_n262), .B2(new_n267), .ZN(new_n303));
  INV_X1    g117(.A(new_n193), .ZN(new_n304));
  AOI21_X1  g118(.A(KEYINPUT29), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n247), .B1(new_n281), .B2(new_n282), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n271), .B(new_n193), .C1(new_n306), .C2(new_n299), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  AOI211_X1 g122(.A(new_n294), .B(new_n295), .C1(new_n302), .C2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(new_n301), .A3(new_n300), .ZN(new_n310));
  AOI21_X1  g124(.A(KEYINPUT71), .B1(new_n310), .B2(G472), .ZN(new_n311));
  OAI22_X1  g125(.A1(new_n288), .A2(new_n293), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G953), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n313), .A2(G221), .A3(G234), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n314), .B(KEYINPUT76), .ZN(new_n315));
  XNOR2_X1  g129(.A(KEYINPUT22), .B(G137), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n315), .B(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  XOR2_X1   g132(.A(KEYINPUT24), .B(G110), .Z(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n234), .A2(G128), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n202), .A2(G119), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT72), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NOR3_X1   g139(.A1(new_n321), .A2(new_n322), .A3(KEYINPUT72), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n320), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G110), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n321), .B1(KEYINPUT73), .B2(KEYINPUT23), .ZN(new_n329));
  OR2_X1    g143(.A1(new_n321), .A2(KEYINPUT73), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT23), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n322), .A2(new_n331), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n328), .B(new_n329), .C1(new_n330), .C2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n327), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(G140), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G125), .ZN(new_n336));
  INV_X1    g150(.A(G125), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G140), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n336), .A2(new_n338), .A3(new_n197), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n334), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT16), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n336), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n338), .A2(KEYINPUT74), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT74), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n344), .A2(new_n337), .A3(G140), .ZN(new_n345));
  AOI22_X1  g159(.A1(new_n343), .A2(new_n345), .B1(G125), .B2(new_n335), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n342), .B1(new_n346), .B2(new_n341), .ZN(new_n347));
  AOI21_X1  g161(.A(KEYINPUT75), .B1(new_n347), .B2(G146), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n347), .A2(KEYINPUT75), .A3(G146), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n340), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n347), .A2(G146), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n197), .B(new_n342), .C1(new_n346), .C2(new_n341), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n325), .A2(new_n326), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n319), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n329), .B1(new_n330), .B2(new_n332), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G110), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n354), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n318), .B1(new_n351), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n350), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n334), .B(new_n339), .C1(new_n361), .C2(new_n348), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n354), .A2(new_n356), .A3(new_n358), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n362), .A2(new_n363), .A3(new_n317), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n360), .A2(new_n364), .A3(new_n301), .ZN(new_n365));
  NOR2_X1   g179(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n366), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n360), .A2(new_n364), .A3(new_n301), .A4(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n367), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G217), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n372), .B1(G234), .B2(new_n301), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  AND2_X1   g188(.A1(new_n360), .A2(new_n364), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n373), .A2(G902), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT13), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n380), .B1(new_n202), .B2(G143), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT90), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n194), .A2(G128), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT90), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n384), .A3(new_n380), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT91), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n202), .A2(G143), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n382), .A2(new_n385), .A3(new_n386), .A4(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n194), .A2(KEYINPUT13), .A3(G128), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  AOI22_X1  g204(.A1(new_n381), .A2(KEYINPUT90), .B1(new_n202), .B2(G143), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n386), .B1(new_n391), .B2(new_n385), .ZN(new_n392));
  OAI21_X1  g206(.A(G134), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT92), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  OAI211_X1 g209(.A(KEYINPUT92), .B(G134), .C1(new_n390), .C2(new_n392), .ZN(new_n396));
  OR2_X1    g210(.A1(new_n236), .A2(G122), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n236), .A2(G122), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  XNOR2_X1  g213(.A(KEYINPUT89), .B(G107), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n399), .B(new_n400), .ZN(new_n401));
  AND3_X1   g215(.A1(new_n383), .A2(new_n387), .A3(new_n204), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n395), .A2(new_n396), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n397), .A2(KEYINPUT14), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n399), .A2(new_n405), .A3(G107), .ZN(new_n406));
  INV_X1    g220(.A(G107), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n397), .B(new_n398), .C1(KEYINPUT14), .C2(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n204), .B1(new_n383), .B2(new_n387), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n406), .B(new_n408), .C1(new_n402), .C2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n404), .A2(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(KEYINPUT9), .B(G234), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n412), .B(KEYINPUT78), .ZN(new_n413));
  NOR3_X1   g227(.A1(new_n413), .A2(new_n372), .A3(G953), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n411), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT93), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n404), .A2(new_n410), .A3(new_n414), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n404), .A2(KEYINPUT93), .A3(new_n410), .A4(new_n414), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n419), .A2(new_n301), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(G478), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n422), .A2(KEYINPUT15), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n423), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n419), .A2(new_n301), .A3(new_n420), .A4(new_n425), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n424), .A2(KEYINPUT94), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(KEYINPUT94), .B1(new_n424), .B2(new_n426), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G475), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n188), .A2(G143), .A3(G214), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(G143), .B1(new_n188), .B2(G214), .ZN(new_n433));
  OAI21_X1  g247(.A(G131), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT17), .ZN(new_n435));
  OR2_X1    g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n433), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n437), .A2(new_n213), .A3(new_n431), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n434), .A2(new_n438), .A3(new_n435), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n352), .A2(new_n436), .A3(new_n353), .A4(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(KEYINPUT18), .A2(G131), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n437), .A2(new_n431), .A3(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n339), .B1(new_n346), .B2(new_n197), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT18), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n442), .B(new_n443), .C1(new_n444), .C2(new_n434), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n440), .A2(new_n445), .ZN(new_n446));
  XNOR2_X1  g260(.A(G113), .B(G122), .ZN(new_n447));
  INV_X1    g261(.A(G104), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n447), .B(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n446), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n440), .A2(new_n449), .A3(new_n445), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n430), .B1(new_n453), .B2(new_n301), .ZN(new_n454));
  NOR2_X1   g268(.A1(G475), .A2(G902), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT19), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n336), .A2(new_n338), .A3(new_n456), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n197), .B(new_n457), .C1(new_n346), .C2(new_n456), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n434), .A2(new_n438), .ZN(new_n459));
  AND2_X1   g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n460), .B1(new_n361), .B2(new_n348), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n449), .B1(new_n461), .B2(new_n445), .ZN(new_n462));
  INV_X1    g276(.A(new_n452), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n455), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT20), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT20), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n466), .B(new_n455), .C1(new_n462), .C2(new_n463), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n454), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(G234), .A2(G237), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n469), .A2(G952), .A3(new_n313), .ZN(new_n470));
  XOR2_X1   g284(.A(KEYINPUT21), .B(G898), .Z(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n469), .A2(G902), .A3(G953), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n470), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n468), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n429), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT3), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n478), .A2(new_n407), .A3(G104), .ZN(new_n479));
  AOI21_X1  g293(.A(KEYINPUT3), .B1(new_n448), .B2(G107), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n448), .A2(G107), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(G101), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n190), .B(new_n479), .C1(new_n480), .C2(new_n481), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n483), .A2(KEYINPUT4), .A3(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT4), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n482), .A2(new_n486), .A3(G101), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n485), .A2(new_n230), .A3(new_n487), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n407), .A2(G104), .ZN(new_n489));
  OAI21_X1  g303(.A(G101), .B1(new_n481), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n484), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(new_n249), .A3(KEYINPUT10), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n488), .A2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  XOR2_X1   g309(.A(KEYINPUT80), .B(KEYINPUT10), .Z(new_n496));
  INV_X1    g310(.A(KEYINPUT79), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n497), .B1(new_n492), .B2(new_n249), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n199), .A2(new_n203), .ZN(new_n499));
  NOR3_X1   g313(.A1(new_n491), .A2(new_n499), .A3(KEYINPUT79), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n496), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n251), .B1(new_n495), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n496), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n492), .A2(new_n249), .A3(new_n497), .ZN(new_n504));
  OAI21_X1  g318(.A(KEYINPUT79), .B1(new_n491), .B2(new_n499), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NOR3_X1   g320(.A1(new_n506), .A2(new_n494), .A3(new_n225), .ZN(new_n507));
  XNOR2_X1  g321(.A(G110), .B(G140), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n313), .A2(G227), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n508), .B(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NOR3_X1   g325(.A1(new_n502), .A2(new_n507), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n491), .A2(new_n499), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n514), .B1(new_n498), .B2(new_n500), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT12), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n516), .B1(new_n251), .B2(KEYINPUT81), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n515), .A2(new_n517), .A3(new_n225), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT81), .ZN(new_n519));
  AOI21_X1  g333(.A(KEYINPUT12), .B1(new_n225), .B2(new_n519), .ZN(new_n520));
  AOI22_X1  g334(.A1(new_n504), .A2(new_n505), .B1(new_n499), .B2(new_n491), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n520), .B1(new_n521), .B2(new_n251), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n507), .B1(new_n518), .B2(new_n522), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n513), .B(KEYINPUT82), .C1(new_n523), .C2(new_n510), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT82), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n522), .A2(new_n518), .ZN(new_n526));
  INV_X1    g340(.A(new_n507), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n510), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n525), .B1(new_n528), .B2(new_n512), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n524), .A2(new_n529), .A3(new_n301), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n506), .A2(new_n494), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n511), .B1(new_n531), .B2(new_n251), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(new_n526), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n511), .B1(new_n502), .B2(new_n507), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(G469), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n535), .A2(new_n536), .A3(new_n301), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(KEYINPUT83), .ZN(new_n538));
  AOI21_X1  g352(.A(G902), .B1(new_n533), .B2(new_n534), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT83), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n539), .A2(new_n540), .A3(new_n536), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n530), .A2(G469), .B1(new_n538), .B2(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(G214), .B1(G237), .B2(G902), .ZN(new_n543));
  XOR2_X1   g357(.A(new_n543), .B(KEYINPUT84), .Z(new_n544));
  XOR2_X1   g358(.A(new_n544), .B(KEYINPUT85), .Z(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  XOR2_X1   g360(.A(G110), .B(G122), .Z(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n258), .A2(new_n485), .A3(new_n259), .A4(new_n487), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT86), .ZN(new_n550));
  OR3_X1    g364(.A1(new_n235), .A2(new_n550), .A3(KEYINPUT5), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n232), .A2(KEYINPUT5), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n550), .B1(new_n235), .B2(KEYINPUT5), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n551), .A2(new_n552), .A3(G113), .A4(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n242), .A2(new_n232), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n492), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n548), .B1(new_n549), .B2(new_n556), .ZN(new_n557));
  OR2_X1    g371(.A1(new_n557), .A2(KEYINPUT6), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n549), .A2(new_n556), .A3(new_n548), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT87), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n549), .A2(KEYINPUT87), .A3(new_n556), .A4(new_n548), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n557), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT6), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n558), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n229), .A2(G125), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n566), .B1(new_n249), .B2(G125), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT88), .B(G224), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n568), .A2(G953), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n567), .B(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n565), .A2(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(G210), .B1(G237), .B2(G902), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT7), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n567), .B1(new_n573), .B2(new_n569), .ZN(new_n574));
  OR2_X1    g388(.A1(new_n567), .A2(new_n569), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n574), .B1(new_n575), .B2(new_n573), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n547), .B(KEYINPUT8), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n554), .A2(new_n555), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n491), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n577), .B1(new_n579), .B2(new_n556), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n561), .A2(new_n562), .ZN(new_n582));
  AOI21_X1  g396(.A(G902), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  AND3_X1   g397(.A1(new_n571), .A2(new_n572), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n572), .B1(new_n571), .B2(new_n583), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n546), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(G221), .B1(new_n413), .B2(G902), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NOR3_X1   g402(.A1(new_n542), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n312), .A2(new_n379), .A3(new_n477), .A4(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(KEYINPUT95), .B(G101), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n590), .B(new_n591), .ZN(G3));
  AOI21_X1  g406(.A(new_n295), .B1(new_n292), .B2(new_n301), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT96), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n292), .A2(new_n301), .ZN(new_n596));
  AOI22_X1  g410(.A1(G472), .A2(new_n596), .B1(new_n287), .B2(new_n594), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NOR3_X1   g412(.A1(new_n542), .A2(new_n378), .A3(new_n588), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(KEYINPUT97), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT33), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n419), .A2(new_n602), .A3(new_n420), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n416), .A2(KEYINPUT33), .A3(new_n418), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n422), .A2(G902), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n421), .A2(new_n422), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n468), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n544), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n611), .B1(new_n584), .B2(new_n585), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT98), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI211_X1 g428(.A(KEYINPUT98), .B(new_n611), .C1(new_n584), .C2(new_n585), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n614), .A2(new_n475), .A3(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NOR3_X1   g431(.A1(new_n601), .A2(new_n610), .A3(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(KEYINPUT34), .B(G104), .Z(new_n619));
  XOR2_X1   g433(.A(new_n619), .B(KEYINPUT99), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n618), .B(new_n620), .ZN(G6));
  INV_X1    g435(.A(KEYINPUT100), .ZN(new_n622));
  OR2_X1    g436(.A1(new_n454), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n465), .A2(new_n467), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n454), .A2(new_n622), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n616), .A2(new_n429), .A3(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n601), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(G107), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT101), .B(KEYINPUT35), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G9));
  NAND2_X1  g446(.A1(new_n362), .A2(new_n363), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n318), .A2(KEYINPUT36), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(new_n635));
  AOI22_X1  g449(.A1(new_n371), .A2(new_n373), .B1(new_n376), .B2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n598), .A2(new_n477), .A3(new_n589), .A4(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT37), .B(G110), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G12));
  NAND2_X1  g454(.A1(new_n571), .A2(new_n583), .ZN(new_n641));
  INV_X1    g455(.A(new_n572), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n571), .A2(new_n572), .A3(new_n583), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(KEYINPUT98), .B1(new_n645), .B2(new_n611), .ZN(new_n646));
  INV_X1    g460(.A(new_n615), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(G900), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n473), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n470), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NOR4_X1   g467(.A1(new_n427), .A2(new_n428), .A3(new_n626), .A4(new_n653), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n542), .A2(new_n588), .A3(new_n636), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n312), .A2(new_n648), .A3(new_n654), .A4(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G128), .ZN(G30));
  NOR3_X1   g471(.A1(new_n427), .A2(new_n428), .A3(new_n468), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n658), .A2(new_n611), .A3(new_n636), .ZN(new_n659));
  XOR2_X1   g473(.A(new_n659), .B(KEYINPUT105), .Z(new_n660));
  XOR2_X1   g474(.A(new_n652), .B(KEYINPUT39), .Z(new_n661));
  OR3_X1    g475(.A1(new_n542), .A2(new_n588), .A3(new_n661), .ZN(new_n662));
  OR2_X1    g476(.A1(new_n662), .A2(KEYINPUT40), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(KEYINPUT40), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT104), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n279), .B1(new_n193), .B2(new_n298), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT103), .ZN(new_n667));
  AOI21_X1  g481(.A(G902), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  OAI211_X1 g482(.A(new_n279), .B(KEYINPUT103), .C1(new_n193), .C2(new_n298), .ZN(new_n669));
  AOI211_X1 g483(.A(new_n665), .B(new_n295), .C1(new_n668), .C2(new_n669), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n283), .A2(new_n193), .A3(new_n278), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n252), .A2(new_n261), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n193), .B1(new_n283), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n667), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n674), .A2(new_n301), .A3(new_n669), .ZN(new_n675));
  AOI21_X1  g489(.A(KEYINPUT104), .B1(new_n675), .B2(G472), .ZN(new_n676));
  OAI22_X1  g490(.A1(new_n293), .A2(new_n288), .B1(new_n670), .B2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n645), .B(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n660), .A2(new_n663), .A3(new_n664), .A4(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G143), .ZN(G45));
  AOI21_X1  g499(.A(new_n468), .B1(new_n606), .B2(new_n607), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT106), .ZN(new_n687));
  AND3_X1   g501(.A1(new_n686), .A2(new_n687), .A3(new_n652), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n687), .B1(new_n686), .B2(new_n652), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n690), .A2(new_n312), .A3(new_n648), .A4(new_n655), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT107), .B(G146), .Z(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G48));
  INV_X1    g507(.A(new_n187), .ZN(new_n694));
  AND2_X1   g508(.A1(new_n280), .A2(new_n285), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n306), .A2(new_n299), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n304), .B1(new_n696), .B2(new_n270), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n694), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n290), .B1(new_n698), .B2(new_n289), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n287), .A2(KEYINPUT70), .A3(KEYINPUT32), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AND2_X1   g515(.A1(new_n305), .A2(new_n307), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n300), .A2(new_n301), .ZN(new_n703));
  OAI21_X1  g517(.A(G472), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n294), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n310), .A2(KEYINPUT71), .A3(G472), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n378), .B1(new_n701), .B2(new_n707), .ZN(new_n708));
  AND4_X1   g522(.A1(new_n475), .A2(new_n614), .A3(new_n686), .A4(new_n615), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n539), .A2(new_n536), .ZN(new_n710));
  AOI211_X1 g524(.A(new_n588), .B(new_n710), .C1(new_n538), .C2(new_n541), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n708), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(KEYINPUT41), .B(G113), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(G15));
  OR2_X1    g528(.A1(new_n539), .A2(new_n536), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n539), .A2(new_n540), .A3(new_n536), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n540), .B1(new_n539), .B2(new_n536), .ZN(new_n717));
  OAI211_X1 g531(.A(new_n587), .B(new_n715), .C1(new_n716), .C2(new_n717), .ZN(new_n718));
  NOR4_X1   g532(.A1(new_n718), .A2(new_n427), .A3(new_n428), .A4(new_n626), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n616), .A2(new_n312), .A3(new_n379), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G116), .ZN(G18));
  AND3_X1   g535(.A1(new_n614), .A2(new_n615), .A3(new_n711), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n722), .A2(new_n312), .A3(new_n477), .A4(new_n637), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G119), .ZN(G21));
  OAI21_X1  g538(.A(new_n271), .B1(new_n298), .B2(new_n299), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT108), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OAI211_X1 g541(.A(KEYINPUT108), .B(new_n271), .C1(new_n298), .C2(new_n299), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n727), .A2(new_n304), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n694), .B1(new_n729), .B2(new_n695), .ZN(new_n730));
  NOR4_X1   g544(.A1(new_n730), .A2(new_n718), .A3(new_n593), .A4(new_n378), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n731), .A2(new_n616), .A3(new_n658), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G122), .ZN(G24));
  NOR3_X1   g547(.A1(new_n730), .A2(new_n593), .A3(new_n636), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n722), .A2(new_n690), .A3(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G125), .ZN(G27));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n528), .A2(new_n512), .ZN(new_n738));
  OAI21_X1  g552(.A(G469), .B1(new_n738), .B2(G902), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n739), .B1(new_n716), .B2(new_n717), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n587), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n643), .A2(new_n611), .A3(new_n644), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n737), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n538), .A2(new_n541), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n588), .B1(new_n744), .B2(new_n739), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n584), .A2(new_n585), .A3(new_n544), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n745), .A2(KEYINPUT109), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n743), .A2(new_n747), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n688), .A2(new_n689), .A3(KEYINPUT42), .ZN(new_n749));
  AND3_X1   g563(.A1(new_n748), .A2(new_n708), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g564(.A(KEYINPUT106), .B1(new_n610), .B2(new_n653), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n686), .A2(new_n687), .A3(new_n652), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n753), .B1(new_n743), .B2(new_n747), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n287), .A2(new_n290), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n698), .A2(KEYINPUT32), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n755), .B(new_n756), .C1(new_n309), .C2(new_n311), .ZN(new_n757));
  AND3_X1   g571(.A1(new_n757), .A2(KEYINPUT110), .A3(new_n379), .ZN(new_n758));
  AOI21_X1  g572(.A(KEYINPUT110), .B1(new_n757), .B2(new_n379), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n754), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n750), .B1(new_n760), .B2(KEYINPUT42), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G131), .ZN(G33));
  NAND3_X1  g576(.A1(new_n748), .A2(new_n708), .A3(new_n654), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G134), .ZN(G36));
  NAND2_X1  g578(.A1(new_n608), .A2(new_n468), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT43), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n765), .B(new_n766), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n767), .B(new_n637), .C1(new_n597), .C2(new_n595), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT44), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(KEYINPUT111), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n536), .B1(new_n738), .B2(KEYINPUT45), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n524), .A2(new_n529), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n772), .B1(new_n773), .B2(KEYINPUT45), .ZN(new_n774));
  NAND2_X1  g588(.A1(G469), .A2(G902), .ZN(new_n775));
  AOI21_X1  g589(.A(KEYINPUT46), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n774), .A2(KEYINPUT46), .A3(new_n775), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n744), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n587), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n779), .A2(new_n661), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n746), .B(KEYINPUT112), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n782), .B1(new_n769), .B2(new_n768), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n771), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G137), .ZN(G39));
  OR2_X1    g599(.A1(new_n779), .A2(KEYINPUT47), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n779), .A2(KEYINPUT47), .ZN(new_n787));
  NOR4_X1   g601(.A1(new_n753), .A2(new_n312), .A3(new_n379), .A4(new_n742), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(KEYINPUT113), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G140), .ZN(G42));
  NAND2_X1  g605(.A1(new_n767), .A2(new_n470), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(KEYINPUT117), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n682), .A2(new_n544), .A3(new_n731), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT50), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n718), .A2(new_n742), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n678), .A2(new_n379), .A3(new_n470), .A4(new_n798), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n799), .A2(new_n609), .A3(new_n608), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n793), .A2(new_n798), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n800), .B1(new_n802), .B2(new_n734), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n710), .B1(new_n538), .B2(new_n541), .ZN(new_n804));
  AOI22_X1  g618(.A1(new_n786), .A2(new_n787), .B1(new_n588), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n730), .A2(new_n593), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n793), .A2(new_n379), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(new_n781), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n797), .B(new_n803), .C1(new_n805), .C2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(KEYINPUT51), .ZN(new_n810));
  OAI211_X1 g624(.A(G952), .B(new_n313), .C1(new_n799), .C2(new_n610), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n811), .B1(new_n807), .B2(new_n722), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT118), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT48), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n758), .A2(new_n759), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n816), .B1(KEYINPUT118), .B2(KEYINPUT48), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n802), .A2(new_n815), .A3(new_n817), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n813), .B(new_n814), .C1(new_n801), .C2(new_n816), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n812), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  XOR2_X1   g634(.A(new_n820), .B(KEYINPUT119), .Z(new_n821));
  NAND2_X1  g635(.A1(new_n810), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n748), .A2(new_n708), .A3(new_n749), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n741), .A2(new_n737), .A3(new_n742), .ZN(new_n824));
  AOI21_X1  g638(.A(KEYINPUT109), .B1(new_n745), .B2(new_n746), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n690), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n309), .A2(new_n311), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n756), .A2(new_n755), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n379), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT110), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n757), .A2(KEYINPUT110), .A3(new_n379), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n826), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT42), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n823), .B(new_n763), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n712), .A2(new_n720), .A3(new_n723), .A4(new_n732), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n734), .A2(new_n752), .A3(new_n751), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(new_n748), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n424), .A2(new_n426), .ZN(new_n840));
  NOR4_X1   g654(.A1(new_n742), .A2(new_n840), .A3(new_n626), .A4(new_n653), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n312), .A2(new_n655), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n840), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n610), .B1(new_n844), .B2(new_n609), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n645), .A2(new_n475), .A3(new_n546), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n598), .A2(new_n599), .A3(new_n845), .A4(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n638), .A2(new_n848), .A3(new_n590), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n837), .A2(new_n843), .A3(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n836), .A2(KEYINPUT114), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT114), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n712), .A2(new_n720), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n638), .A2(new_n848), .A3(new_n590), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n723), .A2(new_n732), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n312), .A2(new_n841), .ZN(new_n856));
  AOI22_X1  g670(.A1(new_n856), .A2(new_n655), .B1(new_n838), .B2(new_n748), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n853), .A2(new_n854), .A3(new_n855), .A4(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n852), .B1(new_n858), .B2(new_n835), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n656), .A2(new_n735), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT115), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n656), .A2(new_n735), .A3(KEYINPUT115), .ZN(new_n863));
  AND4_X1   g677(.A1(new_n587), .A2(new_n740), .A3(new_n636), .A4(new_n652), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n648), .A2(new_n677), .A3(new_n658), .A4(new_n864), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n865), .A2(KEYINPUT52), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n862), .A2(new_n691), .A3(new_n863), .A4(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n656), .A2(new_n691), .A3(new_n865), .A4(new_n735), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT116), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT52), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n869), .B1(new_n868), .B2(new_n870), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n867), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT53), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n851), .A2(new_n859), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n837), .A2(new_n849), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n876), .A2(new_n761), .A3(new_n763), .A4(new_n857), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n868), .B(KEYINPUT52), .ZN(new_n878));
  OAI21_X1  g692(.A(KEYINPUT53), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n875), .A2(KEYINPUT54), .A3(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n858), .A2(new_n835), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n873), .A2(KEYINPUT53), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n874), .B1(new_n877), .B2(new_n878), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT54), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n880), .A2(new_n885), .ZN(new_n886));
  OAI22_X1  g700(.A1(new_n822), .A2(new_n886), .B1(G952), .B2(G953), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n378), .A2(new_n545), .A3(new_n588), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT49), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n888), .B1(new_n804), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n890), .B1(new_n889), .B2(new_n804), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n681), .A2(new_n765), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n891), .A2(new_n678), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n887), .A2(new_n893), .ZN(G75));
  XOR2_X1   g708(.A(new_n565), .B(new_n570), .Z(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  XNOR2_X1  g710(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n301), .B1(new_n882), .B2(new_n883), .ZN(new_n898));
  AOI211_X1 g712(.A(KEYINPUT56), .B(new_n897), .C1(new_n898), .C2(G210), .ZN(new_n899));
  INV_X1    g713(.A(new_n897), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n882), .A2(new_n883), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n901), .A2(G210), .A3(G902), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT56), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n900), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n896), .B1(new_n899), .B2(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n313), .A2(G952), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n906), .B(KEYINPUT121), .Z(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(G210), .ZN(new_n909));
  AOI211_X1 g723(.A(new_n909), .B(new_n301), .C1(new_n882), .C2(new_n883), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n897), .B1(new_n910), .B2(KEYINPUT56), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n902), .A2(new_n903), .A3(new_n900), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n911), .A2(new_n912), .A3(new_n895), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n905), .A2(new_n908), .A3(new_n913), .ZN(G51));
  AOI211_X1 g728(.A(new_n301), .B(new_n774), .C1(new_n882), .C2(new_n883), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n915), .B(KEYINPUT123), .Z(new_n916));
  NAND2_X1  g730(.A1(new_n901), .A2(KEYINPUT54), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(new_n885), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  XNOR2_X1  g733(.A(KEYINPUT122), .B(KEYINPUT57), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(new_n775), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n535), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n906), .B1(new_n916), .B2(new_n922), .ZN(G54));
  AND3_X1   g737(.A1(new_n898), .A2(KEYINPUT58), .A3(G475), .ZN(new_n924));
  OR2_X1    g738(.A1(new_n462), .A2(new_n463), .ZN(new_n925));
  OAI22_X1  g739(.A1(new_n924), .A2(new_n925), .B1(G952), .B2(new_n313), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n924), .A2(new_n925), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(KEYINPUT124), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT124), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n924), .A2(new_n929), .A3(new_n925), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n926), .B1(new_n928), .B2(new_n930), .ZN(G60));
  NAND2_X1  g745(.A1(new_n603), .A2(new_n604), .ZN(new_n932));
  NAND2_X1  g746(.A1(G478), .A2(G902), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT59), .Z(new_n934));
  NOR2_X1   g748(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n907), .B1(new_n918), .B2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(new_n932), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n934), .B1(new_n880), .B2(new_n885), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n936), .B(KEYINPUT125), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT125), .ZN(new_n940));
  INV_X1    g754(.A(new_n885), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n884), .B1(new_n882), .B2(new_n883), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n935), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n908), .ZN(new_n944));
  INV_X1    g758(.A(new_n934), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n937), .B1(new_n886), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n940), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n939), .A2(new_n947), .ZN(G63));
  NAND2_X1  g762(.A1(G217), .A2(G902), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT60), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n950), .B1(new_n882), .B2(new_n883), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n907), .B1(new_n951), .B2(new_n635), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n952), .B1(new_n375), .B2(new_n951), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT61), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(G66));
  OAI21_X1  g769(.A(G953), .B1(new_n472), .B2(new_n568), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n956), .B1(new_n876), .B2(G953), .ZN(new_n957));
  INV_X1    g771(.A(new_n565), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n958), .B1(G898), .B2(new_n313), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n957), .B(new_n959), .ZN(G69));
  AND3_X1   g774(.A1(new_n862), .A2(new_n691), .A3(new_n863), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n684), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT62), .Z(new_n963));
  XNOR2_X1  g777(.A(new_n845), .B(KEYINPUT127), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n662), .A2(new_n742), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n964), .A2(new_n965), .A3(new_n708), .ZN(new_n966));
  AND2_X1   g780(.A1(new_n784), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n963), .A2(new_n790), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n276), .A2(new_n277), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n457), .B1(new_n346), .B2(new_n456), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT126), .Z(new_n971));
  XNOR2_X1  g785(.A(new_n969), .B(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n968), .A2(new_n313), .A3(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(new_n816), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n974), .A2(new_n648), .A3(new_n658), .ZN(new_n975));
  AOI22_X1  g789(.A1(new_n771), .A2(new_n783), .B1(new_n975), .B2(new_n780), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n976), .A2(new_n790), .A3(new_n836), .A4(new_n961), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n313), .ZN(new_n978));
  INV_X1    g792(.A(new_n972), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n978), .B(new_n979), .C1(G227), .C2(new_n313), .ZN(new_n980));
  OAI21_X1  g794(.A(G900), .B1(new_n979), .B2(G227), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(G953), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n973), .A2(new_n980), .A3(new_n982), .ZN(G72));
  NAND2_X1  g797(.A1(G472), .A2(G902), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT63), .Z(new_n985));
  INV_X1    g799(.A(new_n876), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n985), .B1(new_n977), .B2(new_n986), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n303), .A2(new_n193), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n906), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n303), .A2(new_n304), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(new_n279), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n875), .A2(new_n879), .A3(new_n985), .A4(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n985), .B1(new_n968), .B2(new_n986), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n304), .B1(new_n283), .B2(new_n278), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n993), .B1(new_n994), .B2(new_n995), .ZN(G57));
endmodule


