

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584;

  XNOR2_X1 U320 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U321 ( .A(n315), .B(n400), .Z(n288) );
  XOR2_X1 U322 ( .A(n364), .B(KEYINPUT112), .Z(n289) );
  XOR2_X1 U323 ( .A(n329), .B(n328), .Z(n290) );
  INV_X1 U324 ( .A(KEYINPUT11), .ZN(n317) );
  NOR2_X1 U325 ( .A1(n411), .A2(n492), .ZN(n413) );
  XNOR2_X1 U326 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U327 ( .A(n303), .B(n437), .ZN(n304) );
  XNOR2_X1 U328 ( .A(n367), .B(n366), .ZN(n545) );
  XNOR2_X1 U329 ( .A(n305), .B(n304), .ZN(n307) );
  NAND2_X1 U330 ( .A1(n451), .A2(n497), .ZN(n452) );
  XNOR2_X1 U331 ( .A(n359), .B(KEYINPUT74), .ZN(n539) );
  XNOR2_X1 U332 ( .A(n456), .B(G190GAT), .ZN(n457) );
  XNOR2_X1 U333 ( .A(n458), .B(n457), .ZN(G1351GAT) );
  INV_X1 U334 ( .A(G92GAT), .ZN(n291) );
  NAND2_X1 U335 ( .A1(n291), .A2(G85GAT), .ZN(n294) );
  INV_X1 U336 ( .A(G85GAT), .ZN(n292) );
  NAND2_X1 U337 ( .A1(n292), .A2(G92GAT), .ZN(n293) );
  NAND2_X1 U338 ( .A1(n294), .A2(n293), .ZN(n296) );
  XNOR2_X1 U339 ( .A(G99GAT), .B(G106GAT), .ZN(n295) );
  XNOR2_X1 U340 ( .A(n296), .B(n295), .ZN(n315) );
  XNOR2_X1 U341 ( .A(n315), .B(KEYINPUT33), .ZN(n297) );
  XNOR2_X1 U342 ( .A(n297), .B(KEYINPUT31), .ZN(n300) );
  XOR2_X1 U343 ( .A(G176GAT), .B(G64GAT), .Z(n373) );
  XNOR2_X1 U344 ( .A(n373), .B(KEYINPUT70), .ZN(n298) );
  XOR2_X1 U345 ( .A(n298), .B(KEYINPUT32), .Z(n299) );
  XNOR2_X1 U346 ( .A(n300), .B(n299), .ZN(n305) );
  XNOR2_X1 U347 ( .A(G78GAT), .B(G204GAT), .ZN(n301) );
  XNOR2_X1 U348 ( .A(n301), .B(G148GAT), .ZN(n415) );
  XNOR2_X1 U349 ( .A(G57GAT), .B(KEYINPUT69), .ZN(n302) );
  XNOR2_X1 U350 ( .A(n302), .B(KEYINPUT13), .ZN(n351) );
  XNOR2_X1 U351 ( .A(n415), .B(n351), .ZN(n303) );
  XOR2_X1 U352 ( .A(G120GAT), .B(G71GAT), .Z(n437) );
  AND2_X1 U353 ( .A1(G230GAT), .A2(G233GAT), .ZN(n306) );
  XNOR2_X1 U354 ( .A(n307), .B(n306), .ZN(n575) );
  XNOR2_X1 U355 ( .A(KEYINPUT41), .B(n575), .ZN(n551) );
  XNOR2_X1 U356 ( .A(KEYINPUT105), .B(n551), .ZN(n532) );
  XNOR2_X1 U357 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n308) );
  XNOR2_X1 U358 ( .A(n308), .B(G29GAT), .ZN(n309) );
  XOR2_X1 U359 ( .A(n309), .B(KEYINPUT7), .Z(n311) );
  XNOR2_X1 U360 ( .A(G43GAT), .B(G50GAT), .ZN(n310) );
  XNOR2_X1 U361 ( .A(n311), .B(n310), .ZN(n332) );
  XOR2_X1 U362 ( .A(KEYINPUT71), .B(KEYINPUT72), .Z(n313) );
  XNOR2_X1 U363 ( .A(KEYINPUT10), .B(KEYINPUT9), .ZN(n312) );
  XNOR2_X1 U364 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U365 ( .A(n332), .B(n314), .ZN(n322) );
  XOR2_X1 U366 ( .A(G134GAT), .B(KEYINPUT73), .Z(n400) );
  NAND2_X1 U367 ( .A1(G232GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U368 ( .A(n288), .B(n316), .ZN(n320) );
  XOR2_X1 U369 ( .A(G218GAT), .B(G162GAT), .Z(n414) );
  XNOR2_X1 U370 ( .A(G190GAT), .B(n414), .ZN(n318) );
  XNOR2_X1 U371 ( .A(n322), .B(n321), .ZN(n560) );
  INV_X1 U372 ( .A(n560), .ZN(n359) );
  XNOR2_X1 U373 ( .A(G15GAT), .B(G1GAT), .ZN(n323) );
  XNOR2_X1 U374 ( .A(n323), .B(KEYINPUT66), .ZN(n343) );
  XOR2_X1 U375 ( .A(n343), .B(KEYINPUT29), .Z(n325) );
  NAND2_X1 U376 ( .A1(G229GAT), .A2(G233GAT), .ZN(n324) );
  XNOR2_X1 U377 ( .A(n325), .B(n324), .ZN(n329) );
  XOR2_X1 U378 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n327) );
  XNOR2_X1 U379 ( .A(G113GAT), .B(G197GAT), .ZN(n326) );
  XNOR2_X1 U380 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U381 ( .A(G141GAT), .B(G22GAT), .Z(n420) );
  XOR2_X1 U382 ( .A(G169GAT), .B(G8GAT), .Z(n383) );
  XNOR2_X1 U383 ( .A(n420), .B(n383), .ZN(n330) );
  XNOR2_X1 U384 ( .A(n290), .B(n330), .ZN(n331) );
  XOR2_X1 U385 ( .A(n332), .B(n331), .Z(n570) );
  NOR2_X1 U386 ( .A1(n570), .A2(n551), .ZN(n334) );
  XNOR2_X1 U387 ( .A(KEYINPUT111), .B(KEYINPUT46), .ZN(n333) );
  XNOR2_X1 U388 ( .A(n334), .B(n333), .ZN(n356) );
  XOR2_X1 U389 ( .A(KEYINPUT77), .B(KEYINPUT75), .Z(n336) );
  XNOR2_X1 U390 ( .A(G64GAT), .B(KEYINPUT76), .ZN(n335) );
  XNOR2_X1 U391 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U392 ( .A(G78GAT), .B(G155GAT), .Z(n338) );
  XNOR2_X1 U393 ( .A(G8GAT), .B(G211GAT), .ZN(n337) );
  XNOR2_X1 U394 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U395 ( .A(n340), .B(n339), .ZN(n355) );
  XOR2_X1 U396 ( .A(G71GAT), .B(G127GAT), .Z(n342) );
  XNOR2_X1 U397 ( .A(G22GAT), .B(G183GAT), .ZN(n341) );
  XNOR2_X1 U398 ( .A(n342), .B(n341), .ZN(n347) );
  XOR2_X1 U399 ( .A(n343), .B(KEYINPUT14), .Z(n345) );
  NAND2_X1 U400 ( .A1(G231GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U401 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U402 ( .A(n347), .B(n346), .Z(n353) );
  XOR2_X1 U403 ( .A(KEYINPUT79), .B(KEYINPUT12), .Z(n349) );
  XNOR2_X1 U404 ( .A(KEYINPUT15), .B(KEYINPUT78), .ZN(n348) );
  XNOR2_X1 U405 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U406 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U407 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U408 ( .A(n355), .B(n354), .ZN(n557) );
  NAND2_X1 U409 ( .A1(n356), .A2(n557), .ZN(n357) );
  NOR2_X1 U410 ( .A1(n359), .A2(n357), .ZN(n358) );
  XNOR2_X1 U411 ( .A(n358), .B(KEYINPUT47), .ZN(n365) );
  INV_X1 U412 ( .A(KEYINPUT36), .ZN(n360) );
  XNOR2_X1 U413 ( .A(n360), .B(n539), .ZN(n486) );
  NOR2_X1 U414 ( .A1(n486), .A2(n557), .ZN(n361) );
  XNOR2_X1 U415 ( .A(n361), .B(KEYINPUT45), .ZN(n363) );
  XNOR2_X1 U416 ( .A(n570), .B(KEYINPUT68), .ZN(n459) );
  INV_X1 U417 ( .A(n459), .ZN(n563) );
  NOR2_X1 U418 ( .A1(n575), .A2(n563), .ZN(n362) );
  AND2_X1 U419 ( .A1(n363), .A2(n362), .ZN(n364) );
  NAND2_X1 U420 ( .A1(n365), .A2(n289), .ZN(n367) );
  XNOR2_X1 U421 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n366) );
  XOR2_X1 U422 ( .A(G183GAT), .B(KEYINPUT19), .Z(n369) );
  XNOR2_X1 U423 ( .A(KEYINPUT17), .B(KEYINPUT84), .ZN(n368) );
  XNOR2_X1 U424 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U425 ( .A(n370), .B(KEYINPUT83), .Z(n372) );
  XNOR2_X1 U426 ( .A(KEYINPUT18), .B(G190GAT), .ZN(n371) );
  XNOR2_X1 U427 ( .A(n372), .B(n371), .ZN(n448) );
  XOR2_X1 U428 ( .A(n373), .B(KEYINPUT96), .Z(n375) );
  NAND2_X1 U429 ( .A1(G226GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U430 ( .A(n375), .B(n374), .ZN(n379) );
  XOR2_X1 U431 ( .A(G92GAT), .B(G204GAT), .Z(n377) );
  XNOR2_X1 U432 ( .A(G36GAT), .B(G218GAT), .ZN(n376) );
  XNOR2_X1 U433 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U434 ( .A(n379), .B(n378), .Z(n385) );
  XOR2_X1 U435 ( .A(KEYINPUT87), .B(KEYINPUT88), .Z(n381) );
  XNOR2_X1 U436 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n380) );
  XNOR2_X1 U437 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U438 ( .A(G197GAT), .B(n382), .Z(n430) );
  XNOR2_X1 U439 ( .A(n383), .B(n430), .ZN(n384) );
  XNOR2_X1 U440 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U441 ( .A(n448), .B(n386), .Z(n495) );
  NAND2_X1 U442 ( .A1(n545), .A2(n495), .ZN(n388) );
  XOR2_X1 U443 ( .A(KEYINPUT121), .B(KEYINPUT54), .Z(n387) );
  XNOR2_X1 U444 ( .A(n388), .B(n387), .ZN(n411) );
  XOR2_X1 U445 ( .A(KEYINPUT4), .B(KEYINPUT93), .Z(n390) );
  XNOR2_X1 U446 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n389) );
  XNOR2_X1 U447 ( .A(n390), .B(n389), .ZN(n410) );
  XOR2_X1 U448 ( .A(G148GAT), .B(G162GAT), .Z(n392) );
  XNOR2_X1 U449 ( .A(G141GAT), .B(G120GAT), .ZN(n391) );
  XNOR2_X1 U450 ( .A(n392), .B(n391), .ZN(n396) );
  XOR2_X1 U451 ( .A(KEYINPUT94), .B(KEYINPUT5), .Z(n394) );
  XNOR2_X1 U452 ( .A(G1GAT), .B(G57GAT), .ZN(n393) );
  XNOR2_X1 U453 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U454 ( .A(n396), .B(n395), .Z(n408) );
  XNOR2_X1 U455 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n397) );
  XNOR2_X1 U456 ( .A(n397), .B(G127GAT), .ZN(n440) );
  XOR2_X1 U457 ( .A(n440), .B(KEYINPUT95), .Z(n399) );
  NAND2_X1 U458 ( .A1(G225GAT), .A2(G233GAT), .ZN(n398) );
  XNOR2_X1 U459 ( .A(n399), .B(n398), .ZN(n406) );
  XOR2_X1 U460 ( .A(G85GAT), .B(n400), .Z(n404) );
  XOR2_X1 U461 ( .A(G155GAT), .B(KEYINPUT2), .Z(n402) );
  XNOR2_X1 U462 ( .A(KEYINPUT3), .B(KEYINPUT89), .ZN(n401) );
  XNOR2_X1 U463 ( .A(n402), .B(n401), .ZN(n416) );
  XNOR2_X1 U464 ( .A(G29GAT), .B(n416), .ZN(n403) );
  XNOR2_X1 U465 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U466 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U467 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U468 ( .A(n410), .B(n409), .ZN(n492) );
  INV_X1 U469 ( .A(KEYINPUT65), .ZN(n412) );
  XNOR2_X1 U470 ( .A(n413), .B(n412), .ZN(n568) );
  XOR2_X1 U471 ( .A(n415), .B(n414), .Z(n422) );
  XOR2_X1 U472 ( .A(n416), .B(KEYINPUT24), .Z(n418) );
  NAND2_X1 U473 ( .A1(G228GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U474 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U475 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U476 ( .A(n422), .B(n421), .ZN(n426) );
  XOR2_X1 U477 ( .A(KEYINPUT86), .B(KEYINPUT92), .Z(n424) );
  XNOR2_X1 U478 ( .A(G50GAT), .B(G106GAT), .ZN(n423) );
  XNOR2_X1 U479 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U480 ( .A(n426), .B(n425), .Z(n432) );
  XOR2_X1 U481 ( .A(KEYINPUT90), .B(KEYINPUT22), .Z(n428) );
  XNOR2_X1 U482 ( .A(KEYINPUT91), .B(KEYINPUT23), .ZN(n427) );
  XNOR2_X1 U483 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U484 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U485 ( .A(n432), .B(n431), .ZN(n469) );
  NAND2_X1 U486 ( .A1(n568), .A2(n469), .ZN(n433) );
  XNOR2_X1 U487 ( .A(n433), .B(KEYINPUT55), .ZN(n451) );
  XOR2_X1 U488 ( .A(KEYINPUT80), .B(KEYINPUT85), .Z(n435) );
  XNOR2_X1 U489 ( .A(G43GAT), .B(G134GAT), .ZN(n434) );
  XNOR2_X1 U490 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U491 ( .A(n436), .B(G99GAT), .Z(n439) );
  XNOR2_X1 U492 ( .A(G169GAT), .B(n437), .ZN(n438) );
  XNOR2_X1 U493 ( .A(n439), .B(n438), .ZN(n444) );
  XOR2_X1 U494 ( .A(G15GAT), .B(n440), .Z(n442) );
  NAND2_X1 U495 ( .A1(G227GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U496 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U497 ( .A(n444), .B(n443), .Z(n450) );
  XOR2_X1 U498 ( .A(G176GAT), .B(KEYINPUT81), .Z(n446) );
  XNOR2_X1 U499 ( .A(KEYINPUT20), .B(KEYINPUT82), .ZN(n445) );
  XNOR2_X1 U500 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U501 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U502 ( .A(n450), .B(n449), .ZN(n497) );
  XOR2_X2 U503 ( .A(n452), .B(KEYINPUT122), .Z(n565) );
  NAND2_X1 U504 ( .A1(n532), .A2(n565), .ZN(n455) );
  XOR2_X1 U505 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n453) );
  XNOR2_X1 U506 ( .A(n453), .B(G176GAT), .ZN(n454) );
  XNOR2_X1 U507 ( .A(n455), .B(n454), .ZN(G1349GAT) );
  NAND2_X1 U508 ( .A1(n539), .A2(n565), .ZN(n458) );
  XOR2_X1 U509 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n456) );
  INV_X1 U510 ( .A(n492), .ZN(n517) );
  NOR2_X1 U511 ( .A1(n575), .A2(n459), .ZN(n490) );
  NAND2_X1 U512 ( .A1(n497), .A2(n495), .ZN(n460) );
  XNOR2_X1 U513 ( .A(KEYINPUT100), .B(n460), .ZN(n461) );
  NAND2_X1 U514 ( .A1(n461), .A2(n469), .ZN(n462) );
  XOR2_X1 U515 ( .A(KEYINPUT25), .B(n462), .Z(n467) );
  XNOR2_X1 U516 ( .A(KEYINPUT99), .B(KEYINPUT26), .ZN(n464) );
  NOR2_X1 U517 ( .A1(n497), .A2(n469), .ZN(n463) );
  XNOR2_X1 U518 ( .A(n464), .B(n463), .ZN(n465) );
  XOR2_X1 U519 ( .A(KEYINPUT98), .B(n465), .Z(n567) );
  XNOR2_X1 U520 ( .A(n495), .B(KEYINPUT27), .ZN(n470) );
  NAND2_X1 U521 ( .A1(n567), .A2(n470), .ZN(n466) );
  NAND2_X1 U522 ( .A1(n467), .A2(n466), .ZN(n468) );
  NAND2_X1 U523 ( .A1(n517), .A2(n468), .ZN(n473) );
  XOR2_X1 U524 ( .A(n469), .B(KEYINPUT28), .Z(n501) );
  NAND2_X1 U525 ( .A1(n470), .A2(n492), .ZN(n471) );
  XOR2_X1 U526 ( .A(KEYINPUT97), .B(n471), .Z(n546) );
  NOR2_X1 U527 ( .A1(n501), .A2(n546), .ZN(n528) );
  INV_X1 U528 ( .A(n497), .ZN(n530) );
  NAND2_X1 U529 ( .A1(n528), .A2(n530), .ZN(n472) );
  NAND2_X1 U530 ( .A1(n473), .A2(n472), .ZN(n474) );
  XNOR2_X1 U531 ( .A(KEYINPUT101), .B(n474), .ZN(n487) );
  NOR2_X1 U532 ( .A1(n557), .A2(n539), .ZN(n475) );
  XOR2_X1 U533 ( .A(KEYINPUT16), .B(n475), .Z(n476) );
  NOR2_X1 U534 ( .A1(n487), .A2(n476), .ZN(n477) );
  XNOR2_X1 U535 ( .A(KEYINPUT102), .B(n477), .ZN(n504) );
  NAND2_X1 U536 ( .A1(n490), .A2(n504), .ZN(n484) );
  NOR2_X1 U537 ( .A1(n517), .A2(n484), .ZN(n478) );
  XOR2_X1 U538 ( .A(G1GAT), .B(n478), .Z(n479) );
  XNOR2_X1 U539 ( .A(KEYINPUT34), .B(n479), .ZN(G1324GAT) );
  INV_X1 U540 ( .A(n495), .ZN(n519) );
  NOR2_X1 U541 ( .A1(n519), .A2(n484), .ZN(n480) );
  XOR2_X1 U542 ( .A(G8GAT), .B(n480), .Z(G1325GAT) );
  NOR2_X1 U543 ( .A1(n530), .A2(n484), .ZN(n482) );
  XNOR2_X1 U544 ( .A(KEYINPUT103), .B(KEYINPUT35), .ZN(n481) );
  XNOR2_X1 U545 ( .A(n482), .B(n481), .ZN(n483) );
  XOR2_X1 U546 ( .A(G15GAT), .B(n483), .Z(G1326GAT) );
  INV_X1 U547 ( .A(n501), .ZN(n524) );
  NOR2_X1 U548 ( .A1(n524), .A2(n484), .ZN(n485) );
  XOR2_X1 U549 ( .A(G22GAT), .B(n485), .Z(G1327GAT) );
  XOR2_X1 U550 ( .A(G29GAT), .B(KEYINPUT39), .Z(n494) );
  NOR2_X1 U551 ( .A1(n486), .A2(n487), .ZN(n488) );
  NAND2_X1 U552 ( .A1(n557), .A2(n488), .ZN(n489) );
  XNOR2_X1 U553 ( .A(KEYINPUT37), .B(n489), .ZN(n516) );
  NAND2_X1 U554 ( .A1(n490), .A2(n516), .ZN(n491) );
  XOR2_X1 U555 ( .A(KEYINPUT38), .B(n491), .Z(n502) );
  NAND2_X1 U556 ( .A1(n502), .A2(n492), .ZN(n493) );
  XNOR2_X1 U557 ( .A(n494), .B(n493), .ZN(G1328GAT) );
  NAND2_X1 U558 ( .A1(n502), .A2(n495), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n496), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT104), .B(KEYINPUT40), .Z(n499) );
  NAND2_X1 U561 ( .A1(n497), .A2(n502), .ZN(n498) );
  XNOR2_X1 U562 ( .A(n499), .B(n498), .ZN(n500) );
  XOR2_X1 U563 ( .A(G43GAT), .B(n500), .Z(G1330GAT) );
  NAND2_X1 U564 ( .A1(n502), .A2(n501), .ZN(n503) );
  XNOR2_X1 U565 ( .A(n503), .B(G50GAT), .ZN(G1331GAT) );
  AND2_X1 U566 ( .A1(n570), .A2(n532), .ZN(n515) );
  NAND2_X1 U567 ( .A1(n515), .A2(n504), .ZN(n511) );
  NOR2_X1 U568 ( .A1(n517), .A2(n511), .ZN(n505) );
  XOR2_X1 U569 ( .A(KEYINPUT42), .B(n505), .Z(n506) );
  XNOR2_X1 U570 ( .A(G57GAT), .B(n506), .ZN(G1332GAT) );
  NOR2_X1 U571 ( .A1(n519), .A2(n511), .ZN(n508) );
  XNOR2_X1 U572 ( .A(KEYINPUT106), .B(KEYINPUT107), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U574 ( .A(G64GAT), .B(n509), .ZN(G1333GAT) );
  NOR2_X1 U575 ( .A1(n530), .A2(n511), .ZN(n510) );
  XOR2_X1 U576 ( .A(G71GAT), .B(n510), .Z(G1334GAT) );
  NOR2_X1 U577 ( .A1(n524), .A2(n511), .ZN(n513) );
  XNOR2_X1 U578 ( .A(KEYINPUT108), .B(KEYINPUT43), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U580 ( .A(G78GAT), .B(n514), .ZN(G1335GAT) );
  NAND2_X1 U581 ( .A1(n516), .A2(n515), .ZN(n523) );
  NOR2_X1 U582 ( .A1(n517), .A2(n523), .ZN(n518) );
  XOR2_X1 U583 ( .A(G85GAT), .B(n518), .Z(G1336GAT) );
  NOR2_X1 U584 ( .A1(n519), .A2(n523), .ZN(n521) );
  XNOR2_X1 U585 ( .A(G92GAT), .B(KEYINPUT109), .ZN(n520) );
  XNOR2_X1 U586 ( .A(n521), .B(n520), .ZN(G1337GAT) );
  NOR2_X1 U587 ( .A1(n530), .A2(n523), .ZN(n522) );
  XOR2_X1 U588 ( .A(G99GAT), .B(n522), .Z(G1338GAT) );
  NOR2_X1 U589 ( .A1(n524), .A2(n523), .ZN(n526) );
  XNOR2_X1 U590 ( .A(KEYINPUT44), .B(KEYINPUT110), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n526), .B(n525), .ZN(n527) );
  XOR2_X1 U592 ( .A(G106GAT), .B(n527), .Z(G1339GAT) );
  NAND2_X1 U593 ( .A1(n528), .A2(n545), .ZN(n529) );
  NOR2_X1 U594 ( .A1(n530), .A2(n529), .ZN(n540) );
  NAND2_X1 U595 ( .A1(n540), .A2(n563), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n531), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT49), .B(KEYINPUT114), .Z(n534) );
  NAND2_X1 U598 ( .A1(n540), .A2(n532), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n534), .B(n533), .ZN(n536) );
  XOR2_X1 U600 ( .A(G120GAT), .B(KEYINPUT113), .Z(n535) );
  XNOR2_X1 U601 ( .A(n536), .B(n535), .ZN(G1341GAT) );
  INV_X1 U602 ( .A(n557), .ZN(n578) );
  NAND2_X1 U603 ( .A1(n578), .A2(n540), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n537), .B(KEYINPUT50), .ZN(n538) );
  XNOR2_X1 U605 ( .A(G127GAT), .B(n538), .ZN(G1342GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n542) );
  NAND2_X1 U607 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U608 ( .A(n542), .B(n541), .ZN(n544) );
  XOR2_X1 U609 ( .A(G134GAT), .B(KEYINPUT116), .Z(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(G1343GAT) );
  INV_X1 U611 ( .A(n545), .ZN(n547) );
  NOR2_X1 U612 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U613 ( .A1(n567), .A2(n548), .ZN(n559) );
  NOR2_X1 U614 ( .A1(n570), .A2(n559), .ZN(n550) );
  XNOR2_X1 U615 ( .A(G141GAT), .B(KEYINPUT117), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(G1344GAT) );
  NOR2_X1 U617 ( .A1(n551), .A2(n559), .ZN(n556) );
  XOR2_X1 U618 ( .A(KEYINPUT119), .B(KEYINPUT53), .Z(n553) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U621 ( .A(KEYINPUT118), .B(n554), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(G1345GAT) );
  NOR2_X1 U623 ( .A1(n557), .A2(n559), .ZN(n558) );
  XOR2_X1 U624 ( .A(G155GAT), .B(n558), .Z(G1346GAT) );
  NOR2_X1 U625 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U626 ( .A(KEYINPUT120), .B(n561), .Z(n562) );
  XNOR2_X1 U627 ( .A(G162GAT), .B(n562), .ZN(G1347GAT) );
  NAND2_X1 U628 ( .A1(n565), .A2(n563), .ZN(n564) );
  XNOR2_X1 U629 ( .A(n564), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U630 ( .A1(n565), .A2(n578), .ZN(n566) );
  XNOR2_X1 U631 ( .A(n566), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U632 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U633 ( .A(KEYINPUT124), .B(n569), .ZN(n581) );
  NOR2_X1 U634 ( .A1(n581), .A2(n570), .ZN(n574) );
  XOR2_X1 U635 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n572) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  XOR2_X1 U639 ( .A(G204GAT), .B(KEYINPUT61), .Z(n577) );
  INV_X1 U640 ( .A(n581), .ZN(n579) );
  NAND2_X1 U641 ( .A1(n575), .A2(n579), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  NAND2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U644 ( .A(n580), .B(G211GAT), .ZN(G1354GAT) );
  XNOR2_X1 U645 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n583) );
  NOR2_X1 U646 ( .A1(n486), .A2(n581), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(n584) );
  XOR2_X1 U648 ( .A(G218GAT), .B(n584), .Z(G1355GAT) );
endmodule

