//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 0 0 1 1 0 0 0 0 1 0 0 0 1 0 1 0 1 1 0 0 1 0 1 0 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 1 1 0 0 0 0 0 1 1 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:26 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1227, new_n1228, new_n1229, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n203), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n209), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n220), .B1(new_n202), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n211), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n214), .B(new_n219), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G226), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  INV_X1    g0039(.A(G50), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n240), .A2(G68), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n202), .A2(G50), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT66), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT65), .ZN(new_n248));
  XOR2_X1   g0048(.A(G107), .B(G116), .Z(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n246), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(KEYINPUT68), .ZN(new_n252));
  AND2_X1   g0052(.A1(KEYINPUT67), .A2(G45), .ZN(new_n253));
  NOR2_X1   g0053(.A1(KEYINPUT67), .A2(G45), .ZN(new_n254));
  NOR3_X1   g0054(.A1(new_n253), .A2(new_n254), .A3(G41), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n252), .B1(new_n255), .B2(G1), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n257));
  INV_X1    g0057(.A(G274), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT67), .B(G45), .ZN(new_n260));
  OAI211_X1 g0060(.A(KEYINPUT68), .B(new_n208), .C1(new_n260), .C2(G41), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n256), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  INV_X1    g0063(.A(G41), .ZN(new_n264));
  OAI211_X1 g0064(.A(G1), .B(G13), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G226), .ZN(new_n269));
  AND2_X1   g0069(.A1(new_n262), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT3), .B(G33), .ZN(new_n271));
  INV_X1    g0071(.A(G1698), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n271), .A2(G222), .A3(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n271), .A2(G223), .A3(G1698), .ZN(new_n274));
  INV_X1    g0074(.A(G77), .ZN(new_n275));
  OAI211_X1 g0075(.A(new_n273), .B(new_n274), .C1(new_n275), .C2(new_n271), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n257), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n270), .A2(G190), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n277), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n262), .A2(new_n269), .ZN(new_n280));
  OAI21_X1  g0080(.A(G200), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n282));
  INV_X1    g0082(.A(G150), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n209), .A2(new_n263), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT8), .B(G58), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n209), .A2(G33), .ZN(new_n286));
  OAI221_X1 g0086(.A(new_n282), .B1(new_n283), .B2(new_n284), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n217), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n287), .A2(new_n289), .B1(new_n240), .B2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT9), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT70), .ZN(new_n294));
  OAI21_X1  g0094(.A(KEYINPUT69), .B1(new_n209), .B2(G1), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT69), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n296), .A2(new_n208), .A3(G20), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n294), .B1(new_n299), .B2(new_n240), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n290), .A2(new_n217), .A3(new_n288), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n298), .A2(KEYINPUT70), .A3(G50), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n300), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  AND3_X1   g0104(.A1(new_n292), .A2(new_n293), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n293), .B1(new_n292), .B2(new_n304), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n278), .B(new_n281), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT10), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n308), .B1(new_n281), .B2(KEYINPUT72), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n307), .A2(new_n309), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n291), .A2(new_n202), .ZN(new_n314));
  XNOR2_X1  g0114(.A(new_n314), .B(KEYINPUT12), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT73), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n302), .A2(G68), .A3(new_n298), .ZN(new_n317));
  AND3_X1   g0117(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n316), .B1(new_n315), .B2(new_n317), .ZN(new_n319));
  OAI22_X1  g0119(.A1(new_n284), .A2(new_n240), .B1(new_n209), .B2(G68), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n286), .A2(new_n275), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n289), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT11), .ZN(new_n323));
  XNOR2_X1  g0123(.A(new_n322), .B(new_n323), .ZN(new_n324));
  NOR3_X1   g0124(.A1(new_n318), .A2(new_n319), .A3(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT14), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT13), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n267), .A2(new_n221), .ZN(new_n329));
  AND2_X1   g0129(.A1(new_n261), .A2(new_n259), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n329), .B1(new_n330), .B2(new_n256), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n271), .A2(G232), .A3(G1698), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n271), .A2(G226), .A3(new_n272), .ZN(new_n333));
  NAND2_X1  g0133(.A1(G33), .A2(G97), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n257), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n328), .B1(new_n331), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n329), .ZN(new_n338));
  AND4_X1   g0138(.A1(new_n328), .A2(new_n336), .A3(new_n262), .A4(new_n338), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n327), .B(G169), .C1(new_n337), .C2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n331), .A2(new_n328), .A3(new_n336), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n262), .A2(new_n338), .ZN(new_n342));
  AND2_X1   g0142(.A1(new_n335), .A2(new_n257), .ZN(new_n343));
  OAI21_X1  g0143(.A(KEYINPUT13), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n341), .A2(new_n344), .A3(G179), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n340), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n341), .A2(new_n344), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n327), .B1(new_n347), .B2(G169), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n326), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(G190), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n325), .B1(new_n347), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(G200), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n352), .B1(new_n341), .B2(new_n344), .ZN(new_n353));
  OR2_X1    g0153(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n270), .A2(new_n277), .ZN(new_n355));
  INV_X1    g0155(.A(G169), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n292), .A2(new_n304), .ZN(new_n358));
  XNOR2_X1  g0158(.A(KEYINPUT71), .B(G179), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n357), .B(new_n358), .C1(new_n360), .C2(new_n355), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n271), .A2(G232), .A3(new_n272), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n271), .A2(G238), .A3(G1698), .ZN(new_n363));
  INV_X1    g0163(.A(G107), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n362), .B(new_n363), .C1(new_n364), .C2(new_n271), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n257), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n268), .A2(G244), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n366), .A2(new_n262), .A3(new_n367), .ZN(new_n368));
  OR2_X1    g0168(.A1(new_n368), .A2(new_n360), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n356), .ZN(new_n370));
  NOR3_X1   g0170(.A1(new_n299), .A2(new_n275), .A3(new_n301), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n371), .B1(new_n275), .B2(new_n291), .ZN(new_n372));
  OAI22_X1  g0172(.A1(new_n285), .A2(new_n284), .B1(new_n209), .B2(new_n275), .ZN(new_n373));
  XNOR2_X1  g0173(.A(KEYINPUT15), .B(G87), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n374), .A2(new_n286), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n289), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n372), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n369), .A2(new_n370), .A3(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n377), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n368), .A2(G200), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n379), .B(new_n380), .C1(new_n350), .C2(new_n368), .ZN(new_n381));
  AND3_X1   g0181(.A1(new_n361), .A2(new_n378), .A3(new_n381), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n313), .A2(new_n349), .A3(new_n354), .A4(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT77), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT17), .ZN(new_n386));
  AND3_X1   g0186(.A1(new_n265), .A2(G232), .A3(new_n266), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT3), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(G33), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n388), .A2(new_n390), .A3(G226), .A4(G1698), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n388), .A2(new_n390), .A3(G223), .A4(new_n272), .ZN(new_n392));
  NAND2_X1  g0192(.A1(G33), .A2(G87), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n387), .B1(new_n394), .B2(new_n257), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n262), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n352), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n395), .A2(new_n262), .A3(new_n350), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n299), .A2(new_n285), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n400), .A2(new_n302), .B1(new_n291), .B2(new_n285), .ZN(new_n401));
  NAND2_X1  g0201(.A1(G58), .A2(G68), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n209), .B1(new_n203), .B2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(G159), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n284), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(KEYINPUT74), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  AND2_X1   g0206(.A1(G58), .A2(G68), .ZN(new_n407));
  NOR2_X1   g0207(.A1(G58), .A2(G68), .ZN(new_n408));
  OAI21_X1  g0208(.A(G20), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT74), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n409), .B(new_n410), .C1(new_n404), .C2(new_n284), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n406), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT7), .ZN(new_n413));
  NOR3_X1   g0213(.A1(new_n271), .A2(new_n413), .A3(G20), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n388), .A2(new_n390), .ZN(new_n415));
  AOI21_X1  g0215(.A(KEYINPUT7), .B1(new_n415), .B2(new_n209), .ZN(new_n416));
  OAI21_X1  g0216(.A(G68), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n412), .B1(new_n417), .B2(KEYINPUT75), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n413), .B1(new_n271), .B2(G20), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n415), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n202), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT75), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(KEYINPUT16), .B1(new_n418), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n417), .A2(new_n411), .A3(new_n406), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT16), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n289), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n399), .B(new_n401), .C1(new_n424), .C2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT76), .ZN(new_n429));
  INV_X1    g0229(.A(new_n401), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n411), .B(new_n406), .C1(new_n421), .C2(new_n422), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n417), .A2(KEYINPUT75), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n426), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n412), .A2(new_n421), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n434), .A2(KEYINPUT16), .B1(new_n217), .B2(new_n288), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n430), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT76), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n436), .A2(new_n437), .A3(new_n399), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n386), .B1(new_n429), .B2(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n396), .A2(new_n359), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n440), .B1(G169), .B2(new_n396), .ZN(new_n441));
  OAI21_X1  g0241(.A(KEYINPUT18), .B1(new_n436), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n401), .B1(new_n424), .B2(new_n427), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT18), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n396), .A2(G169), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n445), .B1(new_n359), .B2(new_n396), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n443), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n442), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n428), .A2(new_n386), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NOR3_X1   g0250(.A1(new_n439), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n384), .A2(new_n385), .A3(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n428), .A2(KEYINPUT76), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n437), .B1(new_n436), .B2(new_n399), .ZN(new_n454));
  OAI21_X1  g0254(.A(KEYINPUT17), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AND2_X1   g0255(.A1(new_n442), .A2(new_n447), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n455), .A2(new_n456), .A3(new_n449), .ZN(new_n457));
  OAI21_X1  g0257(.A(KEYINPUT77), .B1(new_n383), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n452), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT82), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n264), .A2(KEYINPUT5), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n208), .A2(G45), .ZN(new_n462));
  OAI21_X1  g0262(.A(KEYINPUT79), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT80), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT5), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n464), .B1(new_n465), .B2(G41), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n264), .A2(KEYINPUT80), .A3(KEYINPUT5), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n465), .A2(G41), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT79), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n469), .A2(new_n470), .A3(new_n208), .A4(G45), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n463), .A2(new_n468), .A3(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n472), .A2(G257), .A3(new_n265), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n259), .A2(new_n468), .A3(new_n471), .A4(new_n463), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT81), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n473), .A2(KEYINPUT81), .A3(new_n474), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n271), .A2(G244), .A3(new_n272), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT4), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n271), .A2(KEYINPUT4), .A3(G244), .A4(new_n272), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n271), .A2(G250), .A3(G1698), .ZN(new_n483));
  NAND2_X1  g0283(.A1(G33), .A2(G283), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n481), .A2(new_n482), .A3(new_n483), .A4(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(new_n257), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n477), .A2(G190), .A3(new_n478), .A4(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(G97), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n291), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n208), .A2(G33), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n290), .A2(new_n490), .A3(new_n217), .A4(new_n288), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n489), .B1(new_n491), .B2(new_n488), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n284), .A2(new_n275), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT6), .ZN(new_n495));
  AND2_X1   g0295(.A1(G97), .A2(G107), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n495), .B1(new_n496), .B2(new_n205), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n364), .A2(KEYINPUT6), .A3(G97), .ZN(new_n498));
  AND2_X1   g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI211_X1 g0299(.A(KEYINPUT78), .B(new_n494), .C1(new_n499), .C2(new_n209), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT78), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n209), .B1(new_n497), .B2(new_n498), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n501), .B1(new_n502), .B2(new_n493), .ZN(new_n503));
  OAI21_X1  g0303(.A(G107), .B1(new_n414), .B2(new_n416), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n500), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n492), .B1(new_n505), .B2(new_n289), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n487), .A2(new_n506), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n475), .A2(new_n476), .B1(new_n485), .B2(new_n257), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n352), .B1(new_n508), .B2(new_n478), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n460), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n477), .A2(new_n478), .A3(new_n486), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(G200), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n512), .A2(KEYINPUT82), .A3(new_n506), .A4(new_n487), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n508), .A2(new_n359), .A3(new_n478), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n506), .B1(new_n511), .B2(new_n356), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n510), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n271), .A2(G244), .A3(G1698), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n388), .A2(new_n390), .A3(G238), .A4(new_n272), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G33), .A2(G116), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n257), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n462), .A2(new_n223), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n208), .A2(new_n258), .A3(G45), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n265), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n521), .A2(G190), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(KEYINPUT83), .ZN(new_n526));
  INV_X1    g0326(.A(new_n524), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n527), .B1(new_n520), .B2(new_n257), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT83), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n528), .A2(new_n529), .A3(G190), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n271), .A2(new_n209), .A3(G68), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT19), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n209), .B1(new_n334), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(G87), .B2(new_n206), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n533), .B1(new_n286), .B2(new_n488), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n532), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n537), .A2(new_n289), .B1(new_n291), .B2(new_n374), .ZN(new_n538));
  INV_X1    g0338(.A(new_n491), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(G87), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n538), .B(new_n540), .C1(new_n528), .C2(new_n352), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n528), .ZN(new_n543));
  INV_X1    g0343(.A(new_n374), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n539), .A2(new_n544), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n543), .A2(new_n356), .B1(new_n538), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n528), .A2(new_n359), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n531), .A2(new_n542), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n290), .A2(G116), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n549), .B1(new_n539), .B2(G116), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(G116), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n288), .A2(new_n217), .B1(G20), .B2(new_n552), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n484), .B(new_n209), .C1(G33), .C2(new_n488), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n553), .A2(KEYINPUT20), .A3(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(KEYINPUT20), .B1(new_n553), .B2(new_n554), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n551), .A2(new_n558), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n388), .A2(new_n390), .A3(G264), .A4(G1698), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n388), .A2(new_n390), .A3(G257), .A4(new_n272), .ZN(new_n561));
  INV_X1    g0361(.A(G303), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n560), .B(new_n561), .C1(new_n562), .C2(new_n271), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n257), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n472), .A2(G270), .A3(new_n265), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n564), .A2(new_n565), .A3(new_n474), .ZN(new_n566));
  INV_X1    g0366(.A(G179), .ZN(new_n567));
  NOR3_X1   g0367(.A1(new_n559), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(G169), .B1(new_n551), .B2(new_n558), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n564), .A2(new_n565), .A3(new_n474), .ZN(new_n570));
  OAI21_X1  g0370(.A(KEYINPUT21), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  OR2_X1    g0371(.A1(new_n556), .A2(new_n557), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n356), .B1(new_n572), .B2(new_n550), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT21), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n573), .A2(new_n566), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n568), .B1(new_n571), .B2(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n388), .A2(new_n390), .A3(G257), .A4(G1698), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n388), .A2(new_n390), .A3(G250), .A4(new_n272), .ZN(new_n578));
  NAND2_X1  g0378(.A1(G33), .A2(G294), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT85), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n577), .A2(new_n578), .A3(KEYINPUT85), .A4(new_n579), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n582), .A2(new_n257), .A3(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n472), .A2(G264), .A3(new_n265), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n584), .A2(new_n567), .A3(new_n474), .A4(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n584), .A2(new_n474), .A3(new_n585), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n356), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n222), .A2(KEYINPUT84), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n589), .A2(new_n388), .A3(new_n390), .A4(new_n209), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT22), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n271), .A2(KEYINPUT22), .A3(new_n209), .A4(new_n589), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n519), .A2(G20), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT23), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(new_n209), .B2(G107), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n364), .A2(KEYINPUT23), .A3(G20), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n594), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n592), .A2(new_n593), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(KEYINPUT24), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT24), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n592), .A2(new_n593), .A3(new_n598), .A4(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n603), .A2(new_n289), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n291), .A2(KEYINPUT25), .A3(new_n364), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT25), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(new_n290), .B2(G107), .ZN(new_n607));
  AOI22_X1  g0407(.A1(G107), .A2(new_n539), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n586), .B(new_n588), .C1(new_n604), .C2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n587), .A2(G200), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n609), .B1(new_n603), .B2(new_n289), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n584), .A2(G190), .A3(new_n474), .A4(new_n585), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n566), .A2(G200), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n615), .B(new_n559), .C1(new_n350), .C2(new_n566), .ZN(new_n616));
  AND4_X1   g0416(.A1(new_n576), .A2(new_n610), .A3(new_n614), .A4(new_n616), .ZN(new_n617));
  AND4_X1   g0417(.A1(new_n459), .A2(new_n516), .A3(new_n548), .A4(new_n617), .ZN(G372));
  NAND2_X1  g0418(.A1(new_n429), .A2(new_n438), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n450), .B1(new_n619), .B2(KEYINPUT17), .ZN(new_n620));
  INV_X1    g0420(.A(new_n378), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(new_n351), .B2(new_n353), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n349), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n448), .B1(new_n620), .B2(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(KEYINPUT86), .B1(new_n311), .B2(new_n312), .ZN(new_n625));
  INV_X1    g0425(.A(new_n312), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT86), .ZN(new_n627));
  NOR3_X1   g0427(.A1(new_n626), .A2(new_n310), .A3(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n361), .B1(new_n624), .B2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT87), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  OAI211_X1 g0432(.A(KEYINPUT87), .B(new_n361), .C1(new_n624), .C2(new_n629), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n510), .A2(new_n513), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n612), .A2(new_n613), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n576), .A2(new_n610), .B1(new_n636), .B2(new_n611), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n511), .A2(new_n356), .ZN(new_n638));
  INV_X1    g0438(.A(new_n506), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n638), .A2(new_n514), .A3(new_n639), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n635), .A2(new_n637), .A3(new_n640), .A4(new_n548), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n543), .A2(new_n356), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n538), .A2(new_n545), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n642), .A2(new_n547), .A3(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT26), .ZN(new_n646));
  AND4_X1   g0446(.A1(new_n529), .A2(new_n521), .A3(G190), .A4(new_n524), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n529), .B1(new_n528), .B2(G190), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n644), .B1(new_n649), .B2(new_n541), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n646), .B1(new_n640), .B2(new_n650), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n548), .A2(new_n515), .A3(KEYINPUT26), .A4(new_n514), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n645), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n641), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n459), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n634), .A2(new_n655), .ZN(G369));
  NAND3_X1  g0456(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n657), .A2(KEYINPUT27), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(KEYINPUT27), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(G213), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n660), .B(KEYINPUT88), .ZN(new_n661));
  INV_X1    g0461(.A(G343), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n664), .A2(new_n559), .ZN(new_n665));
  XOR2_X1   g0465(.A(new_n576), .B(new_n665), .Z(new_n666));
  AND2_X1   g0466(.A1(new_n666), .A2(new_n616), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(G330), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n614), .B1(new_n612), .B2(new_n664), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n610), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n610), .A2(new_n663), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n576), .A2(new_n663), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(new_n671), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n677), .B(KEYINPUT89), .ZN(G399));
  INV_X1    g0478(.A(new_n212), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n679), .A2(G41), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NOR3_X1   g0481(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(G1), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n215), .B2(new_n681), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n684), .B(KEYINPUT28), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n654), .A2(new_n664), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT90), .ZN(new_n687));
  AOI21_X1  g0487(.A(KEYINPUT29), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n663), .B1(new_n641), .B2(new_n653), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT29), .ZN(new_n690));
  NOR3_X1   g0490(.A1(new_n689), .A2(KEYINPUT90), .A3(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(G330), .ZN(new_n693));
  AND3_X1   g0493(.A1(new_n477), .A2(new_n478), .A3(new_n486), .ZN(new_n694));
  NOR3_X1   g0494(.A1(new_n543), .A2(new_n566), .A3(new_n567), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n584), .A2(new_n585), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n694), .A2(new_n695), .A3(KEYINPUT30), .A4(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT30), .ZN(new_n698));
  AOI211_X1 g0498(.A(new_n567), .B(new_n527), .C1(new_n520), .C2(new_n257), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n570), .A2(new_n699), .A3(new_n585), .A4(new_n584), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n698), .B1(new_n700), .B2(new_n511), .ZN(new_n701));
  NOR3_X1   g0501(.A1(new_n570), .A2(new_n360), .A3(new_n528), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n702), .A2(new_n511), .A3(new_n587), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n697), .A2(new_n701), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n663), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT31), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n704), .A2(KEYINPUT31), .A3(new_n663), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n516), .A2(new_n548), .A3(new_n617), .A4(new_n664), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n693), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n692), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n685), .B1(new_n714), .B2(G1), .ZN(G364));
  AND2_X1   g0515(.A1(new_n209), .A2(G13), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n208), .B1(new_n716), .B2(G45), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n680), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n668), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n667), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n721), .B1(new_n693), .B2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(G13), .A2(G33), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(G20), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n722), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n217), .B1(G20), .B2(new_n356), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n209), .A2(G190), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n352), .A2(G179), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(G179), .A2(G200), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n730), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AOI22_X1  g0536(.A1(G283), .A2(new_n733), .B1(new_n736), .B2(G329), .ZN(new_n737));
  INV_X1    g0537(.A(G322), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n359), .A2(G200), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n209), .A2(new_n350), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n737), .B1(new_n738), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n740), .A2(new_n731), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n415), .B1(new_n743), .B2(new_n562), .ZN(new_n744));
  XOR2_X1   g0544(.A(new_n744), .B(KEYINPUT98), .Z(new_n745));
  NOR3_X1   g0545(.A1(new_n359), .A2(new_n209), .A3(new_n352), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(new_n350), .ZN(new_n747));
  XOR2_X1   g0547(.A(KEYINPUT33), .B(G317), .Z(new_n748));
  OAI21_X1  g0548(.A(new_n745), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  AND3_X1   g0549(.A1(new_n739), .A2(KEYINPUT93), .A3(new_n730), .ZN(new_n750));
  AOI21_X1  g0550(.A(KEYINPUT93), .B1(new_n739), .B2(new_n730), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  AOI211_X1 g0553(.A(new_n742), .B(new_n749), .C1(G311), .C2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT94), .ZN(new_n755));
  AND3_X1   g0555(.A1(new_n746), .A2(new_n755), .A3(G190), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n755), .B1(new_n746), .B2(G190), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n209), .B1(new_n734), .B2(G190), .ZN(new_n760));
  XOR2_X1   g0560(.A(new_n760), .B(KEYINPUT95), .Z(new_n761));
  AOI22_X1  g0561(.A1(new_n759), .A2(G326), .B1(G294), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(KEYINPUT97), .ZN(new_n763));
  OR2_X1    g0563(.A1(new_n762), .A2(KEYINPUT97), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n754), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  XOR2_X1   g0565(.A(new_n761), .B(KEYINPUT96), .Z(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G97), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n759), .A2(G50), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n753), .A2(G77), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n736), .A2(G159), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(KEYINPUT32), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n747), .A2(new_n202), .B1(new_n741), .B2(new_n201), .ZN(new_n772));
  INV_X1    g0572(.A(new_n743), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G87), .ZN(new_n774));
  OAI211_X1 g0574(.A(new_n774), .B(new_n271), .C1(new_n364), .C2(new_n732), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n771), .A2(new_n772), .A3(new_n775), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n767), .A2(new_n768), .A3(new_n769), .A4(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n729), .B1(new_n765), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n726), .A2(new_n728), .ZN(new_n779));
  XOR2_X1   g0579(.A(new_n779), .B(KEYINPUT92), .Z(new_n780));
  NOR2_X1   g0580(.A1(new_n679), .A2(new_n271), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(new_n215), .B2(new_n260), .ZN(new_n782));
  INV_X1    g0582(.A(G45), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n245), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n679), .A2(new_n415), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G355), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n787), .B1(G116), .B2(new_n212), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n785), .B1(KEYINPUT91), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n789), .B1(KEYINPUT91), .B2(new_n788), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n720), .B(new_n778), .C1(new_n780), .C2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n723), .B1(new_n727), .B2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(G396));
  NOR2_X1   g0593(.A1(new_n728), .A2(new_n724), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n719), .B1(G77), .B2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n747), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n759), .A2(G137), .B1(G150), .B2(new_n797), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n798), .B(KEYINPUT99), .ZN(new_n799));
  INV_X1    g0599(.A(G143), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n799), .B1(new_n800), .B2(new_n741), .C1(new_n404), .C2(new_n752), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT34), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n415), .B1(new_n773), .B2(G50), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n733), .A2(G68), .ZN(new_n804));
  INV_X1    g0604(.A(G132), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n803), .B(new_n804), .C1(new_n805), .C2(new_n735), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(G58), .B2(new_n761), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n802), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n759), .A2(G303), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n753), .A2(G116), .ZN(new_n810));
  AOI22_X1  g0610(.A1(G107), .A2(new_n773), .B1(new_n733), .B2(G87), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n271), .B1(new_n736), .B2(G311), .ZN(new_n812));
  INV_X1    g0612(.A(G294), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n811), .B(new_n812), .C1(new_n813), .C2(new_n741), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(G283), .B2(new_n797), .ZN(new_n815));
  NAND4_X1  g0615(.A1(new_n767), .A2(new_n809), .A3(new_n810), .A4(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n808), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n796), .B1(new_n817), .B2(new_n728), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n378), .A2(new_n663), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n663), .A2(new_n377), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n381), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(new_n378), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n818), .A2(KEYINPUT100), .B1(new_n724), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(KEYINPUT100), .B2(new_n818), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n686), .A2(new_n824), .ZN(new_n827));
  INV_X1    g0627(.A(new_n824), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n689), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n719), .B1(new_n830), .B2(new_n712), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n712), .B2(new_n830), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n826), .A2(new_n832), .ZN(G384));
  INV_X1    g0633(.A(KEYINPUT38), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n434), .A2(KEYINPUT16), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n401), .B1(new_n427), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n661), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n838), .B1(new_n620), .B2(new_n456), .ZN(new_n839));
  AOI21_X1  g0639(.A(KEYINPUT37), .B1(new_n443), .B2(new_n446), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n443), .A2(new_n837), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n619), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n836), .B1(new_n446), .B2(new_n837), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n429), .A2(new_n438), .A3(new_n844), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n842), .A2(new_n843), .B1(new_n845), .B2(KEYINPUT37), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n834), .B1(new_n839), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n845), .A2(KEYINPUT37), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n840), .A2(new_n429), .A3(new_n438), .A4(new_n841), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n850), .B(KEYINPUT38), .C1(new_n451), .C2(new_n838), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n847), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n710), .A2(new_n707), .A3(new_n708), .ZN(new_n853));
  OAI21_X1  g0653(.A(G169), .B1(new_n337), .B2(new_n339), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(KEYINPUT14), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n855), .A2(new_n345), .A3(new_n340), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n351), .A2(new_n353), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n326), .B(new_n663), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n326), .A2(new_n663), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n349), .A2(new_n354), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n824), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  AND2_X1   g0661(.A1(new_n853), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n852), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT40), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n841), .B1(new_n620), .B2(new_n456), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n443), .A2(new_n446), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n866), .A2(new_n841), .A3(new_n428), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(KEYINPUT37), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n868), .A2(new_n849), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n834), .B1(new_n865), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n864), .B1(new_n870), .B2(new_n851), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n863), .A2(new_n864), .B1(new_n871), .B2(new_n862), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n459), .A2(new_n853), .ZN(new_n874));
  OAI21_X1  g0674(.A(G330), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n875), .B1(new_n874), .B2(new_n873), .ZN(new_n876));
  INV_X1    g0676(.A(new_n841), .ZN(new_n877));
  AOI22_X1  g0677(.A1(new_n457), .A2(new_n877), .B1(new_n849), .B2(new_n868), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n851), .B1(new_n878), .B2(KEYINPUT38), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT39), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n856), .A2(new_n326), .A3(new_n664), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n847), .A2(KEYINPUT39), .A3(new_n851), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n881), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n858), .A2(new_n860), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n887), .B1(new_n829), .B2(new_n820), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n888), .A2(new_n852), .B1(new_n448), .B2(new_n661), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n885), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n459), .B1(new_n688), .B2(new_n691), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n634), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n890), .B(new_n892), .ZN(new_n893));
  OAI22_X1  g0693(.A1(new_n876), .A2(new_n893), .B1(new_n208), .B2(new_n716), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n894), .B1(new_n893), .B2(new_n876), .ZN(new_n895));
  INV_X1    g0695(.A(new_n499), .ZN(new_n896));
  OR2_X1    g0696(.A1(new_n896), .A2(KEYINPUT35), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(KEYINPUT35), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n897), .A2(G116), .A3(new_n218), .A4(new_n898), .ZN(new_n899));
  XOR2_X1   g0699(.A(new_n899), .B(KEYINPUT36), .Z(new_n900));
  NAND3_X1  g0700(.A1(new_n216), .A2(G77), .A3(new_n402), .ZN(new_n901));
  AOI211_X1 g0701(.A(new_n208), .B(G13), .C1(new_n901), .C2(new_n241), .ZN(new_n902));
  OR3_X1    g0702(.A1(new_n895), .A2(new_n900), .A3(new_n902), .ZN(G367));
  NOR2_X1   g0703(.A1(new_n640), .A2(new_n664), .ZN(new_n904));
  XOR2_X1   g0704(.A(new_n904), .B(KEYINPUT101), .Z(new_n905));
  OAI21_X1  g0705(.A(new_n516), .B1(new_n506), .B2(new_n664), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n640), .B1(new_n907), .B2(new_n610), .ZN(new_n908));
  OR2_X1    g0708(.A1(new_n908), .A2(KEYINPUT102), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(KEYINPUT102), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n909), .A2(new_n664), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n538), .A2(new_n540), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n663), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n548), .A2(new_n913), .ZN(new_n914));
  OR2_X1    g0714(.A1(new_n913), .A2(new_n644), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n916), .A2(KEYINPUT43), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n907), .A2(new_n675), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n918), .B(KEYINPUT42), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n911), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(KEYINPUT103), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT103), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n911), .A2(new_n922), .A3(new_n917), .A4(new_n919), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n911), .A2(new_n919), .ZN(new_n925));
  XOR2_X1   g0725(.A(new_n916), .B(KEYINPUT43), .Z(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n905), .A2(new_n906), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n673), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n924), .A2(new_n673), .A3(new_n929), .A4(new_n927), .ZN(new_n932));
  XOR2_X1   g0732(.A(new_n680), .B(KEYINPUT41), .Z(new_n933));
  XNOR2_X1  g0733(.A(KEYINPUT105), .B(KEYINPUT44), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n675), .A2(new_n671), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n934), .B1(new_n935), .B2(new_n929), .ZN(new_n936));
  INV_X1    g0736(.A(new_n934), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n907), .A2(new_n676), .A3(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n936), .A2(new_n938), .A3(KEYINPUT106), .ZN(new_n939));
  XOR2_X1   g0739(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n935), .B2(new_n929), .ZN(new_n942));
  NOR3_X1   g0742(.A1(new_n907), .A2(new_n676), .A3(new_n940), .ZN(new_n943));
  OAI221_X1 g0743(.A(new_n939), .B1(KEYINPUT106), .B2(new_n936), .C1(new_n942), .C2(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n944), .A2(new_n673), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n672), .B(new_n674), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n668), .B(new_n946), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n713), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT107), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n944), .A2(new_n950), .A3(new_n673), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n944), .A2(new_n673), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(KEYINPUT107), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n949), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n933), .B1(new_n954), .B2(new_n714), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n931), .B(new_n932), .C1(new_n955), .C2(new_n718), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n766), .A2(G68), .ZN(new_n957));
  AOI22_X1  g0757(.A1(G58), .A2(new_n773), .B1(new_n733), .B2(G77), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n415), .B1(new_n736), .B2(G137), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n958), .B(new_n959), .C1(new_n404), .C2(new_n747), .ZN(new_n960));
  INV_X1    g0760(.A(new_n741), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n960), .B1(G150), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n753), .A2(G50), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n759), .A2(G143), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n957), .A2(new_n962), .A3(new_n963), .A4(new_n964), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n747), .A2(new_n813), .B1(new_n741), .B2(new_n562), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n743), .A2(new_n552), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT46), .ZN(new_n968));
  INV_X1    g0768(.A(G317), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n415), .B1(new_n735), .B2(new_n969), .C1(new_n488), .C2(new_n732), .ZN(new_n970));
  NOR3_X1   g0770(.A1(new_n966), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(G311), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n753), .A2(G283), .B1(G107), .B2(new_n761), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT109), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n971), .B1(new_n972), .B2(new_n758), .C1(new_n973), .C2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n973), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n976), .A2(KEYINPUT109), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n965), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT47), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n729), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n979), .B2(new_n978), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n914), .A2(new_n726), .A3(new_n915), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n781), .A2(new_n238), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n726), .B(new_n728), .C1(new_n679), .C2(new_n544), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n720), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n985), .B(KEYINPUT108), .Z(new_n986));
  NAND3_X1  g0786(.A1(new_n981), .A2(new_n982), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n956), .A2(new_n987), .ZN(G387));
  AOI21_X1  g0788(.A(new_n271), .B1(new_n736), .B2(G326), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n761), .A2(G283), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n813), .B2(new_n743), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n797), .A2(G311), .B1(new_n961), .B2(G317), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n992), .B1(new_n752), .B2(new_n562), .C1(new_n758), .C2(new_n738), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT48), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n991), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n994), .B2(new_n993), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT49), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n989), .B1(new_n552), .B2(new_n732), .C1(new_n996), .C2(new_n997), .ZN(new_n998));
  AND2_X1   g0798(.A1(new_n996), .A2(new_n997), .ZN(new_n999));
  INV_X1    g0799(.A(new_n766), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n1000), .A2(new_n374), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(G77), .A2(new_n773), .B1(new_n736), .B2(G150), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n415), .B1(new_n733), .B2(G97), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n1002), .B(new_n1003), .C1(new_n747), .C2(new_n285), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(G50), .B2(new_n961), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n1005), .B1(new_n202), .B2(new_n752), .C1(new_n404), .C2(new_n758), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n998), .A2(new_n999), .B1(new_n1001), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n728), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n672), .A2(new_n726), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n682), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n786), .A2(new_n1010), .B1(new_n364), .B2(new_n679), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n235), .A2(new_n260), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n285), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n240), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT50), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n682), .B(new_n783), .C1(new_n202), .C2(new_n275), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n781), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1011), .B1(new_n1012), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n720), .B1(new_n1018), .B2(new_n780), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1008), .A2(new_n1009), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n713), .A2(new_n947), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(KEYINPUT110), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1022), .A2(new_n680), .A3(new_n948), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1021), .A2(KEYINPUT110), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1020), .B1(new_n717), .B2(new_n947), .C1(new_n1023), .C2(new_n1024), .ZN(G393));
  INV_X1    g0825(.A(new_n945), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(new_n952), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n948), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1028), .A2(new_n954), .A3(new_n680), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1026), .A2(new_n718), .A3(new_n952), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n779), .B1(new_n488), .B2(new_n212), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(new_n250), .B2(new_n781), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1032), .A2(new_n720), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT111), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n758), .A2(new_n969), .B1(new_n972), .B2(new_n741), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT52), .Z(new_n1036));
  NAND2_X1  g0836(.A1(new_n797), .A2(G303), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n271), .B1(new_n733), .B2(G107), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(G283), .A2(new_n773), .B1(new_n736), .B2(G322), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(G116), .B2(new_n761), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n813), .B2(new_n752), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n758), .A2(new_n283), .B1(new_n404), .B2(new_n741), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT51), .Z(new_n1044));
  NAND2_X1  g0844(.A1(new_n766), .A2(G77), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n271), .B1(new_n732), .B2(new_n222), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n743), .A2(new_n202), .B1(new_n735), .B2(new_n800), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n1046), .B(new_n1047), .C1(new_n797), .C2(G50), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1045), .B(new_n1048), .C1(new_n285), .C2(new_n752), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n1036), .A2(new_n1042), .B1(new_n1044), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT112), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n728), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n726), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1034), .B1(new_n1053), .B2(new_n1054), .C1(new_n929), .C2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1029), .A2(new_n1030), .A3(new_n1056), .ZN(G390));
  AND3_X1   g0857(.A1(new_n847), .A2(KEYINPUT39), .A3(new_n851), .ZN(new_n1058));
  AOI21_X1  g0858(.A(KEYINPUT39), .B1(new_n870), .B2(new_n851), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n1058), .A2(new_n1059), .B1(new_n883), .B2(new_n888), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n663), .B(new_n824), .C1(new_n641), .C2(new_n653), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n886), .B1(new_n1061), .B2(new_n819), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1062), .A2(new_n882), .A3(new_n879), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n853), .A2(G330), .A3(new_n828), .A4(new_n886), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(KEYINPUT113), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT113), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n711), .A2(new_n1066), .A3(new_n828), .A4(new_n886), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n1060), .A2(new_n1063), .A3(new_n1065), .A4(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1064), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n881), .A2(new_n884), .B1(new_n882), .B2(new_n1062), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1063), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1069), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1068), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n459), .A2(new_n711), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n891), .A2(new_n634), .A3(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n886), .B1(new_n711), .B2(new_n828), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n1076), .A2(new_n1069), .B1(new_n819), .B2(new_n1061), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1061), .A2(new_n819), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n853), .A2(G330), .A3(new_n828), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n887), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1067), .A2(new_n1065), .A3(new_n1078), .A4(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1075), .B1(new_n1077), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1073), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1082), .A2(new_n1072), .A3(new_n1068), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1084), .A2(new_n680), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1067), .A2(new_n1065), .ZN(new_n1087));
  NOR3_X1   g0887(.A1(new_n1070), .A2(new_n1071), .A3(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1064), .B1(new_n1060), .B2(new_n1063), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n718), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n724), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n719), .B1(new_n1013), .B2(new_n795), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n741), .A2(new_n552), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n736), .A2(G294), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n774), .A2(new_n804), .A3(new_n1095), .A4(new_n415), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n1094), .B(new_n1096), .C1(G107), .C2(new_n797), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n759), .A2(G283), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n753), .A2(G97), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1045), .A2(new_n1097), .A3(new_n1098), .A4(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n773), .A2(G150), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT53), .ZN(new_n1102));
  INV_X1    g0902(.A(G125), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n271), .B1(new_n735), .B2(new_n1103), .C1(new_n240), .C2(new_n732), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n1102), .B(new_n1104), .C1(new_n766), .C2(G159), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(KEYINPUT54), .B(G143), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT114), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n753), .A2(new_n1107), .B1(G137), .B2(new_n797), .ZN(new_n1108));
  OR2_X1    g0908(.A1(new_n1108), .A2(KEYINPUT115), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(KEYINPUT115), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1105), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(G128), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n758), .A2(new_n1112), .B1(new_n805), .B2(new_n741), .ZN(new_n1113));
  XOR2_X1   g0913(.A(new_n1113), .B(KEYINPUT116), .Z(new_n1114));
  OAI21_X1  g0914(.A(new_n1100), .B1(new_n1111), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1093), .B1(new_n1115), .B2(new_n728), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1092), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1086), .A2(new_n1091), .A3(new_n1117), .ZN(G378));
  NAND2_X1  g0918(.A1(new_n837), .A2(new_n358), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n361), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1120), .B1(new_n629), .B2(new_n1121), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n361), .B(new_n1119), .C1(new_n628), .C2(new_n625), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1122), .A2(new_n1123), .A3(new_n1125), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(new_n872), .B2(G330), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n879), .A2(KEYINPUT40), .A3(new_n862), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n853), .A2(new_n861), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(new_n847), .B2(new_n851), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1131), .B(G330), .C1(KEYINPUT40), .C2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1129), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(KEYINPUT118), .B1(new_n1130), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n885), .A2(new_n889), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(KEYINPUT119), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT119), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n885), .A2(new_n1140), .A3(new_n889), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1137), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n863), .A2(new_n864), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1145), .A2(G330), .A3(new_n1131), .A4(new_n1129), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1147), .A2(KEYINPUT118), .A3(new_n1139), .A4(new_n1141), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1143), .A2(new_n718), .A3(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1135), .A2(new_n724), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n719), .B1(G50), .B2(new_n795), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(G33), .A2(G41), .ZN(new_n1152));
  AOI211_X1 g0952(.A(G50), .B(new_n1152), .C1(new_n415), .C2(new_n264), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n741), .A2(new_n364), .ZN(new_n1154));
  AOI211_X1 g0954(.A(G41), .B(new_n271), .C1(new_n736), .C2(G283), .ZN(new_n1155));
  OAI221_X1 g0955(.A(new_n1155), .B1(new_n201), .B2(new_n732), .C1(new_n275), .C2(new_n743), .ZN(new_n1156));
  AOI211_X1 g0956(.A(new_n1154), .B(new_n1156), .C1(G97), .C2(new_n797), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n753), .A2(new_n544), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n759), .A2(G116), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1157), .A2(new_n957), .A3(new_n1158), .A4(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT58), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1153), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n797), .A2(G132), .B1(new_n773), .B2(new_n1107), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(new_n1112), .B2(new_n741), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(G137), .B2(new_n753), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n1165), .B1(new_n1103), .B2(new_n758), .C1(new_n283), .C2(new_n1000), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(KEYINPUT59), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1152), .B1(new_n732), .B2(new_n404), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(G124), .B2(new_n736), .ZN(new_n1169));
  XOR2_X1   g0969(.A(new_n1169), .B(KEYINPUT117), .Z(new_n1170));
  NAND2_X1  g0970(.A1(new_n1167), .A2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1166), .A2(KEYINPUT59), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n1162), .B1(new_n1161), .B2(new_n1160), .C1(new_n1171), .C2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1151), .B1(new_n1173), .B2(new_n728), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1150), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1149), .A2(new_n1175), .ZN(new_n1176));
  AND3_X1   g0976(.A1(new_n1144), .A2(new_n890), .A3(new_n1146), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n890), .B1(new_n1146), .B2(new_n1144), .ZN(new_n1178));
  OAI21_X1  g0978(.A(KEYINPUT57), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1077), .A2(new_n1081), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1075), .B1(new_n1090), .B2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n680), .B1(new_n1179), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1075), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1085), .A2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1143), .A2(new_n1148), .A3(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT57), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT120), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1182), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1185), .A2(KEYINPUT120), .A3(new_n1186), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1176), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(G375));
  INV_X1    g0992(.A(new_n1180), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(new_n1075), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n933), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1194), .A2(new_n1083), .A3(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n719), .B1(G68), .B2(new_n795), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n961), .A2(G283), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n271), .B1(new_n733), .B2(G77), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1198), .B1(new_n552), .B2(new_n747), .C1(KEYINPUT121), .C2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(KEYINPUT121), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n1201), .B1(new_n488), .B2(new_n743), .C1(new_n562), .C2(new_n735), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1200), .A2(new_n1202), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n1203), .B1(new_n364), .B2(new_n752), .C1(new_n813), .C2(new_n758), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n743), .A2(new_n404), .B1(new_n735), .B2(new_n1112), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n415), .B(new_n1205), .C1(G58), .C2(new_n733), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1206), .B1(new_n283), .B2(new_n752), .C1(new_n1000), .C2(new_n240), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n797), .A2(new_n1107), .B1(new_n961), .B2(G137), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1208), .B1(new_n758), .B2(new_n805), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(KEYINPUT122), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n1204), .A2(new_n1001), .B1(new_n1207), .B2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1197), .B1(new_n1211), .B2(new_n728), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n886), .B2(new_n725), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1213), .B1(new_n1193), .B2(new_n717), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1196), .A2(new_n1215), .ZN(G381));
  OR2_X1    g1016(.A1(G393), .A2(G396), .ZN(new_n1217));
  NOR4_X1   g1017(.A1(G390), .A2(G384), .A3(G381), .A4(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n987), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n954), .A2(new_n714), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(new_n1195), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(new_n717), .ZN(new_n1222));
  AND2_X1   g1022(.A1(new_n931), .A2(new_n932), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1219), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(G378), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1218), .A2(new_n1224), .A3(new_n1225), .A4(new_n1191), .ZN(G407));
  NAND2_X1  g1026(.A1(new_n662), .A2(G213), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1191), .A2(new_n1225), .A3(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(G407), .A2(G213), .A3(new_n1229), .ZN(G409));
  INV_X1    g1030(.A(KEYINPUT60), .ZN(new_n1231));
  NOR3_X1   g1031(.A1(new_n1180), .A2(new_n1183), .A3(new_n1231), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1232), .A2(new_n681), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1194), .B1(new_n1231), .B2(new_n1082), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1214), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  XOR2_X1   g1035(.A(new_n1235), .B(G384), .Z(new_n1236));
  AOI211_X1 g1036(.A(new_n1225), .B(new_n1176), .C1(new_n1189), .C2(new_n1190), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1147), .A2(new_n1138), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1144), .A2(new_n890), .A3(new_n1146), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  OR2_X1    g1040(.A1(new_n1240), .A2(KEYINPUT123), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n717), .B1(new_n1240), .B2(KEYINPUT123), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n1241), .A2(new_n1242), .B1(new_n1150), .B2(new_n1174), .ZN(new_n1243));
  OR2_X1    g1043(.A1(new_n1185), .A2(new_n933), .ZN(new_n1244));
  AOI21_X1  g1044(.A(G378), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1227), .B(new_n1236), .C1(new_n1237), .C2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(KEYINPUT62), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT61), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1228), .A2(G2897), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1236), .B(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1245), .B1(new_n1191), .B2(G378), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1251), .B1(new_n1252), .B2(new_n1228), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1240), .A2(KEYINPUT57), .A3(new_n1184), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1254), .A2(new_n680), .A3(new_n1190), .A4(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1176), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1256), .A2(G378), .A3(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1245), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT62), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1260), .A2(new_n1261), .A3(new_n1227), .A4(new_n1236), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1247), .A2(new_n1248), .A3(new_n1253), .A4(new_n1262), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(G393), .B(G396), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT124), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(new_n1224), .B2(G390), .ZN(new_n1266));
  INV_X1    g1066(.A(G390), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(G387), .A2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1264), .B1(new_n1266), .B2(new_n1268), .ZN(new_n1269));
  NOR3_X1   g1069(.A1(new_n1224), .A2(KEYINPUT124), .A3(G390), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n956), .A2(KEYINPUT125), .A3(G390), .A4(new_n987), .ZN(new_n1272));
  AND3_X1   g1072(.A1(new_n1268), .A2(new_n1272), .A3(new_n1264), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n956), .A2(new_n987), .A3(G390), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT125), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  AOI22_X1  g1076(.A1(new_n1269), .A2(new_n1271), .B1(new_n1273), .B2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1263), .A2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1260), .A2(new_n1227), .ZN(new_n1279));
  AOI21_X1  g1079(.A(KEYINPUT61), .B1(new_n1279), .B2(new_n1251), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1276), .A2(new_n1268), .A3(new_n1272), .A4(new_n1264), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1264), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1274), .A2(KEYINPUT124), .ZN(new_n1283));
  AOI21_X1  g1083(.A(G390), .B1(new_n956), .B2(new_n987), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1282), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1281), .B1(new_n1285), .B2(new_n1270), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT63), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1246), .A2(new_n1287), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1260), .A2(KEYINPUT63), .A3(new_n1227), .A4(new_n1236), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1280), .A2(new_n1286), .A3(new_n1288), .A4(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1278), .A2(new_n1290), .ZN(G405));
  NOR2_X1   g1091(.A1(new_n1191), .A2(G378), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1292), .A2(new_n1237), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT126), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1293), .A2(new_n1294), .A3(new_n1236), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1236), .A2(new_n1294), .ZN(new_n1296));
  OR2_X1    g1096(.A1(new_n1236), .A2(new_n1294), .ZN(new_n1297));
  OAI211_X1 g1097(.A(new_n1296), .B(new_n1297), .C1(new_n1292), .C2(new_n1237), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1277), .A2(new_n1295), .A3(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1295), .A2(new_n1298), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n1286), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1299), .A2(new_n1301), .ZN(G402));
endmodule


