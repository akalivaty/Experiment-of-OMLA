

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587;

  XNOR2_X1 U320 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U321 ( .A(n383), .B(KEYINPUT46), .ZN(n384) );
  XOR2_X1 U322 ( .A(KEYINPUT28), .B(n475), .Z(n536) );
  AND2_X1 U323 ( .A1(G232GAT), .A2(G233GAT), .ZN(n288) );
  XOR2_X1 U324 ( .A(G162GAT), .B(KEYINPUT73), .Z(n289) );
  INV_X1 U325 ( .A(KEYINPUT111), .ZN(n383) );
  XNOR2_X1 U326 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n390) );
  XNOR2_X1 U327 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U328 ( .A(n404), .B(n288), .ZN(n311) );
  XNOR2_X1 U329 ( .A(n429), .B(n311), .ZN(n314) );
  XNOR2_X1 U330 ( .A(n365), .B(n364), .ZN(n371) );
  XNOR2_X1 U331 ( .A(n371), .B(n424), .ZN(n372) );
  XNOR2_X1 U332 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U333 ( .A(n323), .B(n322), .ZN(n328) );
  XNOR2_X1 U334 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U335 ( .A(n382), .B(n381), .ZN(n577) );
  XOR2_X1 U336 ( .A(n452), .B(n451), .Z(n538) );
  XNOR2_X1 U337 ( .A(n458), .B(G190GAT), .ZN(n459) );
  XNOR2_X1 U338 ( .A(n460), .B(n459), .ZN(G1351GAT) );
  XOR2_X1 U339 ( .A(KEYINPUT5), .B(KEYINPUT89), .Z(n291) );
  XNOR2_X1 U340 ( .A(G162GAT), .B(G85GAT), .ZN(n290) );
  XNOR2_X1 U341 ( .A(n291), .B(n290), .ZN(n292) );
  XOR2_X1 U342 ( .A(n292), .B(KEYINPUT6), .Z(n295) );
  INV_X1 U343 ( .A(G148GAT), .ZN(n293) );
  XOR2_X1 U344 ( .A(G120GAT), .B(G57GAT), .Z(n365) );
  XNOR2_X1 U345 ( .A(G148GAT), .B(n365), .ZN(n294) );
  XNOR2_X1 U346 ( .A(n295), .B(n294), .ZN(n298) );
  XOR2_X1 U347 ( .A(G155GAT), .B(KEYINPUT2), .Z(n297) );
  XNOR2_X1 U348 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n296) );
  XNOR2_X1 U349 ( .A(n297), .B(n296), .ZN(n420) );
  XOR2_X1 U350 ( .A(n298), .B(n420), .Z(n300) );
  XOR2_X1 U351 ( .A(G113GAT), .B(G1GAT), .Z(n360) );
  XOR2_X1 U352 ( .A(KEYINPUT0), .B(G127GAT), .Z(n441) );
  XNOR2_X1 U353 ( .A(n360), .B(n441), .ZN(n299) );
  XNOR2_X1 U354 ( .A(n300), .B(n299), .ZN(n309) );
  XOR2_X1 U355 ( .A(KEYINPUT4), .B(KEYINPUT91), .Z(n302) );
  XNOR2_X1 U356 ( .A(KEYINPUT92), .B(KEYINPUT1), .ZN(n301) );
  XNOR2_X1 U357 ( .A(n302), .B(n301), .ZN(n307) );
  XNOR2_X1 U358 ( .A(G29GAT), .B(G134GAT), .ZN(n303) );
  XNOR2_X1 U359 ( .A(n303), .B(KEYINPUT75), .ZN(n326) );
  XOR2_X1 U360 ( .A(KEYINPUT90), .B(n326), .Z(n305) );
  NAND2_X1 U361 ( .A1(G225GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U362 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U363 ( .A(n307), .B(n306), .Z(n308) );
  XNOR2_X1 U364 ( .A(n309), .B(n308), .ZN(n472) );
  XNOR2_X1 U365 ( .A(KEYINPUT93), .B(n472), .ZN(n522) );
  INV_X1 U366 ( .A(KEYINPUT54), .ZN(n416) );
  XNOR2_X1 U367 ( .A(G50GAT), .B(G218GAT), .ZN(n310) );
  XNOR2_X1 U368 ( .A(n289), .B(n310), .ZN(n429) );
  XOR2_X1 U369 ( .A(G36GAT), .B(G190GAT), .Z(n404) );
  INV_X1 U370 ( .A(n314), .ZN(n313) );
  INV_X1 U371 ( .A(KEYINPUT76), .ZN(n312) );
  NAND2_X1 U372 ( .A1(n313), .A2(n312), .ZN(n316) );
  NAND2_X1 U373 ( .A1(n314), .A2(KEYINPUT76), .ZN(n315) );
  NAND2_X1 U374 ( .A1(n316), .A2(n315), .ZN(n323) );
  XNOR2_X1 U375 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n317) );
  XNOR2_X1 U376 ( .A(n317), .B(KEYINPUT7), .ZN(n361) );
  XOR2_X1 U377 ( .A(n361), .B(KEYINPUT11), .Z(n321) );
  XOR2_X1 U378 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n319) );
  XNOR2_X1 U379 ( .A(KEYINPUT64), .B(KEYINPUT74), .ZN(n318) );
  XOR2_X1 U380 ( .A(n319), .B(n318), .Z(n320) );
  XOR2_X1 U381 ( .A(G92GAT), .B(G85GAT), .Z(n325) );
  XNOR2_X1 U382 ( .A(G99GAT), .B(G106GAT), .ZN(n324) );
  XNOR2_X1 U383 ( .A(n325), .B(n324), .ZN(n373) );
  XNOR2_X1 U384 ( .A(n326), .B(n373), .ZN(n327) );
  XNOR2_X1 U385 ( .A(n328), .B(n327), .ZN(n563) );
  XOR2_X1 U386 ( .A(G155GAT), .B(G78GAT), .Z(n330) );
  XNOR2_X1 U387 ( .A(G127GAT), .B(G211GAT), .ZN(n329) );
  XNOR2_X1 U388 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U389 ( .A(n331), .B(G57GAT), .Z(n333) );
  XOR2_X1 U390 ( .A(G15GAT), .B(G22GAT), .Z(n358) );
  XNOR2_X1 U391 ( .A(G1GAT), .B(n358), .ZN(n332) );
  XNOR2_X1 U392 ( .A(n333), .B(n332), .ZN(n338) );
  XNOR2_X1 U393 ( .A(G8GAT), .B(G183GAT), .ZN(n334) );
  XNOR2_X1 U394 ( .A(n334), .B(KEYINPUT78), .ZN(n402) );
  XOR2_X1 U395 ( .A(G71GAT), .B(KEYINPUT13), .Z(n378) );
  XOR2_X1 U396 ( .A(n402), .B(n378), .Z(n336) );
  NAND2_X1 U397 ( .A1(G231GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U398 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U399 ( .A(n338), .B(n337), .Z(n346) );
  XOR2_X1 U400 ( .A(KEYINPUT14), .B(KEYINPUT82), .Z(n340) );
  XNOR2_X1 U401 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n339) );
  XNOR2_X1 U402 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U403 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n342) );
  XNOR2_X1 U404 ( .A(KEYINPUT79), .B(KEYINPUT15), .ZN(n341) );
  XNOR2_X1 U405 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U406 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U407 ( .A(n346), .B(n345), .ZN(n582) );
  NAND2_X1 U408 ( .A1(n563), .A2(n582), .ZN(n387) );
  XOR2_X1 U409 ( .A(KEYINPUT66), .B(KEYINPUT67), .Z(n348) );
  NAND2_X1 U410 ( .A1(G229GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U411 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U412 ( .A(n349), .B(KEYINPUT29), .Z(n357) );
  XOR2_X1 U413 ( .A(G36GAT), .B(G50GAT), .Z(n351) );
  XNOR2_X1 U414 ( .A(G169GAT), .B(G29GAT), .ZN(n350) );
  XNOR2_X1 U415 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U416 ( .A(KEYINPUT30), .B(G8GAT), .Z(n353) );
  XNOR2_X1 U417 ( .A(G197GAT), .B(G141GAT), .ZN(n352) );
  XNOR2_X1 U418 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U419 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U420 ( .A(n357), .B(n356), .ZN(n359) );
  XOR2_X1 U421 ( .A(n359), .B(n358), .Z(n363) );
  XNOR2_X1 U422 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U423 ( .A(n363), .B(n362), .ZN(n571) );
  AND2_X1 U424 ( .A1(G230GAT), .A2(G233GAT), .ZN(n364) );
  NAND2_X1 U425 ( .A1(n293), .A2(G78GAT), .ZN(n368) );
  INV_X1 U426 ( .A(G78GAT), .ZN(n366) );
  NAND2_X1 U427 ( .A1(n366), .A2(G148GAT), .ZN(n367) );
  NAND2_X1 U428 ( .A1(n368), .A2(n367), .ZN(n370) );
  XNOR2_X1 U429 ( .A(G204GAT), .B(KEYINPUT68), .ZN(n369) );
  XNOR2_X1 U430 ( .A(n370), .B(n369), .ZN(n424) );
  XOR2_X1 U431 ( .A(KEYINPUT71), .B(n372), .Z(n375) );
  XNOR2_X1 U432 ( .A(n373), .B(KEYINPUT70), .ZN(n374) );
  XNOR2_X1 U433 ( .A(n375), .B(n374), .ZN(n382) );
  XOR2_X1 U434 ( .A(KEYINPUT31), .B(KEYINPUT69), .Z(n377) );
  XNOR2_X1 U435 ( .A(KEYINPUT32), .B(KEYINPUT33), .ZN(n376) );
  XOR2_X1 U436 ( .A(n377), .B(n376), .Z(n380) );
  XOR2_X1 U437 ( .A(G176GAT), .B(G64GAT), .Z(n405) );
  XNOR2_X1 U438 ( .A(n378), .B(n405), .ZN(n379) );
  XOR2_X1 U439 ( .A(n577), .B(KEYINPUT41), .Z(n556) );
  NOR2_X1 U440 ( .A1(n571), .A2(n556), .ZN(n385) );
  NOR2_X1 U441 ( .A1(n387), .A2(n386), .ZN(n388) );
  XNOR2_X1 U442 ( .A(n388), .B(KEYINPUT47), .ZN(n395) );
  INV_X1 U443 ( .A(n577), .ZN(n461) );
  INV_X1 U444 ( .A(KEYINPUT77), .ZN(n389) );
  XNOR2_X1 U445 ( .A(n389), .B(n563), .ZN(n548) );
  XNOR2_X1 U446 ( .A(KEYINPUT36), .B(n548), .ZN(n490) );
  NOR2_X1 U447 ( .A1(n582), .A2(n490), .ZN(n391) );
  NOR2_X1 U448 ( .A1(n461), .A2(n392), .ZN(n393) );
  NAND2_X1 U449 ( .A1(n393), .A2(n571), .ZN(n394) );
  NAND2_X1 U450 ( .A1(n395), .A2(n394), .ZN(n396) );
  XOR2_X1 U451 ( .A(KEYINPUT48), .B(n396), .Z(n534) );
  XOR2_X1 U452 ( .A(KEYINPUT95), .B(G92GAT), .Z(n398) );
  XNOR2_X1 U453 ( .A(G204GAT), .B(G218GAT), .ZN(n397) );
  XNOR2_X1 U454 ( .A(n398), .B(n397), .ZN(n409) );
  XNOR2_X1 U455 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n399) );
  XNOR2_X1 U456 ( .A(n399), .B(G211GAT), .ZN(n425) );
  XOR2_X1 U457 ( .A(KEYINPUT94), .B(n425), .Z(n401) );
  NAND2_X1 U458 ( .A1(G226GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U459 ( .A(n401), .B(n400), .ZN(n403) );
  XOR2_X1 U460 ( .A(n403), .B(n402), .Z(n407) );
  XNOR2_X1 U461 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U462 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U463 ( .A(n409), .B(n408), .ZN(n414) );
  XOR2_X1 U464 ( .A(KEYINPUT84), .B(KEYINPUT17), .Z(n411) );
  XNOR2_X1 U465 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n410) );
  XNOR2_X1 U466 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U467 ( .A(G169GAT), .B(n412), .Z(n448) );
  INV_X1 U468 ( .A(n448), .ZN(n413) );
  XOR2_X1 U469 ( .A(n414), .B(n413), .Z(n524) );
  INV_X1 U470 ( .A(n524), .ZN(n468) );
  NOR2_X1 U471 ( .A1(n534), .A2(n468), .ZN(n415) );
  XNOR2_X1 U472 ( .A(n416), .B(n415), .ZN(n417) );
  NOR2_X1 U473 ( .A1(n522), .A2(n417), .ZN(n570) );
  XOR2_X1 U474 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n419) );
  XNOR2_X1 U475 ( .A(G22GAT), .B(KEYINPUT23), .ZN(n418) );
  XNOR2_X1 U476 ( .A(n419), .B(n418), .ZN(n433) );
  XOR2_X1 U477 ( .A(KEYINPUT86), .B(n420), .Z(n422) );
  NAND2_X1 U478 ( .A1(G228GAT), .A2(G233GAT), .ZN(n421) );
  XNOR2_X1 U479 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U480 ( .A(n423), .B(G106GAT), .Z(n427) );
  XNOR2_X1 U481 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U482 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U483 ( .A(n428), .B(KEYINPUT88), .Z(n431) );
  XNOR2_X1 U484 ( .A(n429), .B(KEYINPUT87), .ZN(n430) );
  XNOR2_X1 U485 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U486 ( .A(n433), .B(n432), .ZN(n475) );
  NAND2_X1 U487 ( .A1(n570), .A2(n475), .ZN(n435) );
  XOR2_X1 U488 ( .A(KEYINPUT55), .B(KEYINPUT119), .Z(n434) );
  XNOR2_X1 U489 ( .A(n435), .B(n434), .ZN(n453) );
  XOR2_X1 U490 ( .A(G120GAT), .B(G183GAT), .Z(n437) );
  XNOR2_X1 U491 ( .A(G113GAT), .B(G15GAT), .ZN(n436) );
  XNOR2_X1 U492 ( .A(n437), .B(n436), .ZN(n452) );
  XOR2_X1 U493 ( .A(G176GAT), .B(G71GAT), .Z(n439) );
  XNOR2_X1 U494 ( .A(G134GAT), .B(G190GAT), .ZN(n438) );
  XNOR2_X1 U495 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U496 ( .A(n440), .B(G99GAT), .Z(n443) );
  XNOR2_X1 U497 ( .A(G43GAT), .B(n441), .ZN(n442) );
  XNOR2_X1 U498 ( .A(n443), .B(n442), .ZN(n447) );
  XOR2_X1 U499 ( .A(KEYINPUT20), .B(KEYINPUT85), .Z(n445) );
  NAND2_X1 U500 ( .A1(G227GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U501 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U502 ( .A(n447), .B(n446), .Z(n450) );
  XNOR2_X1 U503 ( .A(n448), .B(KEYINPUT83), .ZN(n449) );
  XNOR2_X1 U504 ( .A(n450), .B(n449), .ZN(n451) );
  NAND2_X1 U505 ( .A1(n453), .A2(n538), .ZN(n566) );
  XNOR2_X1 U506 ( .A(n556), .B(KEYINPUT104), .ZN(n540) );
  NOR2_X1 U507 ( .A1(n566), .A2(n540), .ZN(n457) );
  XNOR2_X1 U508 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n455) );
  XNOR2_X1 U509 ( .A(G176GAT), .B(KEYINPUT120), .ZN(n454) );
  XNOR2_X1 U510 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U511 ( .A(n457), .B(n456), .ZN(G1349GAT) );
  NOR2_X1 U512 ( .A1(n548), .A2(n566), .ZN(n460) );
  XNOR2_X1 U513 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n458) );
  NOR2_X1 U514 ( .A1(n461), .A2(n571), .ZN(n462) );
  XOR2_X1 U515 ( .A(n462), .B(KEYINPUT72), .Z(n495) );
  INV_X1 U516 ( .A(n582), .ZN(n463) );
  NAND2_X1 U517 ( .A1(n548), .A2(n463), .ZN(n464) );
  XOR2_X1 U518 ( .A(KEYINPUT16), .B(n464), .Z(n480) );
  NAND2_X1 U519 ( .A1(n538), .A2(n524), .ZN(n465) );
  NAND2_X1 U520 ( .A1(n475), .A2(n465), .ZN(n466) );
  XOR2_X1 U521 ( .A(KEYINPUT25), .B(n466), .Z(n471) );
  XOR2_X1 U522 ( .A(KEYINPUT27), .B(KEYINPUT96), .Z(n467) );
  XNOR2_X1 U523 ( .A(n468), .B(n467), .ZN(n474) );
  NOR2_X1 U524 ( .A1(n475), .A2(n538), .ZN(n469) );
  XNOR2_X1 U525 ( .A(n469), .B(KEYINPUT26), .ZN(n569) );
  NAND2_X1 U526 ( .A1(n474), .A2(n569), .ZN(n470) );
  NAND2_X1 U527 ( .A1(n471), .A2(n470), .ZN(n473) );
  NAND2_X1 U528 ( .A1(n473), .A2(n472), .ZN(n479) );
  NAND2_X1 U529 ( .A1(n522), .A2(n474), .ZN(n533) );
  NOR2_X1 U530 ( .A1(n533), .A2(n536), .ZN(n477) );
  INV_X1 U531 ( .A(n538), .ZN(n476) );
  NAND2_X1 U532 ( .A1(n477), .A2(n476), .ZN(n478) );
  NAND2_X1 U533 ( .A1(n479), .A2(n478), .ZN(n491) );
  NAND2_X1 U534 ( .A1(n480), .A2(n491), .ZN(n509) );
  NOR2_X1 U535 ( .A1(n495), .A2(n509), .ZN(n487) );
  NAND2_X1 U536 ( .A1(n487), .A2(n522), .ZN(n481) );
  XNOR2_X1 U537 ( .A(n481), .B(KEYINPUT34), .ZN(n482) );
  XNOR2_X1 U538 ( .A(G1GAT), .B(n482), .ZN(G1324GAT) );
  NAND2_X1 U539 ( .A1(n487), .A2(n524), .ZN(n483) );
  XNOR2_X1 U540 ( .A(n483), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U541 ( .A(KEYINPUT97), .B(KEYINPUT35), .Z(n485) );
  NAND2_X1 U542 ( .A1(n487), .A2(n538), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n485), .B(n484), .ZN(n486) );
  XOR2_X1 U544 ( .A(G15GAT), .B(n486), .Z(G1326GAT) );
  NAND2_X1 U545 ( .A1(n536), .A2(n487), .ZN(n488) );
  XNOR2_X1 U546 ( .A(n488), .B(KEYINPUT98), .ZN(n489) );
  XNOR2_X1 U547 ( .A(G22GAT), .B(n489), .ZN(G1327GAT) );
  NAND2_X1 U548 ( .A1(n582), .A2(n491), .ZN(n492) );
  NOR2_X1 U549 ( .A1(n490), .A2(n492), .ZN(n494) );
  XNOR2_X1 U550 ( .A(KEYINPUT37), .B(KEYINPUT99), .ZN(n493) );
  XOR2_X1 U551 ( .A(n494), .B(n493), .Z(n521) );
  OR2_X1 U552 ( .A1(n521), .A2(n495), .ZN(n496) );
  XOR2_X1 U553 ( .A(KEYINPUT38), .B(n496), .Z(n505) );
  NAND2_X1 U554 ( .A1(n522), .A2(n505), .ZN(n498) );
  XOR2_X1 U555 ( .A(G29GAT), .B(KEYINPUT39), .Z(n497) );
  XNOR2_X1 U556 ( .A(n498), .B(n497), .ZN(G1328GAT) );
  NAND2_X1 U557 ( .A1(n505), .A2(n524), .ZN(n499) );
  XNOR2_X1 U558 ( .A(n499), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U559 ( .A(KEYINPUT40), .B(KEYINPUT102), .Z(n501) );
  XNOR2_X1 U560 ( .A(G43GAT), .B(KEYINPUT101), .ZN(n500) );
  XNOR2_X1 U561 ( .A(n501), .B(n500), .ZN(n504) );
  NAND2_X1 U562 ( .A1(n505), .A2(n538), .ZN(n502) );
  XNOR2_X1 U563 ( .A(n502), .B(KEYINPUT100), .ZN(n503) );
  XNOR2_X1 U564 ( .A(n504), .B(n503), .ZN(G1330GAT) );
  XOR2_X1 U565 ( .A(G50GAT), .B(KEYINPUT103), .Z(n507) );
  NAND2_X1 U566 ( .A1(n505), .A2(n536), .ZN(n506) );
  XNOR2_X1 U567 ( .A(n507), .B(n506), .ZN(G1331GAT) );
  INV_X1 U568 ( .A(n540), .ZN(n508) );
  NAND2_X1 U569 ( .A1(n571), .A2(n508), .ZN(n520) );
  NOR2_X1 U570 ( .A1(n520), .A2(n509), .ZN(n517) );
  NAND2_X1 U571 ( .A1(n522), .A2(n517), .ZN(n510) );
  XNOR2_X1 U572 ( .A(KEYINPUT42), .B(n510), .ZN(n511) );
  XNOR2_X1 U573 ( .A(G57GAT), .B(n511), .ZN(G1332GAT) );
  XOR2_X1 U574 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n513) );
  NAND2_X1 U575 ( .A1(n517), .A2(n524), .ZN(n512) );
  XNOR2_X1 U576 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U577 ( .A(G64GAT), .B(n514), .ZN(G1333GAT) );
  XOR2_X1 U578 ( .A(G71GAT), .B(KEYINPUT107), .Z(n516) );
  NAND2_X1 U579 ( .A1(n517), .A2(n538), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n516), .B(n515), .ZN(G1334GAT) );
  XOR2_X1 U581 ( .A(G78GAT), .B(KEYINPUT43), .Z(n519) );
  NAND2_X1 U582 ( .A1(n517), .A2(n536), .ZN(n518) );
  XNOR2_X1 U583 ( .A(n519), .B(n518), .ZN(G1335GAT) );
  NOR2_X1 U584 ( .A1(n521), .A2(n520), .ZN(n530) );
  NAND2_X1 U585 ( .A1(n530), .A2(n522), .ZN(n523) );
  XNOR2_X1 U586 ( .A(n523), .B(G85GAT), .ZN(G1336GAT) );
  XOR2_X1 U587 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n526) );
  NAND2_X1 U588 ( .A1(n530), .A2(n524), .ZN(n525) );
  XNOR2_X1 U589 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U590 ( .A(G92GAT), .B(n527), .ZN(G1337GAT) );
  NAND2_X1 U591 ( .A1(n530), .A2(n538), .ZN(n528) );
  XNOR2_X1 U592 ( .A(n528), .B(KEYINPUT110), .ZN(n529) );
  XNOR2_X1 U593 ( .A(G99GAT), .B(n529), .ZN(G1338GAT) );
  NAND2_X1 U594 ( .A1(n536), .A2(n530), .ZN(n531) );
  XNOR2_X1 U595 ( .A(n531), .B(KEYINPUT44), .ZN(n532) );
  XNOR2_X1 U596 ( .A(G106GAT), .B(n532), .ZN(G1339GAT) );
  NOR2_X1 U597 ( .A1(n534), .A2(n533), .ZN(n535) );
  XOR2_X1 U598 ( .A(KEYINPUT112), .B(n535), .Z(n552) );
  NOR2_X1 U599 ( .A1(n552), .A2(n536), .ZN(n537) );
  NAND2_X1 U600 ( .A1(n538), .A2(n537), .ZN(n547) );
  NOR2_X1 U601 ( .A1(n571), .A2(n547), .ZN(n539) );
  XOR2_X1 U602 ( .A(G113GAT), .B(n539), .Z(G1340GAT) );
  NOR2_X1 U603 ( .A1(n540), .A2(n547), .ZN(n542) );
  XNOR2_X1 U604 ( .A(KEYINPUT49), .B(KEYINPUT113), .ZN(n541) );
  XNOR2_X1 U605 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U606 ( .A(G120GAT), .B(n543), .Z(G1341GAT) );
  NOR2_X1 U607 ( .A1(n582), .A2(n547), .ZN(n545) );
  XNOR2_X1 U608 ( .A(KEYINPUT114), .B(KEYINPUT50), .ZN(n544) );
  XNOR2_X1 U609 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U610 ( .A(G127GAT), .B(n546), .Z(G1342GAT) );
  NOR2_X1 U611 ( .A1(n548), .A2(n547), .ZN(n550) );
  XNOR2_X1 U612 ( .A(KEYINPUT115), .B(KEYINPUT51), .ZN(n549) );
  XNOR2_X1 U613 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U614 ( .A(G134GAT), .B(n551), .Z(G1343GAT) );
  INV_X1 U615 ( .A(n552), .ZN(n553) );
  NAND2_X1 U616 ( .A1(n569), .A2(n553), .ZN(n562) );
  NOR2_X1 U617 ( .A1(n571), .A2(n562), .ZN(n554) );
  XOR2_X1 U618 ( .A(n554), .B(KEYINPUT116), .Z(n555) );
  XNOR2_X1 U619 ( .A(G141GAT), .B(n555), .ZN(G1344GAT) );
  NOR2_X1 U620 ( .A1(n556), .A2(n562), .ZN(n558) );
  XNOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n557) );
  XNOR2_X1 U622 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(n559), .ZN(G1345GAT) );
  NOR2_X1 U624 ( .A1(n582), .A2(n562), .ZN(n561) );
  XNOR2_X1 U625 ( .A(G155GAT), .B(KEYINPUT117), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n561), .B(n560), .ZN(G1346GAT) );
  NOR2_X1 U627 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U628 ( .A(KEYINPUT118), .B(n564), .Z(n565) );
  XNOR2_X1 U629 ( .A(G162GAT), .B(n565), .ZN(G1347GAT) );
  NOR2_X1 U630 ( .A1(n571), .A2(n566), .ZN(n567) );
  XOR2_X1 U631 ( .A(G169GAT), .B(n567), .Z(G1348GAT) );
  NOR2_X1 U632 ( .A1(n582), .A2(n566), .ZN(n568) );
  XOR2_X1 U633 ( .A(G183GAT), .B(n568), .Z(G1350GAT) );
  NAND2_X1 U634 ( .A1(n570), .A2(n569), .ZN(n584) );
  NOR2_X1 U635 ( .A1(n571), .A2(n584), .ZN(n576) );
  XOR2_X1 U636 ( .A(KEYINPUT123), .B(KEYINPUT60), .Z(n573) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(KEYINPUT122), .B(n574), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n576), .B(n575), .ZN(G1352GAT) );
  NOR2_X1 U641 ( .A1(n584), .A2(n577), .ZN(n581) );
  XOR2_X1 U642 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n579) );
  XNOR2_X1 U643 ( .A(G204GAT), .B(KEYINPUT125), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(G1353GAT) );
  NOR2_X1 U646 ( .A1(n582), .A2(n584), .ZN(n583) );
  XOR2_X1 U647 ( .A(G211GAT), .B(n583), .Z(G1354GAT) );
  NOR2_X1 U648 ( .A1(n490), .A2(n584), .ZN(n586) );
  XNOR2_X1 U649 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(n587) );
  XOR2_X1 U651 ( .A(G218GAT), .B(n587), .Z(G1355GAT) );
endmodule

