

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U550 ( .A1(n717), .A2(n716), .ZN(n769) );
  BUF_X2 U551 ( .A(n866), .Z(n516) );
  XOR2_X1 U552 ( .A(KEYINPUT17), .B(n518), .Z(n866) );
  NOR2_X1 U553 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U554 ( .A1(n564), .A2(n563), .ZN(n716) );
  AND2_X1 U555 ( .A1(n744), .A2(G1996), .ZN(n718) );
  NAND2_X1 U556 ( .A1(n769), .A2(G1341), .ZN(n517) );
  NOR2_X1 U557 ( .A1(n641), .A2(G651), .ZN(n657) );
  NOR2_X1 U558 ( .A1(n527), .A2(n526), .ZN(G160) );
  NOR2_X1 U559 ( .A1(G2105), .A2(G2104), .ZN(n518) );
  NAND2_X1 U560 ( .A1(n516), .A2(G137), .ZN(n521) );
  INV_X1 U561 ( .A(G2105), .ZN(n522) );
  AND2_X2 U562 ( .A1(n522), .A2(G2104), .ZN(n865) );
  NAND2_X1 U563 ( .A1(G101), .A2(n865), .ZN(n519) );
  XOR2_X1 U564 ( .A(KEYINPUT23), .B(n519), .Z(n520) );
  NAND2_X1 U565 ( .A1(n521), .A2(n520), .ZN(n527) );
  NOR2_X1 U566 ( .A1(G2104), .A2(n522), .ZN(n869) );
  NAND2_X1 U567 ( .A1(n869), .A2(G125), .ZN(n525) );
  NAND2_X1 U568 ( .A1(G2104), .A2(G2105), .ZN(n523) );
  XOR2_X2 U569 ( .A(KEYINPUT64), .B(n523), .Z(n870) );
  NAND2_X1 U570 ( .A1(G113), .A2(n870), .ZN(n524) );
  NAND2_X1 U571 ( .A1(n525), .A2(n524), .ZN(n526) );
  NOR2_X1 U572 ( .A1(G543), .A2(G651), .ZN(n653) );
  NAND2_X1 U573 ( .A1(n653), .A2(G89), .ZN(n528) );
  XNOR2_X1 U574 ( .A(n528), .B(KEYINPUT4), .ZN(n531) );
  XNOR2_X1 U575 ( .A(G543), .B(KEYINPUT0), .ZN(n529) );
  XNOR2_X1 U576 ( .A(n529), .B(KEYINPUT65), .ZN(n641) );
  INV_X1 U577 ( .A(G651), .ZN(n533) );
  NOR2_X1 U578 ( .A1(n641), .A2(n533), .ZN(n647) );
  NAND2_X1 U579 ( .A1(G76), .A2(n647), .ZN(n530) );
  NAND2_X1 U580 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U581 ( .A(KEYINPUT5), .B(n532), .ZN(n540) );
  NAND2_X1 U582 ( .A1(G51), .A2(n657), .ZN(n536) );
  NOR2_X1 U583 ( .A1(G543), .A2(n533), .ZN(n534) );
  XOR2_X1 U584 ( .A(KEYINPUT1), .B(n534), .Z(n649) );
  NAND2_X1 U585 ( .A1(n649), .A2(G63), .ZN(n535) );
  NAND2_X1 U586 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U587 ( .A(n537), .B(KEYINPUT6), .ZN(n538) );
  XOR2_X1 U588 ( .A(KEYINPUT70), .B(n538), .Z(n539) );
  NAND2_X1 U589 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U590 ( .A(KEYINPUT7), .B(n541), .ZN(G168) );
  XOR2_X1 U591 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U592 ( .A1(G85), .A2(n653), .ZN(n543) );
  NAND2_X1 U593 ( .A1(G72), .A2(n647), .ZN(n542) );
  NAND2_X1 U594 ( .A1(n543), .A2(n542), .ZN(n547) );
  NAND2_X1 U595 ( .A1(G60), .A2(n649), .ZN(n545) );
  NAND2_X1 U596 ( .A1(G47), .A2(n657), .ZN(n544) );
  NAND2_X1 U597 ( .A1(n545), .A2(n544), .ZN(n546) );
  OR2_X1 U598 ( .A1(n547), .A2(n546), .ZN(G290) );
  XOR2_X1 U599 ( .A(G2427), .B(G2435), .Z(n549) );
  XNOR2_X1 U600 ( .A(G2454), .B(G2443), .ZN(n548) );
  XNOR2_X1 U601 ( .A(n549), .B(n548), .ZN(n556) );
  XOR2_X1 U602 ( .A(G2451), .B(KEYINPUT105), .Z(n551) );
  XNOR2_X1 U603 ( .A(G2430), .B(G2438), .ZN(n550) );
  XNOR2_X1 U604 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U605 ( .A(n552), .B(G2446), .Z(n554) );
  XNOR2_X1 U606 ( .A(G1341), .B(G1348), .ZN(n553) );
  XNOR2_X1 U607 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U608 ( .A(n556), .B(n555), .ZN(n557) );
  AND2_X1 U609 ( .A1(n557), .A2(G14), .ZN(G401) );
  AND2_X1 U610 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U611 ( .A(G57), .ZN(G237) );
  INV_X1 U612 ( .A(G69), .ZN(G235) );
  INV_X1 U613 ( .A(G108), .ZN(G238) );
  INV_X1 U614 ( .A(G120), .ZN(G236) );
  INV_X1 U615 ( .A(G132), .ZN(G219) );
  INV_X1 U616 ( .A(G82), .ZN(G220) );
  NAND2_X1 U617 ( .A1(n865), .A2(G102), .ZN(n560) );
  NAND2_X1 U618 ( .A1(G138), .A2(n516), .ZN(n558) );
  XOR2_X1 U619 ( .A(n558), .B(KEYINPUT87), .Z(n559) );
  AND2_X1 U620 ( .A1(n560), .A2(n559), .ZN(n564) );
  NAND2_X1 U621 ( .A1(n869), .A2(G126), .ZN(n562) );
  NAND2_X1 U622 ( .A1(G114), .A2(n870), .ZN(n561) );
  AND2_X1 U623 ( .A1(n562), .A2(n561), .ZN(n563) );
  INV_X1 U624 ( .A(n716), .ZN(G164) );
  NAND2_X1 U625 ( .A1(G88), .A2(n653), .ZN(n566) );
  NAND2_X1 U626 ( .A1(G75), .A2(n647), .ZN(n565) );
  NAND2_X1 U627 ( .A1(n566), .A2(n565), .ZN(n572) );
  NAND2_X1 U628 ( .A1(n657), .A2(G50), .ZN(n567) );
  XNOR2_X1 U629 ( .A(n567), .B(KEYINPUT78), .ZN(n569) );
  NAND2_X1 U630 ( .A1(G62), .A2(n649), .ZN(n568) );
  NAND2_X1 U631 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U632 ( .A(KEYINPUT79), .B(n570), .Z(n571) );
  NOR2_X1 U633 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U634 ( .A(KEYINPUT80), .B(n573), .Z(G303) );
  NAND2_X1 U635 ( .A1(G7), .A2(G661), .ZN(n574) );
  XNOR2_X1 U636 ( .A(n574), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U637 ( .A(G223), .ZN(n832) );
  AND2_X1 U638 ( .A1(G567), .A2(n832), .ZN(n575) );
  XNOR2_X1 U639 ( .A(n575), .B(KEYINPUT11), .ZN(G234) );
  XNOR2_X1 U640 ( .A(KEYINPUT67), .B(KEYINPUT13), .ZN(n580) );
  NAND2_X1 U641 ( .A1(n653), .A2(G81), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n576), .B(KEYINPUT12), .ZN(n578) );
  NAND2_X1 U643 ( .A1(G68), .A2(n647), .ZN(n577) );
  NAND2_X1 U644 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n583) );
  NAND2_X1 U646 ( .A1(n649), .A2(G56), .ZN(n581) );
  XOR2_X1 U647 ( .A(KEYINPUT14), .B(n581), .Z(n582) );
  NOR2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n585) );
  NAND2_X1 U649 ( .A1(n657), .A2(G43), .ZN(n584) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n969) );
  INV_X1 U651 ( .A(G860), .ZN(n614) );
  OR2_X1 U652 ( .A1(n969), .A2(n614), .ZN(G153) );
  NAND2_X1 U653 ( .A1(G90), .A2(n653), .ZN(n587) );
  NAND2_X1 U654 ( .A1(G77), .A2(n647), .ZN(n586) );
  NAND2_X1 U655 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U656 ( .A(KEYINPUT9), .B(n588), .ZN(n592) );
  NAND2_X1 U657 ( .A1(G64), .A2(n649), .ZN(n590) );
  NAND2_X1 U658 ( .A1(G52), .A2(n657), .ZN(n589) );
  AND2_X1 U659 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U660 ( .A1(n592), .A2(n591), .ZN(G301) );
  NAND2_X1 U661 ( .A1(G868), .A2(G301), .ZN(n593) );
  XNOR2_X1 U662 ( .A(n593), .B(KEYINPUT68), .ZN(n603) );
  INV_X1 U663 ( .A(G868), .ZN(n660) );
  NAND2_X1 U664 ( .A1(G54), .A2(n657), .ZN(n600) );
  NAND2_X1 U665 ( .A1(G79), .A2(n647), .ZN(n595) );
  NAND2_X1 U666 ( .A1(G66), .A2(n649), .ZN(n594) );
  NAND2_X1 U667 ( .A1(n595), .A2(n594), .ZN(n598) );
  NAND2_X1 U668 ( .A1(G92), .A2(n653), .ZN(n596) );
  XNOR2_X1 U669 ( .A(KEYINPUT69), .B(n596), .ZN(n597) );
  NOR2_X1 U670 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U671 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U672 ( .A(n601), .B(KEYINPUT15), .ZN(n882) );
  INV_X1 U673 ( .A(n882), .ZN(n972) );
  NAND2_X1 U674 ( .A1(n660), .A2(n972), .ZN(n602) );
  NAND2_X1 U675 ( .A1(n603), .A2(n602), .ZN(G284) );
  NAND2_X1 U676 ( .A1(G91), .A2(n653), .ZN(n605) );
  NAND2_X1 U677 ( .A1(G78), .A2(n647), .ZN(n604) );
  NAND2_X1 U678 ( .A1(n605), .A2(n604), .ZN(n609) );
  NAND2_X1 U679 ( .A1(G65), .A2(n649), .ZN(n607) );
  NAND2_X1 U680 ( .A1(G53), .A2(n657), .ZN(n606) );
  NAND2_X1 U681 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U682 ( .A1(n609), .A2(n608), .ZN(n610) );
  XOR2_X1 U683 ( .A(KEYINPUT66), .B(n610), .Z(G299) );
  NOR2_X1 U684 ( .A1(G299), .A2(G868), .ZN(n611) );
  XOR2_X1 U685 ( .A(KEYINPUT71), .B(n611), .Z(n613) );
  NOR2_X1 U686 ( .A1(G286), .A2(n660), .ZN(n612) );
  NOR2_X1 U687 ( .A1(n613), .A2(n612), .ZN(G297) );
  NAND2_X1 U688 ( .A1(n614), .A2(G559), .ZN(n615) );
  NAND2_X1 U689 ( .A1(n615), .A2(n882), .ZN(n616) );
  XNOR2_X1 U690 ( .A(n616), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U691 ( .A1(G868), .A2(n969), .ZN(n619) );
  NAND2_X1 U692 ( .A1(n882), .A2(G868), .ZN(n617) );
  NOR2_X1 U693 ( .A1(G559), .A2(n617), .ZN(n618) );
  NOR2_X1 U694 ( .A1(n619), .A2(n618), .ZN(G282) );
  NAND2_X1 U695 ( .A1(G99), .A2(n865), .ZN(n621) );
  NAND2_X1 U696 ( .A1(G135), .A2(n516), .ZN(n620) );
  NAND2_X1 U697 ( .A1(n621), .A2(n620), .ZN(n627) );
  NAND2_X1 U698 ( .A1(G123), .A2(n869), .ZN(n622) );
  XNOR2_X1 U699 ( .A(n622), .B(KEYINPUT18), .ZN(n625) );
  NAND2_X1 U700 ( .A1(n870), .A2(G111), .ZN(n623) );
  XNOR2_X1 U701 ( .A(n623), .B(KEYINPUT72), .ZN(n624) );
  NAND2_X1 U702 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U703 ( .A1(n627), .A2(n626), .ZN(n931) );
  XNOR2_X1 U704 ( .A(G2096), .B(n931), .ZN(n629) );
  INV_X1 U705 ( .A(G2100), .ZN(n628) );
  NAND2_X1 U706 ( .A1(n629), .A2(n628), .ZN(G156) );
  NAND2_X1 U707 ( .A1(G93), .A2(n653), .ZN(n630) );
  XNOR2_X1 U708 ( .A(n630), .B(KEYINPUT74), .ZN(n637) );
  NAND2_X1 U709 ( .A1(G80), .A2(n647), .ZN(n632) );
  NAND2_X1 U710 ( .A1(G55), .A2(n657), .ZN(n631) );
  NAND2_X1 U711 ( .A1(n632), .A2(n631), .ZN(n635) );
  NAND2_X1 U712 ( .A1(G67), .A2(n649), .ZN(n633) );
  XNOR2_X1 U713 ( .A(KEYINPUT75), .B(n633), .ZN(n634) );
  NOR2_X1 U714 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U715 ( .A1(n637), .A2(n636), .ZN(n664) );
  NAND2_X1 U716 ( .A1(n882), .A2(G559), .ZN(n671) );
  XOR2_X1 U717 ( .A(KEYINPUT73), .B(n969), .Z(n638) );
  XNOR2_X1 U718 ( .A(n671), .B(n638), .ZN(n639) );
  NOR2_X1 U719 ( .A1(G860), .A2(n639), .ZN(n640) );
  XOR2_X1 U720 ( .A(n664), .B(n640), .Z(G145) );
  NAND2_X1 U721 ( .A1(G49), .A2(n657), .ZN(n643) );
  NAND2_X1 U722 ( .A1(G87), .A2(n641), .ZN(n642) );
  NAND2_X1 U723 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U724 ( .A1(n649), .A2(n644), .ZN(n646) );
  NAND2_X1 U725 ( .A1(G651), .A2(G74), .ZN(n645) );
  NAND2_X1 U726 ( .A1(n646), .A2(n645), .ZN(G288) );
  NAND2_X1 U727 ( .A1(G73), .A2(n647), .ZN(n648) );
  XOR2_X1 U728 ( .A(KEYINPUT2), .B(n648), .Z(n652) );
  NAND2_X1 U729 ( .A1(n649), .A2(G61), .ZN(n650) );
  XOR2_X1 U730 ( .A(KEYINPUT76), .B(n650), .Z(n651) );
  NOR2_X1 U731 ( .A1(n652), .A2(n651), .ZN(n655) );
  NAND2_X1 U732 ( .A1(n653), .A2(G86), .ZN(n654) );
  NAND2_X1 U733 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U734 ( .A(n656), .B(KEYINPUT77), .ZN(n659) );
  NAND2_X1 U735 ( .A1(G48), .A2(n657), .ZN(n658) );
  NAND2_X1 U736 ( .A1(n659), .A2(n658), .ZN(G305) );
  AND2_X1 U737 ( .A1(n660), .A2(n664), .ZN(n661) );
  XNOR2_X1 U738 ( .A(n661), .B(KEYINPUT83), .ZN(n674) );
  XNOR2_X1 U739 ( .A(KEYINPUT81), .B(KEYINPUT82), .ZN(n663) );
  XNOR2_X1 U740 ( .A(G288), .B(KEYINPUT19), .ZN(n662) );
  XNOR2_X1 U741 ( .A(n663), .B(n662), .ZN(n667) );
  XNOR2_X1 U742 ( .A(G299), .B(G290), .ZN(n665) );
  XNOR2_X1 U743 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U744 ( .A(n667), .B(n666), .ZN(n669) );
  XNOR2_X1 U745 ( .A(n969), .B(G303), .ZN(n668) );
  XNOR2_X1 U746 ( .A(n669), .B(n668), .ZN(n670) );
  XOR2_X1 U747 ( .A(n670), .B(G305), .Z(n885) );
  XOR2_X1 U748 ( .A(n885), .B(n671), .Z(n672) );
  NAND2_X1 U749 ( .A1(G868), .A2(n672), .ZN(n673) );
  NAND2_X1 U750 ( .A1(n674), .A2(n673), .ZN(G295) );
  NAND2_X1 U751 ( .A1(G2084), .A2(G2078), .ZN(n675) );
  XOR2_X1 U752 ( .A(KEYINPUT20), .B(n675), .Z(n676) );
  NAND2_X1 U753 ( .A1(G2090), .A2(n676), .ZN(n677) );
  XNOR2_X1 U754 ( .A(KEYINPUT21), .B(n677), .ZN(n678) );
  NAND2_X1 U755 ( .A1(n678), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U756 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U757 ( .A1(G220), .A2(G219), .ZN(n679) );
  XOR2_X1 U758 ( .A(KEYINPUT22), .B(n679), .Z(n680) );
  NOR2_X1 U759 ( .A1(G218), .A2(n680), .ZN(n681) );
  NAND2_X1 U760 ( .A1(G96), .A2(n681), .ZN(n839) );
  NAND2_X1 U761 ( .A1(G2106), .A2(n839), .ZN(n682) );
  XOR2_X1 U762 ( .A(KEYINPUT84), .B(n682), .Z(n687) );
  NOR2_X1 U763 ( .A1(G236), .A2(G238), .ZN(n684) );
  NOR2_X1 U764 ( .A1(G235), .A2(G237), .ZN(n683) );
  NAND2_X1 U765 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U766 ( .A(KEYINPUT85), .B(n685), .Z(n840) );
  AND2_X1 U767 ( .A1(n840), .A2(G567), .ZN(n686) );
  NOR2_X1 U768 ( .A1(n687), .A2(n686), .ZN(G319) );
  INV_X1 U769 ( .A(G319), .ZN(n910) );
  NAND2_X1 U770 ( .A1(G661), .A2(G483), .ZN(n688) );
  NOR2_X1 U771 ( .A1(n910), .A2(n688), .ZN(n836) );
  NAND2_X1 U772 ( .A1(G36), .A2(n836), .ZN(n689) );
  XNOR2_X1 U773 ( .A(n689), .B(KEYINPUT86), .ZN(G176) );
  INV_X1 U774 ( .A(G1384), .ZN(n714) );
  AND2_X1 U775 ( .A1(n716), .A2(n714), .ZN(n690) );
  NAND2_X1 U776 ( .A1(G160), .A2(G40), .ZN(n713) );
  NOR2_X1 U777 ( .A1(n690), .A2(n713), .ZN(n827) );
  XNOR2_X1 U778 ( .A(G1986), .B(G290), .ZN(n978) );
  NAND2_X1 U779 ( .A1(n827), .A2(n978), .ZN(n712) );
  NAND2_X1 U780 ( .A1(G141), .A2(n516), .ZN(n692) );
  NAND2_X1 U781 ( .A1(G117), .A2(n870), .ZN(n691) );
  NAND2_X1 U782 ( .A1(n692), .A2(n691), .ZN(n695) );
  NAND2_X1 U783 ( .A1(n865), .A2(G105), .ZN(n693) );
  XOR2_X1 U784 ( .A(KEYINPUT38), .B(n693), .Z(n694) );
  NOR2_X1 U785 ( .A1(n695), .A2(n694), .ZN(n697) );
  NAND2_X1 U786 ( .A1(n869), .A2(G129), .ZN(n696) );
  NAND2_X1 U787 ( .A1(n697), .A2(n696), .ZN(n855) );
  NAND2_X1 U788 ( .A1(G1996), .A2(n855), .ZN(n698) );
  XNOR2_X1 U789 ( .A(n698), .B(KEYINPUT92), .ZN(n709) );
  NAND2_X1 U790 ( .A1(G107), .A2(n870), .ZN(n699) );
  XOR2_X1 U791 ( .A(KEYINPUT89), .B(n699), .Z(n701) );
  NAND2_X1 U792 ( .A1(n869), .A2(G119), .ZN(n700) );
  NAND2_X1 U793 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U794 ( .A(KEYINPUT90), .B(n702), .ZN(n705) );
  NAND2_X1 U795 ( .A1(G95), .A2(n865), .ZN(n703) );
  XNOR2_X1 U796 ( .A(KEYINPUT91), .B(n703), .ZN(n704) );
  NOR2_X1 U797 ( .A1(n705), .A2(n704), .ZN(n707) );
  NAND2_X1 U798 ( .A1(n516), .A2(G131), .ZN(n706) );
  NAND2_X1 U799 ( .A1(n707), .A2(n706), .ZN(n876) );
  NAND2_X1 U800 ( .A1(G1991), .A2(n876), .ZN(n708) );
  NAND2_X1 U801 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U802 ( .A(KEYINPUT93), .B(n710), .ZN(n935) );
  INV_X1 U803 ( .A(n935), .ZN(n711) );
  NAND2_X1 U804 ( .A1(n711), .A2(n827), .ZN(n816) );
  NAND2_X1 U805 ( .A1(n712), .A2(n816), .ZN(n804) );
  INV_X1 U806 ( .A(n713), .ZN(n715) );
  AND2_X1 U807 ( .A1(n715), .A2(n714), .ZN(n717) );
  NOR2_X1 U808 ( .A1(G2084), .A2(n769), .ZN(n753) );
  NAND2_X1 U809 ( .A1(G8), .A2(n753), .ZN(n767) );
  NAND2_X1 U810 ( .A1(G8), .A2(n769), .ZN(n798) );
  NOR2_X1 U811 ( .A1(G1966), .A2(n798), .ZN(n765) );
  INV_X2 U812 ( .A(n769), .ZN(n744) );
  XNOR2_X1 U813 ( .A(n718), .B(KEYINPUT26), .ZN(n719) );
  INV_X1 U814 ( .A(n719), .ZN(n720) );
  NAND2_X1 U815 ( .A1(n720), .A2(n517), .ZN(n721) );
  NOR2_X2 U816 ( .A1(n969), .A2(n721), .ZN(n728) );
  NAND2_X1 U817 ( .A1(n728), .A2(n882), .ZN(n726) );
  INV_X1 U818 ( .A(G1348), .ZN(n993) );
  NOR2_X1 U819 ( .A1(n744), .A2(n993), .ZN(n722) );
  XNOR2_X1 U820 ( .A(n722), .B(KEYINPUT97), .ZN(n724) );
  NAND2_X1 U821 ( .A1(n744), .A2(G2067), .ZN(n723) );
  NAND2_X1 U822 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U823 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U824 ( .A(n727), .B(KEYINPUT98), .ZN(n730) );
  OR2_X1 U825 ( .A1(n728), .A2(n882), .ZN(n729) );
  NAND2_X1 U826 ( .A1(n730), .A2(n729), .ZN(n736) );
  NAND2_X1 U827 ( .A1(G2072), .A2(n744), .ZN(n731) );
  XOR2_X1 U828 ( .A(KEYINPUT95), .B(n731), .Z(n732) );
  XNOR2_X1 U829 ( .A(KEYINPUT27), .B(n732), .ZN(n734) );
  INV_X1 U830 ( .A(G1956), .ZN(n995) );
  NOR2_X1 U831 ( .A1(n744), .A2(n995), .ZN(n733) );
  NOR2_X1 U832 ( .A1(n734), .A2(n733), .ZN(n738) );
  INV_X1 U833 ( .A(G299), .ZN(n737) );
  NAND2_X1 U834 ( .A1(n738), .A2(n737), .ZN(n735) );
  NAND2_X1 U835 ( .A1(n736), .A2(n735), .ZN(n742) );
  NOR2_X1 U836 ( .A1(n738), .A2(n737), .ZN(n740) );
  XOR2_X1 U837 ( .A(KEYINPUT28), .B(KEYINPUT96), .Z(n739) );
  XNOR2_X1 U838 ( .A(n740), .B(n739), .ZN(n741) );
  NAND2_X1 U839 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U840 ( .A(KEYINPUT29), .B(n743), .ZN(n749) );
  NAND2_X1 U841 ( .A1(G1961), .A2(n769), .ZN(n746) );
  XOR2_X1 U842 ( .A(KEYINPUT25), .B(G2078), .Z(n944) );
  NAND2_X1 U843 ( .A1(n744), .A2(n944), .ZN(n745) );
  NAND2_X1 U844 ( .A1(n746), .A2(n745), .ZN(n751) );
  NOR2_X1 U845 ( .A1(G301), .A2(n751), .ZN(n747) );
  XNOR2_X1 U846 ( .A(n747), .B(KEYINPUT94), .ZN(n748) );
  XNOR2_X1 U847 ( .A(n750), .B(KEYINPUT99), .ZN(n762) );
  NAND2_X1 U848 ( .A1(G301), .A2(n751), .ZN(n752) );
  XOR2_X1 U849 ( .A(KEYINPUT100), .B(n752), .Z(n758) );
  NOR2_X1 U850 ( .A1(n765), .A2(n753), .ZN(n754) );
  NAND2_X1 U851 ( .A1(G8), .A2(n754), .ZN(n755) );
  XNOR2_X1 U852 ( .A(KEYINPUT30), .B(n755), .ZN(n756) );
  NOR2_X1 U853 ( .A1(G168), .A2(n756), .ZN(n757) );
  NOR2_X1 U854 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U855 ( .A(n759), .B(KEYINPUT101), .ZN(n760) );
  XNOR2_X1 U856 ( .A(n760), .B(KEYINPUT31), .ZN(n761) );
  NAND2_X1 U857 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U858 ( .A(n763), .B(KEYINPUT102), .ZN(n768) );
  INV_X1 U859 ( .A(n768), .ZN(n764) );
  NOR2_X1 U860 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U861 ( .A1(n767), .A2(n766), .ZN(n779) );
  NAND2_X1 U862 ( .A1(n768), .A2(G286), .ZN(n774) );
  NOR2_X1 U863 ( .A1(G1971), .A2(n798), .ZN(n771) );
  NOR2_X1 U864 ( .A1(G2090), .A2(n769), .ZN(n770) );
  NOR2_X1 U865 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U866 ( .A1(n772), .A2(G303), .ZN(n773) );
  NAND2_X1 U867 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U868 ( .A1(n775), .A2(G8), .ZN(n777) );
  XOR2_X1 U869 ( .A(KEYINPUT32), .B(KEYINPUT103), .Z(n776) );
  XNOR2_X1 U870 ( .A(n777), .B(n776), .ZN(n778) );
  NAND2_X1 U871 ( .A1(n779), .A2(n778), .ZN(n794) );
  NOR2_X1 U872 ( .A1(G1976), .A2(G288), .ZN(n785) );
  NOR2_X1 U873 ( .A1(G303), .A2(G1971), .ZN(n780) );
  NOR2_X1 U874 ( .A1(n785), .A2(n780), .ZN(n982) );
  INV_X1 U875 ( .A(KEYINPUT33), .ZN(n781) );
  AND2_X1 U876 ( .A1(n982), .A2(n781), .ZN(n782) );
  AND2_X1 U877 ( .A1(n794), .A2(n782), .ZN(n791) );
  INV_X1 U878 ( .A(n798), .ZN(n783) );
  NAND2_X1 U879 ( .A1(G1976), .A2(G288), .ZN(n975) );
  AND2_X1 U880 ( .A1(n783), .A2(n975), .ZN(n784) );
  NOR2_X1 U881 ( .A1(KEYINPUT33), .A2(n784), .ZN(n788) );
  NAND2_X1 U882 ( .A1(n785), .A2(KEYINPUT33), .ZN(n786) );
  NOR2_X1 U883 ( .A1(n798), .A2(n786), .ZN(n787) );
  NOR2_X1 U884 ( .A1(n788), .A2(n787), .ZN(n789) );
  XOR2_X1 U885 ( .A(G1981), .B(G305), .Z(n964) );
  NAND2_X1 U886 ( .A1(n789), .A2(n964), .ZN(n790) );
  NOR2_X1 U887 ( .A1(n791), .A2(n790), .ZN(n802) );
  NOR2_X1 U888 ( .A1(G2090), .A2(G303), .ZN(n792) );
  NAND2_X1 U889 ( .A1(G8), .A2(n792), .ZN(n793) );
  NAND2_X1 U890 ( .A1(n794), .A2(n793), .ZN(n795) );
  NAND2_X1 U891 ( .A1(n795), .A2(n798), .ZN(n800) );
  NOR2_X1 U892 ( .A1(G1981), .A2(G305), .ZN(n796) );
  XOR2_X1 U893 ( .A(n796), .B(KEYINPUT24), .Z(n797) );
  OR2_X1 U894 ( .A1(n798), .A2(n797), .ZN(n799) );
  NAND2_X1 U895 ( .A1(n800), .A2(n799), .ZN(n801) );
  NOR2_X1 U896 ( .A1(n802), .A2(n801), .ZN(n803) );
  NOR2_X1 U897 ( .A1(n804), .A2(n803), .ZN(n815) );
  NAND2_X1 U898 ( .A1(G104), .A2(n865), .ZN(n806) );
  NAND2_X1 U899 ( .A1(G140), .A2(n516), .ZN(n805) );
  NAND2_X1 U900 ( .A1(n806), .A2(n805), .ZN(n807) );
  XNOR2_X1 U901 ( .A(KEYINPUT34), .B(n807), .ZN(n813) );
  NAND2_X1 U902 ( .A1(n869), .A2(G128), .ZN(n809) );
  NAND2_X1 U903 ( .A1(G116), .A2(n870), .ZN(n808) );
  NAND2_X1 U904 ( .A1(n809), .A2(n808), .ZN(n810) );
  XOR2_X1 U905 ( .A(KEYINPUT35), .B(n810), .Z(n811) );
  XNOR2_X1 U906 ( .A(KEYINPUT88), .B(n811), .ZN(n812) );
  NOR2_X1 U907 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U908 ( .A(KEYINPUT36), .B(n814), .ZN(n879) );
  XNOR2_X1 U909 ( .A(G2067), .B(KEYINPUT37), .ZN(n824) );
  NOR2_X1 U910 ( .A1(n879), .A2(n824), .ZN(n928) );
  NAND2_X1 U911 ( .A1(n827), .A2(n928), .ZN(n822) );
  NAND2_X1 U912 ( .A1(n815), .A2(n822), .ZN(n830) );
  NOR2_X1 U913 ( .A1(G1996), .A2(n855), .ZN(n921) );
  INV_X1 U914 ( .A(n816), .ZN(n819) );
  NOR2_X1 U915 ( .A1(G1986), .A2(G290), .ZN(n817) );
  NOR2_X1 U916 ( .A1(G1991), .A2(n876), .ZN(n932) );
  NOR2_X1 U917 ( .A1(n817), .A2(n932), .ZN(n818) );
  NOR2_X1 U918 ( .A1(n819), .A2(n818), .ZN(n820) );
  NOR2_X1 U919 ( .A1(n921), .A2(n820), .ZN(n821) );
  XNOR2_X1 U920 ( .A(n821), .B(KEYINPUT39), .ZN(n823) );
  NAND2_X1 U921 ( .A1(n823), .A2(n822), .ZN(n825) );
  NAND2_X1 U922 ( .A1(n879), .A2(n824), .ZN(n925) );
  NAND2_X1 U923 ( .A1(n825), .A2(n925), .ZN(n826) );
  NAND2_X1 U924 ( .A1(n827), .A2(n826), .ZN(n828) );
  XNOR2_X1 U925 ( .A(n828), .B(KEYINPUT104), .ZN(n829) );
  NAND2_X1 U926 ( .A1(n830), .A2(n829), .ZN(n831) );
  XNOR2_X1 U927 ( .A(KEYINPUT40), .B(n831), .ZN(G329) );
  NAND2_X1 U928 ( .A1(n832), .A2(G2106), .ZN(n833) );
  XNOR2_X1 U929 ( .A(n833), .B(KEYINPUT106), .ZN(G217) );
  NAND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n834) );
  XNOR2_X1 U931 ( .A(KEYINPUT107), .B(n834), .ZN(n835) );
  NAND2_X1 U932 ( .A1(n835), .A2(G661), .ZN(G259) );
  NAND2_X1 U933 ( .A1(G3), .A2(G1), .ZN(n837) );
  NAND2_X1 U934 ( .A1(n837), .A2(n836), .ZN(n838) );
  XNOR2_X1 U935 ( .A(n838), .B(KEYINPUT108), .ZN(G188) );
  XNOR2_X1 U936 ( .A(G96), .B(KEYINPUT109), .ZN(G221) );
  NOR2_X1 U938 ( .A1(n840), .A2(n839), .ZN(G325) );
  INV_X1 U939 ( .A(G325), .ZN(G261) );
  NAND2_X1 U940 ( .A1(G124), .A2(n869), .ZN(n841) );
  XNOR2_X1 U941 ( .A(n841), .B(KEYINPUT44), .ZN(n843) );
  NAND2_X1 U942 ( .A1(n865), .A2(G100), .ZN(n842) );
  NAND2_X1 U943 ( .A1(n843), .A2(n842), .ZN(n847) );
  NAND2_X1 U944 ( .A1(G136), .A2(n516), .ZN(n845) );
  NAND2_X1 U945 ( .A1(G112), .A2(n870), .ZN(n844) );
  NAND2_X1 U946 ( .A1(n845), .A2(n844), .ZN(n846) );
  NOR2_X1 U947 ( .A1(n847), .A2(n846), .ZN(G162) );
  NAND2_X1 U948 ( .A1(n869), .A2(G130), .ZN(n849) );
  NAND2_X1 U949 ( .A1(G118), .A2(n870), .ZN(n848) );
  NAND2_X1 U950 ( .A1(n849), .A2(n848), .ZN(n854) );
  NAND2_X1 U951 ( .A1(G106), .A2(n865), .ZN(n851) );
  NAND2_X1 U952 ( .A1(G142), .A2(n516), .ZN(n850) );
  NAND2_X1 U953 ( .A1(n851), .A2(n850), .ZN(n852) );
  XOR2_X1 U954 ( .A(KEYINPUT45), .B(n852), .Z(n853) );
  NOR2_X1 U955 ( .A1(n854), .A2(n853), .ZN(n864) );
  XNOR2_X1 U956 ( .A(G164), .B(n931), .ZN(n862) );
  XNOR2_X1 U957 ( .A(KEYINPUT114), .B(KEYINPUT113), .ZN(n857) );
  XNOR2_X1 U958 ( .A(n855), .B(KEYINPUT48), .ZN(n856) );
  XNOR2_X1 U959 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U960 ( .A(n858), .B(KEYINPUT46), .Z(n860) );
  XNOR2_X1 U961 ( .A(G160), .B(G162), .ZN(n859) );
  XNOR2_X1 U962 ( .A(n860), .B(n859), .ZN(n861) );
  XNOR2_X1 U963 ( .A(n862), .B(n861), .ZN(n863) );
  XNOR2_X1 U964 ( .A(n864), .B(n863), .ZN(n878) );
  NAND2_X1 U965 ( .A1(G103), .A2(n865), .ZN(n868) );
  NAND2_X1 U966 ( .A1(G139), .A2(n516), .ZN(n867) );
  NAND2_X1 U967 ( .A1(n868), .A2(n867), .ZN(n875) );
  NAND2_X1 U968 ( .A1(n869), .A2(G127), .ZN(n872) );
  NAND2_X1 U969 ( .A1(G115), .A2(n870), .ZN(n871) );
  NAND2_X1 U970 ( .A1(n872), .A2(n871), .ZN(n873) );
  XOR2_X1 U971 ( .A(KEYINPUT47), .B(n873), .Z(n874) );
  NOR2_X1 U972 ( .A1(n875), .A2(n874), .ZN(n916) );
  XNOR2_X1 U973 ( .A(n876), .B(n916), .ZN(n877) );
  XNOR2_X1 U974 ( .A(n878), .B(n877), .ZN(n880) );
  XNOR2_X1 U975 ( .A(n880), .B(n879), .ZN(n881) );
  NOR2_X1 U976 ( .A1(G37), .A2(n881), .ZN(G395) );
  INV_X1 U977 ( .A(G301), .ZN(G171) );
  XOR2_X1 U978 ( .A(KEYINPUT115), .B(G286), .Z(n884) );
  XNOR2_X1 U979 ( .A(G171), .B(n882), .ZN(n883) );
  XNOR2_X1 U980 ( .A(n884), .B(n883), .ZN(n886) );
  XNOR2_X1 U981 ( .A(n886), .B(n885), .ZN(n887) );
  NOR2_X1 U982 ( .A1(G37), .A2(n887), .ZN(G397) );
  XOR2_X1 U983 ( .A(KEYINPUT111), .B(G1981), .Z(n889) );
  XNOR2_X1 U984 ( .A(G1966), .B(G1956), .ZN(n888) );
  XNOR2_X1 U985 ( .A(n889), .B(n888), .ZN(n890) );
  XOR2_X1 U986 ( .A(n890), .B(KEYINPUT41), .Z(n892) );
  XNOR2_X1 U987 ( .A(G1996), .B(G1991), .ZN(n891) );
  XNOR2_X1 U988 ( .A(n892), .B(n891), .ZN(n896) );
  XOR2_X1 U989 ( .A(G1986), .B(G1976), .Z(n894) );
  XNOR2_X1 U990 ( .A(G1961), .B(G1971), .ZN(n893) );
  XNOR2_X1 U991 ( .A(n894), .B(n893), .ZN(n895) );
  XOR2_X1 U992 ( .A(n896), .B(n895), .Z(n898) );
  XNOR2_X1 U993 ( .A(KEYINPUT112), .B(G2474), .ZN(n897) );
  XNOR2_X1 U994 ( .A(n898), .B(n897), .ZN(G229) );
  XOR2_X1 U995 ( .A(G2096), .B(KEYINPUT43), .Z(n900) );
  XNOR2_X1 U996 ( .A(G2090), .B(KEYINPUT110), .ZN(n899) );
  XNOR2_X1 U997 ( .A(n900), .B(n899), .ZN(n901) );
  XOR2_X1 U998 ( .A(n901), .B(G2678), .Z(n903) );
  XNOR2_X1 U999 ( .A(G2072), .B(G2067), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(n903), .B(n902), .ZN(n907) );
  XOR2_X1 U1001 ( .A(KEYINPUT42), .B(G2100), .Z(n905) );
  XNOR2_X1 U1002 ( .A(G2084), .B(G2078), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(n907), .B(n906), .ZN(G227) );
  NOR2_X1 U1005 ( .A1(G229), .A2(G227), .ZN(n908) );
  XNOR2_X1 U1006 ( .A(KEYINPUT49), .B(n908), .ZN(n909) );
  NOR2_X1 U1007 ( .A1(G397), .A2(n909), .ZN(n913) );
  NOR2_X1 U1008 ( .A1(G401), .A2(n910), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(n911), .B(KEYINPUT116), .ZN(n912) );
  NAND2_X1 U1010 ( .A1(n913), .A2(n912), .ZN(n914) );
  NOR2_X1 U1011 ( .A1(G395), .A2(n914), .ZN(n915) );
  XNOR2_X1 U1012 ( .A(KEYINPUT117), .B(n915), .ZN(G225) );
  INV_X1 U1013 ( .A(G225), .ZN(G308) );
  INV_X1 U1014 ( .A(G303), .ZN(G166) );
  XOR2_X1 U1015 ( .A(G2072), .B(n916), .Z(n918) );
  XOR2_X1 U1016 ( .A(G164), .B(G2078), .Z(n917) );
  NOR2_X1 U1017 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1018 ( .A(KEYINPUT50), .B(n919), .ZN(n930) );
  XOR2_X1 U1019 ( .A(G160), .B(G2084), .Z(n924) );
  XOR2_X1 U1020 ( .A(G2090), .B(G162), .Z(n920) );
  NOR2_X1 U1021 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1022 ( .A(KEYINPUT51), .B(n922), .ZN(n923) );
  NOR2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n926) );
  NAND2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n927) );
  NOR2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1026 ( .A1(n930), .A2(n929), .ZN(n937) );
  NOR2_X1 U1027 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1028 ( .A(n933), .B(KEYINPUT118), .ZN(n934) );
  NAND2_X1 U1029 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1030 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1031 ( .A(KEYINPUT52), .B(n938), .ZN(n940) );
  INV_X1 U1032 ( .A(KEYINPUT55), .ZN(n939) );
  NAND2_X1 U1033 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1034 ( .A1(n941), .A2(G29), .ZN(n942) );
  XNOR2_X1 U1035 ( .A(n942), .B(KEYINPUT119), .ZN(n963) );
  XNOR2_X1 U1036 ( .A(G2090), .B(G35), .ZN(n956) );
  XOR2_X1 U1037 ( .A(G1991), .B(G25), .Z(n943) );
  NAND2_X1 U1038 ( .A1(n943), .A2(G28), .ZN(n953) );
  XNOR2_X1 U1039 ( .A(n944), .B(G27), .ZN(n946) );
  XNOR2_X1 U1040 ( .A(G32), .B(G1996), .ZN(n945) );
  NOR2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1042 ( .A(KEYINPUT120), .B(n947), .ZN(n951) );
  XNOR2_X1 U1043 ( .A(G2072), .B(G33), .ZN(n949) );
  XNOR2_X1 U1044 ( .A(G2067), .B(G26), .ZN(n948) );
  NOR2_X1 U1045 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1046 ( .A1(n951), .A2(n950), .ZN(n952) );
  NOR2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(KEYINPUT53), .B(n954), .ZN(n955) );
  NOR2_X1 U1049 ( .A1(n956), .A2(n955), .ZN(n959) );
  XOR2_X1 U1050 ( .A(G2084), .B(G34), .Z(n957) );
  XNOR2_X1 U1051 ( .A(KEYINPUT54), .B(n957), .ZN(n958) );
  NAND2_X1 U1052 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1053 ( .A(KEYINPUT55), .B(n960), .ZN(n961) );
  NOR2_X1 U1054 ( .A1(n961), .A2(G29), .ZN(n962) );
  NOR2_X1 U1055 ( .A1(n963), .A2(n962), .ZN(n992) );
  XNOR2_X1 U1056 ( .A(KEYINPUT121), .B(KEYINPUT122), .ZN(n968) );
  XNOR2_X1 U1057 ( .A(G1966), .B(G168), .ZN(n965) );
  NAND2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1059 ( .A(n966), .B(KEYINPUT57), .ZN(n967) );
  XNOR2_X1 U1060 ( .A(n968), .B(n967), .ZN(n987) );
  XNOR2_X1 U1061 ( .A(n969), .B(G1341), .ZN(n971) );
  XNOR2_X1 U1062 ( .A(G299), .B(G1956), .ZN(n970) );
  NOR2_X1 U1063 ( .A1(n971), .A2(n970), .ZN(n980) );
  XNOR2_X1 U1064 ( .A(G301), .B(G1961), .ZN(n974) );
  XNOR2_X1 U1065 ( .A(n972), .B(G1348), .ZN(n973) );
  NOR2_X1 U1066 ( .A1(n974), .A2(n973), .ZN(n976) );
  NAND2_X1 U1067 ( .A1(n976), .A2(n975), .ZN(n977) );
  NOR2_X1 U1068 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1069 ( .A1(n980), .A2(n979), .ZN(n984) );
  NAND2_X1 U1070 ( .A1(G303), .A2(G1971), .ZN(n981) );
  NAND2_X1 U1071 ( .A1(n982), .A2(n981), .ZN(n983) );
  NOR2_X1 U1072 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1073 ( .A(n985), .B(KEYINPUT123), .ZN(n986) );
  NOR2_X1 U1074 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1075 ( .A(KEYINPUT124), .B(n988), .Z(n990) );
  XNOR2_X1 U1076 ( .A(G16), .B(KEYINPUT56), .ZN(n989) );
  NAND2_X1 U1077 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1078 ( .A1(n992), .A2(n991), .ZN(n1021) );
  XOR2_X1 U1079 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n1016) );
  XOR2_X1 U1080 ( .A(G1966), .B(G21), .Z(n1005) );
  XNOR2_X1 U1081 ( .A(G4), .B(KEYINPUT59), .ZN(n994) );
  XNOR2_X1 U1082 ( .A(n994), .B(n993), .ZN(n1002) );
  XNOR2_X1 U1083 ( .A(G20), .B(n995), .ZN(n999) );
  XNOR2_X1 U1084 ( .A(G1341), .B(G19), .ZN(n997) );
  XNOR2_X1 U1085 ( .A(G1981), .B(G6), .ZN(n996) );
  NOR2_X1 U1086 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1087 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1088 ( .A(KEYINPUT125), .B(n1000), .Z(n1001) );
  NOR2_X1 U1089 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1090 ( .A(KEYINPUT60), .B(n1003), .ZN(n1004) );
  NAND2_X1 U1091 ( .A1(n1005), .A2(n1004), .ZN(n1012) );
  XNOR2_X1 U1092 ( .A(G1971), .B(G22), .ZN(n1007) );
  XNOR2_X1 U1093 ( .A(G23), .B(G1976), .ZN(n1006) );
  NOR2_X1 U1094 ( .A1(n1007), .A2(n1006), .ZN(n1009) );
  XOR2_X1 U1095 ( .A(G1986), .B(G24), .Z(n1008) );
  NAND2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1097 ( .A(KEYINPUT58), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1098 ( .A1(n1012), .A2(n1011), .ZN(n1014) );
  XOR2_X1 U1099 ( .A(G1961), .B(G5), .Z(n1013) );
  NAND2_X1 U1100 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1101 ( .A(n1016), .B(n1015), .ZN(n1018) );
  INV_X1 U1102 ( .A(G16), .ZN(n1017) );
  NAND2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1104 ( .A1(G11), .A2(n1019), .ZN(n1020) );
  NOR2_X1 U1105 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1106 ( .A(n1022), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1107 ( .A(G311), .ZN(G150) );
endmodule

