//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 1 1 0 1 1 1 0 0 0 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 1 1 0 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:24 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047;
  INV_X1    g000(.A(KEYINPUT30), .ZN(new_n187));
  NAND2_X1  g001(.A1(KEYINPUT68), .A2(KEYINPUT11), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G134), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G137), .ZN(new_n191));
  OR2_X1    g005(.A1(KEYINPUT68), .A2(KEYINPUT11), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n189), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n190), .A2(G137), .ZN(new_n194));
  INV_X1    g008(.A(G137), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G134), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n194), .B1(new_n196), .B2(new_n188), .ZN(new_n197));
  OAI21_X1  g011(.A(G131), .B1(new_n193), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT69), .ZN(new_n199));
  NOR2_X1   g013(.A1(KEYINPUT68), .A2(KEYINPUT11), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n188), .B1(new_n196), .B2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n191), .A2(new_n189), .ZN(new_n202));
  INV_X1    g016(.A(G131), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n201), .A2(new_n202), .A3(new_n203), .A4(new_n194), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n198), .A2(new_n199), .A3(new_n204), .ZN(new_n205));
  OAI211_X1 g019(.A(KEYINPUT69), .B(G131), .C1(new_n193), .C2(new_n197), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT64), .ZN(new_n208));
  INV_X1    g022(.A(G143), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(KEYINPUT64), .A2(G143), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(G146), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(KEYINPUT67), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT67), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n210), .A2(new_n214), .A3(G146), .A4(new_n211), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n209), .A2(G146), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  AND2_X1   g031(.A1(KEYINPUT0), .A2(G128), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n213), .A2(new_n215), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G146), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT66), .B1(new_n220), .B2(G143), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n222), .A2(new_n209), .A3(G146), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  AND2_X1   g038(.A1(KEYINPUT64), .A2(G143), .ZN(new_n225));
  NOR2_X1   g039(.A1(KEYINPUT64), .A2(G143), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n220), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(KEYINPUT65), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT65), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n229), .B(new_n220), .C1(new_n225), .C2(new_n226), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n224), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g045(.A(KEYINPUT0), .B(G128), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n219), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n207), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n196), .A2(new_n194), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G131), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n204), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n224), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n210), .A2(new_n211), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n229), .B1(new_n239), .B2(new_n220), .ZN(new_n240));
  INV_X1    g054(.A(new_n230), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n238), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G128), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n243), .B1(new_n217), .B2(KEYINPUT1), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n242), .A2(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n243), .A2(KEYINPUT1), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n213), .A2(new_n215), .A3(new_n217), .A4(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n237), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n187), .B1(new_n234), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G116), .ZN(new_n251));
  INV_X1    g065(.A(G119), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(G116), .A2(G119), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(KEYINPUT2), .B(G113), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n255), .A2(KEYINPUT70), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT70), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n253), .A2(new_n260), .A3(new_n254), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n258), .B1(new_n262), .B2(new_n257), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n232), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n242), .A2(new_n265), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n266), .A2(new_n219), .A3(new_n206), .A4(new_n205), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n248), .B1(new_n231), .B2(new_n244), .ZN(new_n268));
  INV_X1    g082(.A(new_n237), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n267), .A2(KEYINPUT30), .A3(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n250), .A2(new_n264), .A3(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT31), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n267), .A2(new_n263), .A3(new_n270), .ZN(new_n274));
  INV_X1    g088(.A(G101), .ZN(new_n275));
  OR2_X1    g089(.A1(KEYINPUT71), .A2(G237), .ZN(new_n276));
  NAND2_X1  g090(.A1(KEYINPUT71), .A2(G237), .ZN(new_n277));
  AOI21_X1  g091(.A(G953), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G210), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT27), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT26), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT27), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n278), .A2(new_n282), .A3(G210), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n280), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n281), .B1(new_n280), .B2(new_n283), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n275), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(new_n286), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n288), .A2(G101), .A3(new_n284), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n272), .A2(new_n273), .A3(new_n274), .A4(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT72), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n272), .A2(new_n274), .A3(new_n291), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(KEYINPUT31), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n294), .A2(KEYINPUT72), .A3(KEYINPUT31), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT28), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n274), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n264), .B1(new_n234), .B2(new_n249), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n298), .B1(new_n300), .B2(new_n274), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT73), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n299), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  AOI211_X1 g117(.A(KEYINPUT73), .B(new_n298), .C1(new_n300), .C2(new_n274), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n290), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n296), .A2(new_n297), .A3(new_n305), .ZN(new_n306));
  NOR2_X1   g120(.A1(G472), .A2(G902), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT32), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n291), .B1(new_n303), .B2(new_n304), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n272), .A2(new_n274), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(new_n290), .ZN(new_n314));
  AOI21_X1  g128(.A(KEYINPUT29), .B1(new_n311), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G902), .ZN(new_n316));
  AND3_X1   g130(.A1(new_n267), .A2(new_n263), .A3(new_n270), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n263), .B1(new_n267), .B2(new_n270), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT28), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT74), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n299), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n274), .A2(KEYINPUT74), .A3(new_n298), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n319), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n291), .A2(KEYINPUT29), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n316), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(G472), .B1(new_n315), .B2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n306), .A2(KEYINPUT32), .A3(new_n307), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n310), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n248), .A2(KEYINPUT79), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n216), .B1(new_n212), .B2(KEYINPUT67), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT79), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n330), .A2(new_n331), .A3(new_n215), .A4(new_n247), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n213), .A2(new_n215), .A3(new_n217), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n227), .A2(KEYINPUT1), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G128), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n329), .A2(new_n332), .A3(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(G107), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G104), .ZN(new_n339));
  INV_X1    g153(.A(G104), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G107), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n275), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT3), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n343), .A2(new_n338), .A3(G104), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n344), .A2(new_n341), .ZN(new_n345));
  OAI21_X1  g159(.A(KEYINPUT3), .B1(new_n340), .B2(G107), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n345), .A2(KEYINPUT78), .A3(new_n275), .A4(new_n346), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n346), .A2(new_n344), .A3(new_n275), .A4(new_n341), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT78), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n342), .B1(new_n347), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n337), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT10), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n346), .A2(new_n344), .A3(new_n341), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(G101), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT4), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n357), .B1(new_n347), .B2(new_n350), .ZN(new_n360));
  INV_X1    g174(.A(new_n356), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(new_n219), .A3(new_n266), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n268), .A2(KEYINPUT10), .A3(new_n351), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n354), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n207), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(G110), .B(G140), .ZN(new_n368));
  INV_X1    g182(.A(G227), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n369), .A2(G953), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n368), .B(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n354), .A2(new_n207), .A3(new_n363), .A4(new_n364), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n367), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n373), .ZN(new_n375));
  INV_X1    g189(.A(new_n342), .ZN(new_n376));
  INV_X1    g190(.A(new_n350), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n348), .A2(new_n349), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n379), .A2(new_n246), .A3(new_n248), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n207), .B1(new_n352), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(KEYINPUT81), .B1(new_n381), .B2(KEYINPUT12), .ZN(new_n382));
  AOI22_X1  g196(.A1(KEYINPUT79), .A2(new_n248), .B1(new_n333), .B2(new_n335), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n379), .B1(new_n383), .B2(new_n332), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n268), .A2(new_n351), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n366), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT81), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT12), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n382), .A2(new_n389), .ZN(new_n390));
  OAI211_X1 g204(.A(KEYINPUT12), .B(new_n366), .C1(new_n384), .C2(new_n385), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(KEYINPUT80), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT80), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n381), .A2(new_n393), .A3(KEYINPUT12), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n375), .B1(new_n390), .B2(new_n395), .ZN(new_n396));
  OAI211_X1 g210(.A(G469), .B(new_n374), .C1(new_n396), .C2(new_n372), .ZN(new_n397));
  INV_X1    g211(.A(G469), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n373), .A2(new_n372), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n399), .B1(new_n390), .B2(new_n395), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n372), .B1(new_n367), .B2(new_n373), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n398), .B(new_n316), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n398), .A2(new_n316), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n397), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(G214), .B1(G237), .B2(G902), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n406), .B(KEYINPUT82), .ZN(new_n407));
  OAI21_X1  g221(.A(G210), .B1(G237), .B2(G902), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(KEYINPUT4), .B1(new_n377), .B2(new_n378), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n358), .B1(new_n410), .B2(new_n356), .ZN(new_n411));
  INV_X1    g225(.A(new_n258), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT5), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n413), .B1(new_n259), .B2(new_n261), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(new_n252), .A3(G116), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(G113), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n412), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  OAI22_X1  g231(.A1(new_n411), .A2(new_n263), .B1(new_n379), .B2(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(G110), .B(G122), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n417), .ZN(new_n422));
  AOI22_X1  g236(.A1(new_n362), .A2(new_n264), .B1(new_n422), .B2(new_n351), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n419), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n421), .A2(KEYINPUT6), .A3(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n266), .A2(G125), .A3(new_n219), .ZN(new_n426));
  INV_X1    g240(.A(G125), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n268), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G224), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n430), .A2(G953), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n431), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n426), .A2(new_n428), .A3(new_n433), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  OR3_X1    g249(.A1(new_n423), .A2(KEYINPUT6), .A3(new_n419), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n425), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT7), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n433), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n432), .A2(new_n434), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n416), .B1(KEYINPUT5), .B2(new_n255), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n351), .B1(new_n258), .B2(new_n441), .ZN(new_n442));
  XOR2_X1   g256(.A(KEYINPUT83), .B(KEYINPUT8), .Z(new_n443));
  XNOR2_X1  g257(.A(new_n443), .B(new_n419), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n442), .B(new_n444), .C1(new_n351), .C2(new_n417), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n426), .A2(new_n428), .A3(new_n438), .A4(new_n433), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n440), .A2(new_n424), .A3(new_n445), .A4(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n316), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n409), .B1(new_n437), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n425), .A2(new_n435), .A3(new_n436), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n450), .A2(new_n316), .A3(new_n408), .A4(new_n447), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n407), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  XOR2_X1   g266(.A(KEYINPUT9), .B(G234), .Z(new_n453));
  XNOR2_X1  g267(.A(new_n453), .B(KEYINPUT77), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n316), .ZN(new_n455));
  AND2_X1   g269(.A1(new_n455), .A2(G221), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  AND3_X1   g271(.A1(new_n405), .A2(new_n452), .A3(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(G953), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n454), .A2(G217), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n251), .A2(G122), .ZN(new_n461));
  INV_X1    g275(.A(G122), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(G116), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  AND2_X1   g278(.A1(new_n464), .A2(new_n338), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT90), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n466), .B1(new_n461), .B2(KEYINPUT14), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT14), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n468), .A2(new_n251), .A3(KEYINPUT90), .A4(G122), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n461), .A2(KEYINPUT14), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n467), .A2(new_n463), .A3(new_n469), .A4(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n465), .B1(new_n471), .B2(G107), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n210), .A2(G128), .A3(new_n211), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT88), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n210), .A2(KEYINPUT88), .A3(G128), .A4(new_n211), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n209), .A2(G128), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n190), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  AOI211_X1 g294(.A(G134), .B(new_n478), .C1(new_n475), .C2(new_n476), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n472), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT91), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  OAI211_X1 g298(.A(KEYINPUT91), .B(new_n472), .C1(new_n480), .C2(new_n481), .ZN(new_n485));
  AND2_X1   g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT92), .ZN(new_n487));
  AOI21_X1  g301(.A(KEYINPUT13), .B1(new_n475), .B2(new_n476), .ZN(new_n488));
  OAI21_X1  g302(.A(KEYINPUT89), .B1(new_n488), .B2(new_n478), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT13), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n225), .A2(new_n226), .ZN(new_n491));
  AOI21_X1  g305(.A(KEYINPUT88), .B1(new_n491), .B2(G128), .ZN(new_n492));
  INV_X1    g306(.A(new_n476), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n490), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT89), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n494), .A2(new_n495), .A3(new_n479), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n475), .A2(KEYINPUT13), .A3(new_n476), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n489), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G134), .ZN(new_n499));
  INV_X1    g313(.A(new_n481), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n464), .B(new_n338), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n486), .A2(new_n487), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n484), .A2(new_n485), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n502), .B1(new_n498), .B2(G134), .ZN(new_n507));
  OAI21_X1  g321(.A(KEYINPUT92), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n460), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  NOR3_X1   g323(.A1(new_n506), .A2(new_n507), .A3(KEYINPUT92), .ZN(new_n510));
  INV_X1    g324(.A(new_n460), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n316), .B1(new_n509), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(G478), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n514), .A2(KEYINPUT15), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n515), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n316), .B(new_n517), .C1(new_n509), .C2(new_n512), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(G140), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(G125), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n427), .A2(G140), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n521), .A2(new_n522), .A3(KEYINPUT16), .ZN(new_n523));
  OR3_X1    g337(.A1(new_n427), .A2(KEYINPUT16), .A3(G140), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n523), .A2(new_n524), .A3(G146), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(G146), .B1(new_n523), .B2(new_n524), .ZN(new_n527));
  OAI21_X1  g341(.A(KEYINPUT86), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AND2_X1   g342(.A1(KEYINPUT71), .A2(G237), .ZN(new_n529));
  NOR2_X1   g343(.A1(KEYINPUT71), .A2(G237), .ZN(new_n530));
  OAI211_X1 g344(.A(G214), .B(new_n459), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n491), .ZN(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT71), .B(G237), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n533), .A2(G143), .A3(G214), .A4(new_n459), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n535), .A2(KEYINPUT17), .A3(G131), .ZN(new_n536));
  INV_X1    g350(.A(new_n527), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT86), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n537), .A2(new_n538), .A3(new_n525), .ZN(new_n539));
  AND3_X1   g353(.A1(new_n528), .A2(new_n536), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n535), .A2(G131), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT17), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n532), .A2(new_n534), .A3(new_n203), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n521), .A2(new_n522), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(KEYINPUT84), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(G146), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n521), .A2(new_n522), .A3(new_n220), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(KEYINPUT18), .A2(G131), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n550), .B1(new_n535), .B2(KEYINPUT85), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT85), .ZN(new_n552));
  INV_X1    g366(.A(new_n550), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n532), .A2(new_n534), .A3(new_n552), .A4(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  AOI22_X1  g369(.A1(new_n540), .A2(new_n544), .B1(new_n549), .B2(new_n555), .ZN(new_n556));
  XNOR2_X1  g370(.A(G113), .B(G122), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n557), .B(new_n340), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n544), .A2(new_n536), .A3(new_n528), .A4(new_n539), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n555), .A2(new_n549), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT87), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n560), .A2(new_n561), .A3(new_n562), .A4(new_n558), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n560), .A2(new_n558), .A3(new_n561), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(KEYINPUT87), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n559), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(G475), .B1(new_n566), .B2(G902), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT20), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n565), .A2(new_n563), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n545), .A2(KEYINPUT19), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n570), .B1(new_n546), .B2(KEYINPUT19), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n220), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n541), .A2(new_n543), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n572), .A2(new_n573), .A3(new_n525), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n558), .B1(new_n574), .B2(new_n561), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n569), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(G475), .A2(G902), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n568), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n575), .B1(new_n565), .B2(new_n563), .ZN(new_n580));
  INV_X1    g394(.A(new_n578), .ZN(new_n581));
  NOR3_X1   g395(.A1(new_n580), .A2(KEYINPUT20), .A3(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n567), .B1(new_n579), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(G234), .A2(G237), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n584), .A2(G952), .A3(new_n459), .ZN(new_n585));
  XOR2_X1   g399(.A(KEYINPUT21), .B(G898), .Z(new_n586));
  NAND3_X1  g400(.A1(new_n584), .A2(G902), .A3(G953), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  XOR2_X1   g402(.A(new_n588), .B(KEYINPUT93), .Z(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NOR3_X1   g404(.A1(new_n519), .A2(new_n583), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n252), .A2(G128), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n243), .A2(KEYINPUT23), .A3(G119), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n252), .A2(G128), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n592), .B(new_n593), .C1(new_n594), .C2(KEYINPUT23), .ZN(new_n595));
  XNOR2_X1  g409(.A(KEYINPUT24), .B(G110), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n243), .A2(G119), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n598), .A2(new_n592), .ZN(new_n599));
  AOI22_X1  g413(.A1(new_n595), .A2(G110), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n600), .B1(new_n526), .B2(new_n527), .ZN(new_n601));
  OAI22_X1  g415(.A1(new_n595), .A2(G110), .B1(new_n597), .B2(new_n599), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n602), .A2(new_n525), .A3(new_n548), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n459), .A2(G221), .A3(G234), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(KEYINPUT22), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(G137), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n604), .B(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n316), .ZN(new_n609));
  NOR2_X1   g423(.A1(KEYINPUT75), .A2(KEYINPUT25), .ZN(new_n610));
  OR2_X1    g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(KEYINPUT75), .A2(KEYINPUT25), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n609), .A2(new_n610), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(G217), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n615), .B1(G234), .B2(new_n316), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n616), .A2(G902), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(KEYINPUT76), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n608), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n328), .A2(new_n458), .A3(new_n591), .A4(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(G101), .ZN(G3));
  INV_X1    g438(.A(G472), .ZN(new_n625));
  OR2_X1    g439(.A1(new_n625), .A2(KEYINPUT94), .ZN(new_n626));
  AND3_X1   g440(.A1(new_n306), .A2(new_n316), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n626), .B1(new_n306), .B2(new_n316), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n627), .A2(new_n628), .A3(new_n621), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n405), .A2(new_n457), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n452), .A2(new_n589), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n514), .A2(G902), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n487), .B1(new_n486), .B2(new_n504), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n511), .B1(new_n635), .B2(new_n510), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT33), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n505), .A2(new_n460), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n486), .B(new_n504), .C1(KEYINPUT95), .C2(new_n511), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n511), .A2(KEYINPUT95), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n641), .B1(new_n506), .B2(new_n507), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n637), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n634), .B1(new_n639), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n636), .A2(new_n638), .ZN(new_n646));
  AOI21_X1  g460(.A(G478), .B1(new_n646), .B2(new_n316), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n583), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n632), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n631), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT34), .B(G104), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G6));
  INV_X1    g466(.A(new_n519), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n632), .A2(new_n653), .A3(new_n583), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n631), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT35), .B(G107), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G9));
  NOR2_X1   g471(.A1(new_n627), .A2(new_n628), .ZN(new_n658));
  INV_X1    g472(.A(new_n607), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n659), .A2(KEYINPUT36), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(new_n604), .ZN(new_n661));
  AOI22_X1  g475(.A1(new_n614), .A2(new_n616), .B1(new_n619), .B2(new_n661), .ZN(new_n662));
  NOR4_X1   g476(.A1(new_n519), .A2(new_n583), .A3(new_n662), .A4(new_n590), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n458), .A2(new_n658), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(KEYINPUT37), .B(G110), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT96), .B(KEYINPUT97), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G12));
  INV_X1    g482(.A(new_n662), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n452), .A2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n587), .A2(G900), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  OR2_X1    g487(.A1(new_n673), .A2(KEYINPUT98), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(KEYINPUT98), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n674), .A2(new_n585), .A3(new_n675), .ZN(new_n676));
  OAI211_X1 g490(.A(new_n567), .B(new_n676), .C1(new_n579), .C2(new_n582), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n653), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n328), .A2(new_n630), .A3(new_n671), .A4(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT99), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n677), .ZN(new_n682));
  AND4_X1   g496(.A1(new_n457), .A2(new_n405), .A3(new_n682), .A4(new_n519), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n683), .A2(KEYINPUT99), .A3(new_n328), .A4(new_n671), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G128), .ZN(G30));
  XNOR2_X1  g500(.A(new_n676), .B(KEYINPUT39), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n630), .A2(new_n687), .ZN(new_n688));
  XOR2_X1   g502(.A(new_n688), .B(KEYINPUT40), .Z(new_n689));
  AND3_X1   g503(.A1(new_n306), .A2(KEYINPUT32), .A3(new_n307), .ZN(new_n690));
  AOI21_X1  g504(.A(KEYINPUT32), .B1(new_n306), .B2(new_n307), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n313), .A2(new_n290), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n300), .A2(new_n290), .A3(new_n274), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n316), .ZN(new_n695));
  OAI21_X1  g509(.A(G472), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n449), .A2(new_n451), .ZN(new_n698));
  XOR2_X1   g512(.A(new_n698), .B(KEYINPUT38), .Z(new_n699));
  OR2_X1    g513(.A1(new_n566), .A2(G902), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n577), .A2(new_n568), .A3(new_n578), .ZN(new_n701));
  OAI21_X1  g515(.A(KEYINPUT20), .B1(new_n580), .B2(new_n581), .ZN(new_n702));
  AOI22_X1  g516(.A1(new_n700), .A2(G475), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NOR4_X1   g517(.A1(new_n699), .A2(new_n407), .A3(new_n653), .A4(new_n703), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n689), .A2(new_n662), .A3(new_n697), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(new_n239), .ZN(G45));
  NAND2_X1  g520(.A1(new_n405), .A2(new_n457), .ZN(new_n707));
  OAI211_X1 g521(.A(new_n583), .B(new_n676), .C1(new_n645), .C2(new_n647), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n709), .A2(new_n328), .A3(new_n671), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(new_n220), .ZN(G48));
  OAI21_X1  g525(.A(new_n316), .B1(new_n400), .B2(new_n401), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT100), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n713), .A2(new_n398), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  OAI221_X1 g529(.A(new_n316), .B1(new_n713), .B2(new_n398), .C1(new_n400), .C2(new_n401), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n717), .A2(new_n456), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n649), .A2(new_n328), .A3(new_n622), .A4(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(KEYINPUT101), .ZN(new_n720));
  XNOR2_X1  g534(.A(KEYINPUT41), .B(G113), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n720), .B(new_n721), .ZN(G15));
  NAND4_X1  g536(.A1(new_n654), .A2(new_n328), .A3(new_n622), .A4(new_n718), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G116), .ZN(G18));
  AND4_X1   g538(.A1(new_n452), .A2(new_n715), .A3(new_n457), .A4(new_n716), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n328), .A2(new_n725), .A3(new_n663), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G119), .ZN(G21));
  NAND2_X1  g541(.A1(new_n701), .A2(new_n702), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n407), .B1(new_n728), .B2(new_n567), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n729), .A2(new_n519), .A3(new_n698), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT103), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n729), .A2(new_n519), .A3(KEYINPUT103), .A4(new_n698), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n306), .A2(new_n316), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(G472), .ZN(new_n736));
  AOI22_X1  g550(.A1(new_n323), .A2(new_n290), .B1(new_n294), .B2(KEYINPUT31), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT102), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n292), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n323), .A2(new_n290), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n740), .A2(new_n738), .A3(new_n295), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n307), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n736), .A2(new_n622), .A3(new_n742), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n717), .A2(new_n456), .A3(new_n590), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n734), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G122), .ZN(G24));
  NAND2_X1  g560(.A1(new_n740), .A2(new_n295), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(KEYINPUT102), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n737), .A2(new_n738), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n748), .A2(new_n292), .A3(new_n749), .ZN(new_n750));
  AOI22_X1  g564(.A1(new_n307), .A2(new_n750), .B1(new_n735), .B2(G472), .ZN(new_n751));
  INV_X1    g565(.A(new_n708), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n725), .A2(new_n751), .A3(new_n752), .A4(new_n669), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(KEYINPUT104), .ZN(new_n754));
  AOI22_X1  g568(.A1(new_n319), .A2(KEYINPUT73), .B1(new_n298), .B2(new_n274), .ZN(new_n755));
  INV_X1    g569(.A(new_n304), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n291), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n297), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g573(.A(G902), .B1(new_n759), .B2(new_n296), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n742), .B(new_n669), .C1(new_n760), .C2(new_n625), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT104), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n762), .A2(new_n763), .A3(new_n752), .A4(new_n725), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n754), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G125), .ZN(G27));
  AOI21_X1  g580(.A(new_n621), .B1(new_n692), .B2(new_n326), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n698), .A2(new_n407), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n767), .A2(KEYINPUT42), .A3(new_n709), .A4(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT42), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n328), .A2(new_n622), .A3(new_n768), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n630), .A2(new_n752), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n769), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G131), .ZN(G33));
  NAND4_X1  g589(.A1(new_n683), .A2(new_n622), .A3(new_n328), .A4(new_n768), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G134), .ZN(G36));
  NOR3_X1   g591(.A1(new_n509), .A2(new_n512), .A3(KEYINPUT33), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n633), .B1(new_n778), .B2(new_n643), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n513), .A2(new_n514), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(new_n703), .ZN(new_n782));
  OR2_X1    g596(.A1(new_n782), .A2(KEYINPUT43), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n658), .A2(new_n662), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n782), .A2(KEYINPUT43), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n783), .A2(new_n784), .A3(KEYINPUT44), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n768), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT105), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT44), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n783), .A2(new_n785), .ZN(new_n791));
  INV_X1    g605(.A(new_n784), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n786), .A2(KEYINPUT105), .A3(new_n768), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n789), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(KEYINPUT106), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT106), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n789), .A2(new_n797), .A3(new_n793), .A4(new_n794), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n374), .B1(new_n396), .B2(new_n372), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT45), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n398), .B1(new_n799), .B2(new_n800), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n403), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n803), .A2(KEYINPUT46), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n402), .B1(new_n803), .B2(KEYINPUT46), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n457), .B(new_n687), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n796), .A2(new_n798), .A3(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(KEYINPUT107), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G137), .ZN(G39));
  OAI21_X1  g624(.A(new_n457), .B1(new_n804), .B2(new_n805), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n811), .A2(KEYINPUT47), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(KEYINPUT47), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n768), .A2(new_n621), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n328), .A2(new_n708), .A3(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n812), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(KEYINPUT108), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT108), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n812), .A2(new_n818), .A3(new_n813), .A4(new_n815), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(G140), .ZN(G42));
  XOR2_X1   g635(.A(KEYINPUT116), .B(KEYINPUT48), .Z(new_n822));
  NOR2_X1   g636(.A1(new_n791), .A2(new_n585), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n823), .A2(new_n718), .A3(new_n768), .ZN(new_n824));
  INV_X1    g638(.A(new_n767), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n822), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n824), .A2(new_n825), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n827), .A2(KEYINPUT116), .A3(KEYINPUT48), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n823), .A2(new_n743), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(new_n725), .ZN(new_n831));
  INV_X1    g645(.A(G952), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n718), .A2(new_n768), .ZN(new_n833));
  NOR4_X1   g647(.A1(new_n697), .A2(new_n833), .A3(new_n585), .A4(new_n621), .ZN(new_n834));
  INV_X1    g648(.A(new_n648), .ZN(new_n835));
  AOI211_X1 g649(.A(new_n832), .B(G953), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  AND4_X1   g650(.A1(new_n826), .A2(new_n828), .A3(new_n831), .A4(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT113), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n699), .A2(new_n407), .A3(new_n718), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n838), .B1(new_n829), .B2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT50), .ZN(new_n841));
  INV_X1    g655(.A(new_n839), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n823), .A2(KEYINPUT113), .A3(new_n743), .A4(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n840), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT114), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT114), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n840), .A2(new_n846), .A3(new_n841), .A4(new_n843), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n829), .A2(new_n839), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT50), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n845), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n717), .A2(new_n457), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n851), .B1(new_n812), .B2(new_n813), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n830), .A2(new_n768), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n834), .A2(new_n703), .A3(new_n780), .A4(new_n779), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n855), .B1(new_n824), .B2(new_n761), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n850), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT51), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n837), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT115), .ZN(new_n861));
  OAI221_X1 g675(.A(new_n855), .B1(new_n761), .B2(new_n824), .C1(new_n852), .C2(new_n853), .ZN(new_n862));
  AOI22_X1  g676(.A1(new_n844), .A2(KEYINPUT114), .B1(KEYINPUT50), .B2(new_n848), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n862), .B1(new_n863), .B2(new_n847), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n861), .B1(new_n864), .B2(KEYINPUT51), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n858), .A2(KEYINPUT115), .A3(new_n859), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n860), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT52), .ZN(new_n868));
  INV_X1    g682(.A(new_n710), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n670), .B1(new_n692), .B2(new_n326), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT99), .B1(new_n870), .B2(new_n683), .ZN(new_n871));
  INV_X1    g685(.A(new_n684), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n869), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n405), .A2(new_n457), .A3(new_n676), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n734), .A2(new_n697), .A3(new_n662), .A4(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n761), .A2(new_n708), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n763), .B1(new_n876), .B2(new_n725), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n452), .A2(new_n715), .A3(new_n457), .A4(new_n716), .ZN(new_n878));
  NOR4_X1   g692(.A1(new_n761), .A2(new_n878), .A3(KEYINPUT104), .A4(new_n708), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n875), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n868), .B1(new_n873), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n710), .B1(new_n681), .B2(new_n684), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n882), .A2(KEYINPUT52), .A3(new_n765), .A4(new_n875), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n881), .A2(KEYINPUT111), .A3(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT109), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n517), .B1(new_n646), .B2(new_n316), .ZN(new_n886));
  INV_X1    g700(.A(new_n518), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n516), .A2(KEYINPUT109), .A3(new_n518), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n677), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n328), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n751), .A2(new_n752), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n630), .A2(new_n669), .A3(new_n768), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(KEYINPUT110), .B1(new_n896), .B2(new_n776), .ZN(new_n897));
  AOI22_X1  g711(.A1(new_n328), .A2(new_n890), .B1(new_n751), .B2(new_n752), .ZN(new_n898));
  OAI211_X1 g712(.A(KEYINPUT110), .B(new_n776), .C1(new_n898), .C2(new_n894), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n888), .A2(new_n703), .A3(new_n889), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n648), .ZN(new_n903));
  INV_X1    g717(.A(new_n632), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n903), .A2(new_n630), .A3(new_n904), .A4(new_n629), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n745), .A2(new_n723), .A3(new_n905), .ZN(new_n906));
  AND4_X1   g720(.A1(new_n623), .A2(new_n719), .A3(new_n664), .A4(new_n726), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n906), .A2(new_n907), .A3(new_n774), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n901), .A2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT111), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n910), .B(new_n868), .C1(new_n873), .C2(new_n880), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n884), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT53), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n912), .A2(KEYINPUT112), .A3(new_n913), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n734), .A2(new_n662), .A3(new_n697), .ZN(new_n915));
  AOI22_X1  g729(.A1(new_n915), .A2(new_n874), .B1(new_n754), .B2(new_n764), .ZN(new_n916));
  AOI21_X1  g730(.A(KEYINPUT52), .B1(new_n916), .B2(new_n882), .ZN(new_n917));
  AND4_X1   g731(.A1(KEYINPUT52), .A2(new_n882), .A3(new_n765), .A4(new_n875), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n909), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n914), .B1(new_n913), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(KEYINPUT112), .B1(new_n912), .B2(new_n913), .ZN(new_n921));
  OAI21_X1  g735(.A(KEYINPUT54), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n918), .A2(new_n917), .ZN(new_n923));
  INV_X1    g737(.A(new_n908), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n896), .A2(new_n776), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT110), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n899), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n924), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n913), .B1(new_n923), .B2(new_n929), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n884), .A2(new_n909), .A3(KEYINPUT53), .A4(new_n911), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  OR2_X1    g746(.A1(new_n932), .A2(KEYINPUT54), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n867), .A2(new_n922), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n832), .A2(new_n459), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n621), .A2(new_n407), .A3(new_n456), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n699), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n717), .B(KEYINPUT49), .ZN(new_n939));
  OR4_X1    g753(.A1(new_n697), .A2(new_n938), .A3(new_n782), .A4(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n936), .A2(new_n940), .ZN(G75));
  AOI21_X1  g755(.A(new_n316), .B1(new_n930), .B2(new_n931), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(G210), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT56), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n425), .A2(new_n436), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(new_n435), .Z(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT55), .ZN(new_n948));
  OAI21_X1  g762(.A(KEYINPUT118), .B1(new_n945), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(KEYINPUT56), .B1(new_n942), .B2(G210), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT118), .ZN(new_n951));
  INV_X1    g765(.A(new_n948), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n949), .A2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT117), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n945), .A2(new_n955), .A3(new_n948), .ZN(new_n956));
  OAI21_X1  g770(.A(KEYINPUT117), .B1(new_n950), .B2(new_n952), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n459), .A2(G952), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n954), .A2(new_n958), .A3(new_n960), .ZN(G51));
  XNOR2_X1  g775(.A(new_n932), .B(KEYINPUT54), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n403), .B(KEYINPUT57), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n964), .B1(new_n401), .B2(new_n400), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n942), .A2(new_n801), .A3(new_n802), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(KEYINPUT119), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n959), .B1(new_n965), .B2(new_n967), .ZN(G54));
  NAND3_X1  g782(.A1(new_n942), .A2(KEYINPUT58), .A3(G475), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT120), .ZN(new_n970));
  AND3_X1   g784(.A1(new_n969), .A2(new_n970), .A3(new_n580), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n960), .B1(new_n969), .B2(new_n580), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n970), .B1(new_n969), .B2(new_n580), .ZN(new_n973));
  NOR3_X1   g787(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(G60));
  NOR2_X1   g788(.A1(new_n778), .A2(new_n643), .ZN(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n922), .A2(new_n933), .ZN(new_n977));
  NAND2_X1  g791(.A1(G478), .A2(G902), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT59), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n976), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n962), .A2(new_n976), .A3(new_n979), .ZN(new_n981));
  NOR3_X1   g795(.A1(new_n980), .A2(new_n959), .A3(new_n981), .ZN(G63));
  XNOR2_X1  g796(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT121), .ZN(new_n984));
  NAND2_X1  g798(.A1(G217), .A2(G902), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(KEYINPUT60), .ZN(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n984), .B1(new_n932), .B2(new_n987), .ZN(new_n988));
  AOI211_X1 g802(.A(KEYINPUT121), .B(new_n986), .C1(new_n930), .C2(new_n931), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n608), .B(KEYINPUT123), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n959), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n661), .B(KEYINPUT122), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n993), .B1(new_n988), .B2(new_n989), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n983), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n932), .A2(new_n987), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(KEYINPUT121), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n932), .A2(new_n984), .A3(new_n987), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n997), .A2(new_n998), .A3(new_n991), .ZN(new_n999));
  AND4_X1   g813(.A1(new_n960), .A2(new_n999), .A3(new_n983), .A4(new_n994), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n995), .A2(new_n1000), .ZN(G66));
  AND2_X1   g815(.A1(new_n906), .A2(new_n907), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n430), .A2(new_n459), .ZN(new_n1003));
  AOI22_X1  g817(.A1(new_n1002), .A2(new_n459), .B1(new_n586), .B2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n946), .B1(G898), .B2(new_n459), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1004), .B(new_n1005), .ZN(G69));
  AND2_X1   g820(.A1(new_n882), .A2(new_n765), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1007), .A2(new_n705), .ZN(new_n1008));
  INV_X1    g822(.A(KEYINPUT62), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n1007), .A2(new_n705), .A3(KEYINPUT62), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(new_n903), .ZN(new_n1013));
  NOR3_X1   g827(.A1(new_n1013), .A2(new_n771), .A3(new_n688), .ZN(new_n1014));
  INV_X1    g828(.A(new_n1014), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n1012), .A2(new_n808), .A3(new_n820), .A4(new_n1015), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(KEYINPUT125), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1014), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1018));
  INV_X1    g832(.A(KEYINPUT125), .ZN(new_n1019));
  NAND4_X1  g833(.A1(new_n1018), .A2(new_n1019), .A3(new_n808), .A4(new_n820), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n250), .A2(new_n271), .ZN(new_n1022));
  XNOR2_X1  g836(.A(new_n1022), .B(new_n571), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n1021), .A2(new_n459), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g838(.A(G900), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1025), .B1(new_n1023), .B2(new_n369), .ZN(new_n1026));
  AND2_X1   g840(.A1(new_n767), .A2(new_n734), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n807), .A2(new_n1027), .ZN(new_n1028));
  NAND4_X1  g842(.A1(new_n808), .A2(new_n820), .A3(new_n1007), .A4(new_n1028), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n774), .A2(new_n459), .A3(new_n776), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1031), .B1(G227), .B2(G953), .ZN(new_n1032));
  OAI221_X1 g846(.A(new_n1024), .B1(new_n459), .B2(new_n1026), .C1(new_n1032), .C2(new_n1023), .ZN(G72));
  NAND2_X1  g847(.A1(G472), .A2(G902), .ZN(new_n1034));
  XOR2_X1   g848(.A(new_n1034), .B(KEYINPUT63), .Z(new_n1035));
  NAND2_X1  g849(.A1(new_n924), .A2(new_n776), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1035), .B1(new_n1029), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g851(.A(new_n314), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n959), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g853(.A(new_n693), .ZN(new_n1040));
  NAND3_X1  g854(.A1(new_n1040), .A2(new_n314), .A3(new_n1035), .ZN(new_n1041));
  XOR2_X1   g855(.A(new_n1041), .B(KEYINPUT127), .Z(new_n1042));
  OAI21_X1  g856(.A(new_n1042), .B1(new_n920), .B2(new_n921), .ZN(new_n1043));
  NAND3_X1  g857(.A1(new_n1017), .A2(new_n1020), .A3(new_n1002), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n1040), .B1(new_n1044), .B2(new_n1035), .ZN(new_n1045));
  OAI211_X1 g859(.A(new_n1039), .B(new_n1043), .C1(new_n1045), .C2(KEYINPUT126), .ZN(new_n1046));
  AND2_X1   g860(.A1(new_n1045), .A2(KEYINPUT126), .ZN(new_n1047));
  NOR2_X1   g861(.A1(new_n1046), .A2(new_n1047), .ZN(G57));
endmodule


