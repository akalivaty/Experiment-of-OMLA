

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728;

  NOR2_X1 U368 ( .A1(n534), .A2(n470), .ZN(n471) );
  NOR2_X1 U369 ( .A1(n572), .A2(n571), .ZN(n641) );
  NOR2_X2 U370 ( .A1(n607), .A2(n714), .ZN(n608) );
  NOR2_X2 U371 ( .A1(n612), .A2(n714), .ZN(n614) );
  XNOR2_X1 U372 ( .A(n395), .B(n394), .ZN(n508) );
  XNOR2_X1 U373 ( .A(n375), .B(n593), .ZN(n598) );
  XNOR2_X1 U374 ( .A(n516), .B(n515), .ZN(n727) );
  NAND2_X1 U375 ( .A1(n390), .A2(n389), .ZN(n388) );
  NOR2_X1 U376 ( .A1(n509), .A2(n508), .ZN(n673) );
  XNOR2_X1 U377 ( .A(KEYINPUT93), .B(KEYINPUT15), .ZN(n409) );
  INV_X2 U378 ( .A(G953), .ZN(n718) );
  INV_X1 U379 ( .A(G143), .ZN(n404) );
  NOR2_X2 U380 ( .A1(n618), .A2(n714), .ZN(n619) );
  BUF_X1 U381 ( .A(n699), .Z(n710) );
  XNOR2_X2 U382 ( .A(n716), .B(G146), .ZN(n464) );
  NOR2_X1 U383 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U384 ( .A(n360), .B(n396), .ZN(n436) );
  XNOR2_X1 U385 ( .A(G122), .B(G116), .ZN(n360) );
  NAND2_X1 U386 ( .A1(n387), .A2(n551), .ZN(n570) );
  XNOR2_X1 U387 ( .A(n550), .B(n549), .ZN(n387) );
  INV_X1 U388 ( .A(KEYINPUT77), .ZN(n549) );
  XNOR2_X1 U389 ( .A(n521), .B(KEYINPUT106), .ZN(n661) );
  NOR2_X1 U390 ( .A1(n647), .A2(n644), .ZN(n521) );
  XNOR2_X1 U391 ( .A(n350), .B(n430), .ZN(n431) );
  XNOR2_X1 U392 ( .A(G131), .B(G143), .ZN(n427) );
  XNOR2_X1 U393 ( .A(n426), .B(n384), .ZN(n383) );
  INV_X1 U394 ( .A(G140), .ZN(n384) );
  XNOR2_X1 U395 ( .A(G113), .B(G104), .ZN(n426) );
  XNOR2_X1 U396 ( .A(n423), .B(n378), .ZN(n482) );
  INV_X1 U397 ( .A(KEYINPUT10), .ZN(n378) );
  NAND2_X1 U398 ( .A1(n587), .A2(n376), .ZN(n375) );
  AND2_X1 U399 ( .A1(n586), .A2(n355), .ZN(n376) );
  INV_X1 U400 ( .A(KEYINPUT108), .ZN(n391) );
  INV_X1 U401 ( .A(n531), .ZN(n389) );
  XNOR2_X1 U402 ( .A(n393), .B(n392), .ZN(n477) );
  INV_X1 U403 ( .A(KEYINPUT8), .ZN(n392) );
  NAND2_X1 U404 ( .A1(n718), .A2(G234), .ZN(n393) );
  XNOR2_X1 U405 ( .A(n437), .B(n436), .ZN(n358) );
  XNOR2_X1 U406 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n402) );
  XOR2_X1 U407 ( .A(KEYINPUT91), .B(KEYINPUT79), .Z(n403) );
  XNOR2_X1 U408 ( .A(KEYINPUT94), .B(KEYINPUT4), .ZN(n400) );
  XNOR2_X1 U409 ( .A(n379), .B(G125), .ZN(n423) );
  INV_X1 U410 ( .A(G146), .ZN(n379) );
  XNOR2_X1 U411 ( .A(n361), .B(n436), .ZN(n621) );
  XNOR2_X1 U412 ( .A(n398), .B(n458), .ZN(n361) );
  NOR2_X2 U413 ( .A1(n654), .A2(n600), .ZN(n699) );
  BUF_X1 U414 ( .A(n510), .Z(n502) );
  AND2_X1 U415 ( .A1(n663), .A2(n655), .ZN(n559) );
  XNOR2_X1 U416 ( .A(n554), .B(n553), .ZN(n595) );
  INV_X1 U417 ( .A(KEYINPUT39), .ZN(n553) );
  XNOR2_X1 U418 ( .A(n502), .B(KEYINPUT92), .ZN(n591) );
  NOR2_X1 U419 ( .A1(n570), .A2(n588), .ZN(n386) );
  XNOR2_X1 U420 ( .A(n416), .B(n415), .ZN(n574) );
  OR2_X1 U421 ( .A1(n712), .A2(G902), .ZN(n395) );
  XNOR2_X1 U422 ( .A(n485), .B(n351), .ZN(n394) );
  XNOR2_X1 U423 ( .A(n354), .B(n433), .ZN(n520) );
  XNOR2_X1 U424 ( .A(n432), .B(G475), .ZN(n433) );
  NAND2_X1 U425 ( .A1(n368), .A2(n366), .ZN(n534) );
  AND2_X1 U426 ( .A1(n370), .A2(n369), .ZN(n368) );
  NAND2_X1 U427 ( .A1(n367), .A2(n371), .ZN(n366) );
  XNOR2_X1 U428 ( .A(n377), .B(n464), .ZN(n701) );
  XNOR2_X1 U429 ( .A(n453), .B(n359), .ZN(n377) );
  XNOR2_X1 U430 ( .A(n396), .B(G101), .ZN(n359) );
  AND2_X1 U431 ( .A1(n606), .A2(G953), .ZN(n714) );
  NOR2_X1 U432 ( .A1(G237), .A2(G953), .ZN(n429) );
  NOR2_X1 U433 ( .A1(n548), .A2(n547), .ZN(n550) );
  XNOR2_X1 U434 ( .A(n454), .B(G469), .ZN(n525) );
  NOR2_X1 U435 ( .A1(n701), .A2(G902), .ZN(n454) );
  XNOR2_X1 U436 ( .A(n449), .B(n448), .ZN(n716) );
  AND2_X1 U437 ( .A1(n520), .A2(n518), .ZN(n655) );
  XOR2_X1 U438 ( .A(n544), .B(n569), .Z(n657) );
  AND2_X1 U439 ( .A1(n347), .A2(n447), .ZN(n371) );
  XNOR2_X1 U440 ( .A(n382), .B(n425), .ZN(n609) );
  XNOR2_X1 U441 ( .A(n431), .B(n383), .ZN(n382) );
  XNOR2_X1 U442 ( .A(KEYINPUT12), .B(KEYINPUT102), .ZN(n424) );
  XNOR2_X1 U443 ( .A(n522), .B(n391), .ZN(n390) );
  BUF_X1 U444 ( .A(n500), .Z(n569) );
  OR2_X1 U445 ( .A1(n574), .A2(n353), .ZN(n364) );
  AND2_X1 U446 ( .A1(n373), .A2(n372), .ZN(n365) );
  XNOR2_X1 U447 ( .A(n483), .B(n715), .ZN(n712) );
  XNOR2_X1 U448 ( .A(n476), .B(n475), .ZN(n479) );
  XNOR2_X1 U449 ( .A(n438), .B(n358), .ZN(n440) );
  XNOR2_X1 U450 ( .A(n621), .B(n408), .ZN(n603) );
  XNOR2_X1 U451 ( .A(n565), .B(n357), .ZN(n726) );
  INV_X1 U452 ( .A(KEYINPUT42), .ZN(n357) );
  NOR2_X1 U453 ( .A1(n595), .A2(n555), .ZN(n557) );
  INV_X1 U454 ( .A(KEYINPUT32), .ZN(n504) );
  INV_X1 U455 ( .A(KEYINPUT112), .ZN(n385) );
  XNOR2_X1 U456 ( .A(n490), .B(KEYINPUT105), .ZN(n644) );
  XNOR2_X1 U457 ( .A(n703), .B(n702), .ZN(n704) );
  XNOR2_X1 U458 ( .A(n701), .B(n700), .ZN(n702) );
  AND2_X1 U459 ( .A1(n655), .A2(n669), .ZN(n347) );
  XOR2_X1 U460 ( .A(KEYINPUT67), .B(KEYINPUT0), .Z(n348) );
  NOR2_X1 U461 ( .A1(n534), .A2(n533), .ZN(n349) );
  XNOR2_X1 U462 ( .A(n434), .B(G134), .ZN(n449) );
  XOR2_X1 U463 ( .A(n428), .B(n427), .Z(n350) );
  NAND2_X2 U464 ( .A1(n365), .A2(n364), .ZN(n528) );
  XOR2_X1 U465 ( .A(n487), .B(n486), .Z(n351) );
  XOR2_X1 U466 ( .A(KEYINPUT97), .B(KEYINPUT23), .Z(n352) );
  OR2_X1 U467 ( .A1(n422), .A2(n348), .ZN(n353) );
  NOR2_X1 U468 ( .A1(n609), .A2(G902), .ZN(n354) );
  AND2_X1 U469 ( .A1(n651), .A2(n585), .ZN(n355) );
  INV_X1 U470 ( .A(G107), .ZN(n396) );
  XOR2_X1 U471 ( .A(KEYINPUT33), .B(KEYINPUT109), .Z(n356) );
  INV_X1 U472 ( .A(n447), .ZN(n374) );
  NAND2_X1 U473 ( .A1(n726), .A2(n725), .ZN(n567) );
  OR2_X1 U474 ( .A1(n347), .A2(n447), .ZN(n369) );
  XNOR2_X2 U475 ( .A(n363), .B(n362), .ZN(n458) );
  XNOR2_X2 U476 ( .A(KEYINPUT3), .B(G119), .ZN(n362) );
  XNOR2_X2 U477 ( .A(G113), .B(G101), .ZN(n363) );
  INV_X1 U478 ( .A(n528), .ZN(n367) );
  NAND2_X1 U479 ( .A1(n528), .A2(n374), .ZN(n370) );
  NAND2_X1 U480 ( .A1(n422), .A2(n348), .ZN(n372) );
  NAND2_X1 U481 ( .A1(n574), .A2(n348), .ZN(n373) );
  NOR2_X1 U482 ( .A1(n534), .A2(n380), .ZN(n505) );
  NAND2_X1 U483 ( .A1(n591), .A2(n381), .ZN(n380) );
  AND2_X1 U484 ( .A1(n531), .A2(n503), .ZN(n381) );
  XNOR2_X1 U485 ( .A(n386), .B(n385), .ZN(n571) );
  NAND2_X1 U486 ( .A1(n691), .A2(n367), .ZN(n512) );
  XNOR2_X2 U487 ( .A(n388), .B(n356), .ZN(n691) );
  XNOR2_X2 U488 ( .A(n469), .B(n468), .ZN(n672) );
  XNOR2_X1 U489 ( .A(KEYINPUT46), .B(KEYINPUT87), .ZN(n566) );
  XNOR2_X1 U490 ( .A(n482), .B(n424), .ZN(n425) );
  INV_X1 U491 ( .A(KEYINPUT24), .ZN(n473) );
  XNOR2_X1 U492 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U493 ( .A(n525), .B(n455), .ZN(n510) );
  INV_X1 U494 ( .A(KEYINPUT34), .ZN(n511) );
  XNOR2_X1 U495 ( .A(n706), .B(n705), .ZN(n707) );
  XNOR2_X1 U496 ( .A(n708), .B(n707), .ZN(n709) );
  XNOR2_X2 U497 ( .A(G110), .B(G104), .ZN(n451) );
  XNOR2_X1 U498 ( .A(KEYINPUT73), .B(KEYINPUT16), .ZN(n397) );
  XNOR2_X1 U499 ( .A(n451), .B(n397), .ZN(n398) );
  NAND2_X1 U500 ( .A1(n718), .A2(G224), .ZN(n399) );
  XNOR2_X1 U501 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U502 ( .A(n423), .B(n401), .ZN(n407) );
  XNOR2_X1 U503 ( .A(n403), .B(n402), .ZN(n405) );
  XNOR2_X2 U504 ( .A(n404), .B(G128), .ZN(n434) );
  XNOR2_X1 U505 ( .A(n405), .B(n434), .ZN(n406) );
  XNOR2_X1 U506 ( .A(n407), .B(n406), .ZN(n408) );
  INV_X1 U507 ( .A(G902), .ZN(n465) );
  XNOR2_X1 U508 ( .A(n409), .B(n465), .ZN(n600) );
  NAND2_X1 U509 ( .A1(n603), .A2(n600), .ZN(n413) );
  INV_X1 U510 ( .A(G237), .ZN(n410) );
  NAND2_X1 U511 ( .A1(n465), .A2(n410), .ZN(n414) );
  NAND2_X1 U512 ( .A1(n414), .A2(G210), .ZN(n411) );
  XNOR2_X1 U513 ( .A(n411), .B(KEYINPUT95), .ZN(n412) );
  XNOR2_X2 U514 ( .A(n413), .B(n412), .ZN(n500) );
  NAND2_X1 U515 ( .A1(n414), .A2(G214), .ZN(n656) );
  NAND2_X1 U516 ( .A1(n500), .A2(n656), .ZN(n416) );
  INV_X1 U517 ( .A(KEYINPUT19), .ZN(n415) );
  NAND2_X1 U518 ( .A1(G234), .A2(G237), .ZN(n417) );
  XNOR2_X1 U519 ( .A(KEYINPUT14), .B(n417), .ZN(n419) );
  NAND2_X1 U520 ( .A1(n419), .A2(G952), .ZN(n418) );
  XNOR2_X1 U521 ( .A(n418), .B(KEYINPUT96), .ZN(n688) );
  NOR2_X1 U522 ( .A1(n688), .A2(G953), .ZN(n493) );
  AND2_X1 U523 ( .A1(G953), .A2(n419), .ZN(n420) );
  NAND2_X1 U524 ( .A1(G902), .A2(n420), .ZN(n491) );
  NOR2_X1 U525 ( .A1(n491), .A2(G898), .ZN(n421) );
  NOR2_X1 U526 ( .A1(n493), .A2(n421), .ZN(n422) );
  XOR2_X1 U527 ( .A(KEYINPUT11), .B(G122), .Z(n428) );
  XNOR2_X1 U528 ( .A(n429), .B(KEYINPUT76), .ZN(n456) );
  NAND2_X1 U529 ( .A1(G214), .A2(n456), .ZN(n430) );
  XNOR2_X1 U530 ( .A(KEYINPUT13), .B(KEYINPUT103), .ZN(n432) );
  INV_X1 U531 ( .A(n449), .ZN(n438) );
  XOR2_X1 U532 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n435) );
  XNOR2_X1 U533 ( .A(n435), .B(KEYINPUT104), .ZN(n437) );
  NAND2_X1 U534 ( .A1(G217), .A2(n477), .ZN(n439) );
  XNOR2_X1 U535 ( .A(n440), .B(n439), .ZN(n706) );
  NOR2_X1 U536 ( .A1(G902), .A2(n706), .ZN(n441) );
  XNOR2_X1 U537 ( .A(n441), .B(G478), .ZN(n518) );
  NAND2_X1 U538 ( .A1(G234), .A2(n600), .ZN(n442) );
  XNOR2_X1 U539 ( .A(KEYINPUT20), .B(n442), .ZN(n484) );
  AND2_X1 U540 ( .A1(n484), .A2(G221), .ZN(n445) );
  INV_X1 U541 ( .A(KEYINPUT99), .ZN(n443) );
  XNOR2_X1 U542 ( .A(n443), .B(KEYINPUT21), .ZN(n444) );
  XNOR2_X1 U543 ( .A(n445), .B(n444), .ZN(n669) );
  INV_X1 U544 ( .A(n669), .ZN(n509) );
  XNOR2_X1 U545 ( .A(KEYINPUT72), .B(KEYINPUT22), .ZN(n446) );
  XNOR2_X1 U546 ( .A(n446), .B(KEYINPUT71), .ZN(n447) );
  XNOR2_X1 U547 ( .A(KEYINPUT4), .B(G131), .ZN(n448) );
  XOR2_X1 U548 ( .A(G137), .B(G140), .Z(n480) );
  NAND2_X1 U549 ( .A1(G227), .A2(n718), .ZN(n450) );
  XNOR2_X1 U550 ( .A(n450), .B(n451), .ZN(n452) );
  XNOR2_X1 U551 ( .A(n480), .B(n452), .ZN(n453) );
  XNOR2_X1 U552 ( .A(KEYINPUT65), .B(KEYINPUT1), .ZN(n455) );
  INV_X1 U553 ( .A(n502), .ZN(n530) );
  NAND2_X1 U554 ( .A1(G210), .A2(n456), .ZN(n457) );
  XNOR2_X1 U555 ( .A(n458), .B(n457), .ZN(n462) );
  XOR2_X1 U556 ( .A(KEYINPUT75), .B(KEYINPUT5), .Z(n460) );
  XNOR2_X1 U557 ( .A(G116), .B(G137), .ZN(n459) );
  XNOR2_X1 U558 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U559 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U560 ( .A(n464), .B(n463), .ZN(n615) );
  NAND2_X1 U561 ( .A1(n615), .A2(n465), .ZN(n469) );
  XNOR2_X1 U562 ( .A(G472), .B(KEYINPUT100), .ZN(n467) );
  INV_X1 U563 ( .A(KEYINPUT70), .ZN(n466) );
  XNOR2_X1 U564 ( .A(n467), .B(n466), .ZN(n468) );
  NAND2_X1 U565 ( .A1(n530), .A2(n672), .ZN(n470) );
  XNOR2_X1 U566 ( .A(n471), .B(KEYINPUT64), .ZN(n488) );
  XNOR2_X1 U567 ( .A(G128), .B(KEYINPUT69), .ZN(n472) );
  XNOR2_X1 U568 ( .A(n352), .B(n472), .ZN(n476) );
  XNOR2_X1 U569 ( .A(G119), .B(G110), .ZN(n474) );
  NAND2_X1 U570 ( .A1(n477), .A2(G221), .ZN(n478) );
  XNOR2_X1 U571 ( .A(n479), .B(n478), .ZN(n483) );
  INV_X1 U572 ( .A(n480), .ZN(n481) );
  XNOR2_X1 U573 ( .A(n482), .B(n481), .ZN(n715) );
  NAND2_X1 U574 ( .A1(n484), .A2(G217), .ZN(n485) );
  XNOR2_X1 U575 ( .A(KEYINPUT98), .B(KEYINPUT25), .ZN(n487) );
  INV_X1 U576 ( .A(KEYINPUT78), .ZN(n486) );
  NAND2_X1 U577 ( .A1(n488), .A2(n508), .ZN(n506) );
  XNOR2_X1 U578 ( .A(n506), .B(G110), .ZN(G12) );
  INV_X1 U579 ( .A(n520), .ZN(n489) );
  NAND2_X1 U580 ( .A1(n518), .A2(n489), .ZN(n490) );
  INV_X1 U581 ( .A(n644), .ZN(n555) );
  NOR2_X1 U582 ( .A1(G900), .A2(n491), .ZN(n492) );
  NOR2_X1 U583 ( .A1(n493), .A2(n492), .ZN(n547) );
  NOR2_X1 U584 ( .A1(n509), .A2(n547), .ZN(n494) );
  NAND2_X1 U585 ( .A1(n508), .A2(n494), .ZN(n561) );
  INV_X1 U586 ( .A(KEYINPUT6), .ZN(n495) );
  XNOR2_X1 U587 ( .A(n672), .B(n495), .ZN(n531) );
  NOR2_X1 U588 ( .A1(n561), .A2(n531), .ZN(n496) );
  XNOR2_X1 U589 ( .A(n496), .B(KEYINPUT111), .ZN(n497) );
  NOR2_X1 U590 ( .A1(n555), .A2(n497), .ZN(n498) );
  NAND2_X1 U591 ( .A1(n498), .A2(n656), .ZN(n589) );
  NOR2_X1 U592 ( .A1(n502), .A2(n589), .ZN(n499) );
  XNOR2_X1 U593 ( .A(n499), .B(KEYINPUT43), .ZN(n501) );
  NOR2_X1 U594 ( .A1(n501), .A2(n569), .ZN(n596) );
  XOR2_X1 U595 ( .A(G140), .B(n596), .Z(G42) );
  XNOR2_X1 U596 ( .A(n508), .B(KEYINPUT107), .ZN(n668) );
  INV_X1 U597 ( .A(n668), .ZN(n503) );
  XNOR2_X1 U598 ( .A(n505), .B(n504), .ZN(n728) );
  NAND2_X1 U599 ( .A1(n506), .A2(n728), .ZN(n507) );
  XNOR2_X1 U600 ( .A(n507), .B(KEYINPUT89), .ZN(n517) );
  NAND2_X1 U601 ( .A1(n673), .A2(n510), .ZN(n522) );
  XNOR2_X1 U602 ( .A(n512), .B(n511), .ZN(n514) );
  NOR2_X1 U603 ( .A1(n518), .A2(n520), .ZN(n513) );
  XNOR2_X1 U604 ( .A(n513), .B(KEYINPUT110), .ZN(n568) );
  NAND2_X1 U605 ( .A1(n514), .A2(n568), .ZN(n516) );
  XOR2_X1 U606 ( .A(KEYINPUT80), .B(KEYINPUT35), .Z(n515) );
  NAND2_X1 U607 ( .A1(n517), .A2(n727), .ZN(n539) );
  NAND2_X1 U608 ( .A1(n539), .A2(KEYINPUT44), .ZN(n537) );
  INV_X1 U609 ( .A(n518), .ZN(n519) );
  AND2_X1 U610 ( .A1(n520), .A2(n519), .ZN(n647) );
  XNOR2_X1 U611 ( .A(KEYINPUT84), .B(n661), .ZN(n583) );
  NOR2_X1 U612 ( .A1(n672), .A2(n522), .ZN(n523) );
  XOR2_X1 U613 ( .A(KEYINPUT101), .B(n523), .Z(n679) );
  NAND2_X1 U614 ( .A1(n679), .A2(n367), .ZN(n524) );
  XNOR2_X1 U615 ( .A(n524), .B(KEYINPUT31), .ZN(n648) );
  INV_X1 U616 ( .A(n525), .ZN(n563) );
  NAND2_X1 U617 ( .A1(n563), .A2(n673), .ZN(n548) );
  INV_X1 U618 ( .A(n548), .ZN(n526) );
  NAND2_X1 U619 ( .A1(n526), .A2(n672), .ZN(n527) );
  NOR2_X1 U620 ( .A1(n528), .A2(n527), .ZN(n633) );
  NOR2_X1 U621 ( .A1(n648), .A2(n633), .ZN(n529) );
  NOR2_X1 U622 ( .A1(n583), .A2(n529), .ZN(n535) );
  AND2_X1 U623 ( .A1(n530), .A2(n668), .ZN(n532) );
  NAND2_X1 U624 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X1 U625 ( .A1(n535), .A2(n349), .ZN(n536) );
  NAND2_X1 U626 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U627 ( .A(n538), .B(KEYINPUT88), .ZN(n541) );
  NOR2_X1 U628 ( .A1(n539), .A2(KEYINPUT44), .ZN(n540) );
  NOR2_X2 U629 ( .A1(n541), .A2(n540), .ZN(n543) );
  XNOR2_X1 U630 ( .A(KEYINPUT86), .B(KEYINPUT45), .ZN(n542) );
  XNOR2_X1 U631 ( .A(n543), .B(n542), .ZN(n624) );
  XNOR2_X1 U632 ( .A(KEYINPUT38), .B(KEYINPUT74), .ZN(n544) );
  INV_X1 U633 ( .A(n672), .ZN(n545) );
  NAND2_X1 U634 ( .A1(n545), .A2(n656), .ZN(n546) );
  XOR2_X1 U635 ( .A(KEYINPUT30), .B(n546), .Z(n551) );
  INV_X1 U636 ( .A(n570), .ZN(n552) );
  NAND2_X1 U637 ( .A1(n657), .A2(n552), .ZN(n554) );
  INV_X1 U638 ( .A(KEYINPUT40), .ZN(n556) );
  XNOR2_X1 U639 ( .A(n557), .B(n556), .ZN(n725) );
  XNOR2_X1 U640 ( .A(KEYINPUT114), .B(KEYINPUT41), .ZN(n560) );
  NAND2_X1 U641 ( .A1(n657), .A2(n656), .ZN(n558) );
  XNOR2_X1 U642 ( .A(n558), .B(KEYINPUT113), .ZN(n663) );
  XNOR2_X1 U643 ( .A(n560), .B(n559), .ZN(n681) );
  NOR2_X1 U644 ( .A1(n672), .A2(n561), .ZN(n562) );
  XNOR2_X1 U645 ( .A(KEYINPUT28), .B(n562), .ZN(n564) );
  NAND2_X1 U646 ( .A1(n564), .A2(n563), .ZN(n575) );
  NOR2_X1 U647 ( .A1(n681), .A2(n575), .ZN(n565) );
  XNOR2_X1 U648 ( .A(n567), .B(n566), .ZN(n587) );
  INV_X1 U649 ( .A(n568), .ZN(n572) );
  INV_X1 U650 ( .A(n569), .ZN(n588) );
  XNOR2_X1 U651 ( .A(n641), .B(KEYINPUT85), .ZN(n581) );
  NAND2_X1 U652 ( .A1(n661), .A2(KEYINPUT47), .ZN(n573) );
  XNOR2_X1 U653 ( .A(n573), .B(KEYINPUT83), .ZN(n579) );
  NOR2_X1 U654 ( .A1(n575), .A2(n574), .ZN(n642) );
  INV_X1 U655 ( .A(n642), .ZN(n576) );
  NAND2_X1 U656 ( .A1(n576), .A2(KEYINPUT47), .ZN(n577) );
  XOR2_X1 U657 ( .A(KEYINPUT82), .B(n577), .Z(n578) );
  NAND2_X1 U658 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U659 ( .A(n582), .B(KEYINPUT81), .ZN(n586) );
  NOR2_X1 U660 ( .A1(KEYINPUT47), .A2(n583), .ZN(n584) );
  NAND2_X1 U661 ( .A1(n642), .A2(n584), .ZN(n585) );
  NOR2_X1 U662 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U663 ( .A(n590), .B(KEYINPUT36), .ZN(n592) );
  NAND2_X1 U664 ( .A1(n592), .A2(n591), .ZN(n651) );
  XOR2_X1 U665 ( .A(KEYINPUT48), .B(KEYINPUT68), .Z(n593) );
  INV_X1 U666 ( .A(n647), .ZN(n594) );
  NOR2_X1 U667 ( .A1(n595), .A2(n594), .ZN(n653) );
  NOR2_X1 U668 ( .A1(n596), .A2(n653), .ZN(n597) );
  NAND2_X1 U669 ( .A1(n598), .A2(n597), .ZN(n717) );
  NOR2_X1 U670 ( .A1(n624), .A2(n717), .ZN(n599) );
  XNOR2_X1 U671 ( .A(n599), .B(KEYINPUT2), .ZN(n654) );
  NAND2_X1 U672 ( .A1(n699), .A2(G210), .ZN(n605) );
  XNOR2_X1 U673 ( .A(KEYINPUT90), .B(KEYINPUT54), .ZN(n601) );
  XNOR2_X1 U674 ( .A(n601), .B(KEYINPUT55), .ZN(n602) );
  XNOR2_X1 U675 ( .A(n603), .B(n602), .ZN(n604) );
  XNOR2_X1 U676 ( .A(n605), .B(n604), .ZN(n607) );
  INV_X1 U677 ( .A(G952), .ZN(n606) );
  XNOR2_X1 U678 ( .A(n608), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U679 ( .A1(n699), .A2(G475), .ZN(n611) );
  XOR2_X1 U680 ( .A(n609), .B(KEYINPUT59), .Z(n610) );
  XNOR2_X1 U681 ( .A(n611), .B(n610), .ZN(n612) );
  XNOR2_X1 U682 ( .A(KEYINPUT66), .B(KEYINPUT60), .ZN(n613) );
  XNOR2_X1 U683 ( .A(n614), .B(n613), .ZN(G60) );
  INV_X1 U684 ( .A(KEYINPUT63), .ZN(n620) );
  NAND2_X1 U685 ( .A1(n699), .A2(G472), .ZN(n617) );
  XOR2_X1 U686 ( .A(KEYINPUT62), .B(n615), .Z(n616) );
  XNOR2_X1 U687 ( .A(n617), .B(n616), .ZN(n618) );
  XNOR2_X1 U688 ( .A(n620), .B(n619), .ZN(G57) );
  INV_X1 U689 ( .A(n621), .ZN(n623) );
  OR2_X1 U690 ( .A1(n718), .A2(G898), .ZN(n622) );
  NAND2_X1 U691 ( .A1(n623), .A2(n622), .ZN(n631) );
  NOR2_X1 U692 ( .A1(n624), .A2(G953), .ZN(n625) );
  XNOR2_X1 U693 ( .A(n625), .B(KEYINPUT127), .ZN(n629) );
  NAND2_X1 U694 ( .A1(G953), .A2(G224), .ZN(n626) );
  XNOR2_X1 U695 ( .A(KEYINPUT61), .B(n626), .ZN(n627) );
  NAND2_X1 U696 ( .A1(n627), .A2(G898), .ZN(n628) );
  NAND2_X1 U697 ( .A1(n629), .A2(n628), .ZN(n630) );
  XOR2_X1 U698 ( .A(n631), .B(n630), .Z(G69) );
  XOR2_X1 U699 ( .A(G101), .B(n349), .Z(G3) );
  NAND2_X1 U700 ( .A1(n633), .A2(n644), .ZN(n632) );
  XNOR2_X1 U701 ( .A(n632), .B(G104), .ZN(G6) );
  XOR2_X1 U702 ( .A(KEYINPUT115), .B(KEYINPUT27), .Z(n635) );
  NAND2_X1 U703 ( .A1(n633), .A2(n647), .ZN(n634) );
  XNOR2_X1 U704 ( .A(n635), .B(n634), .ZN(n637) );
  XOR2_X1 U705 ( .A(G107), .B(KEYINPUT26), .Z(n636) );
  XNOR2_X1 U706 ( .A(n637), .B(n636), .ZN(G9) );
  XOR2_X1 U707 ( .A(KEYINPUT116), .B(KEYINPUT29), .Z(n639) );
  NAND2_X1 U708 ( .A1(n642), .A2(n647), .ZN(n638) );
  XNOR2_X1 U709 ( .A(n639), .B(n638), .ZN(n640) );
  XNOR2_X1 U710 ( .A(G128), .B(n640), .ZN(G30) );
  XOR2_X1 U711 ( .A(G143), .B(n641), .Z(G45) );
  NAND2_X1 U712 ( .A1(n644), .A2(n642), .ZN(n643) );
  XNOR2_X1 U713 ( .A(n643), .B(G146), .ZN(G48) );
  XOR2_X1 U714 ( .A(G113), .B(KEYINPUT117), .Z(n646) );
  NAND2_X1 U715 ( .A1(n648), .A2(n644), .ZN(n645) );
  XNOR2_X1 U716 ( .A(n646), .B(n645), .ZN(G15) );
  NAND2_X1 U717 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U718 ( .A(n649), .B(G116), .ZN(G18) );
  XOR2_X1 U719 ( .A(KEYINPUT37), .B(KEYINPUT118), .Z(n650) );
  XNOR2_X1 U720 ( .A(n651), .B(n650), .ZN(n652) );
  XNOR2_X1 U721 ( .A(G125), .B(n652), .ZN(G27) );
  XOR2_X1 U722 ( .A(G134), .B(n653), .Z(G36) );
  INV_X1 U723 ( .A(n654), .ZN(n697) );
  INV_X1 U724 ( .A(n655), .ZN(n659) );
  NOR2_X1 U725 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U726 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U727 ( .A(KEYINPUT120), .B(n660), .Z(n665) );
  INV_X1 U728 ( .A(n661), .ZN(n662) );
  NAND2_X1 U729 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U730 ( .A1(n665), .A2(n664), .ZN(n666) );
  XOR2_X1 U731 ( .A(KEYINPUT121), .B(n666), .Z(n667) );
  NAND2_X1 U732 ( .A1(n667), .A2(n691), .ZN(n684) );
  NOR2_X1 U733 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U734 ( .A(n670), .B(KEYINPUT49), .ZN(n671) );
  NAND2_X1 U735 ( .A1(n672), .A2(n671), .ZN(n676) );
  NOR2_X1 U736 ( .A1(n673), .A2(n502), .ZN(n674) );
  XNOR2_X1 U737 ( .A(n674), .B(KEYINPUT50), .ZN(n675) );
  NOR2_X1 U738 ( .A1(n676), .A2(n675), .ZN(n677) );
  XOR2_X1 U739 ( .A(KEYINPUT119), .B(n677), .Z(n678) );
  NOR2_X1 U740 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U741 ( .A(n680), .B(KEYINPUT51), .ZN(n682) );
  INV_X1 U742 ( .A(n681), .ZN(n690) );
  NAND2_X1 U743 ( .A1(n682), .A2(n690), .ZN(n683) );
  NAND2_X1 U744 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U745 ( .A(n685), .B(KEYINPUT122), .ZN(n686) );
  XOR2_X1 U746 ( .A(KEYINPUT52), .B(n686), .Z(n687) );
  NOR2_X1 U747 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U748 ( .A(KEYINPUT123), .B(n689), .Z(n694) );
  NAND2_X1 U749 ( .A1(n691), .A2(n690), .ZN(n692) );
  XOR2_X1 U750 ( .A(KEYINPUT124), .B(n692), .Z(n693) );
  NOR2_X1 U751 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U752 ( .A1(n695), .A2(n718), .ZN(n696) );
  NOR2_X1 U753 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U754 ( .A(n698), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U755 ( .A1(n710), .A2(G469), .ZN(n703) );
  XOR2_X1 U756 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n700) );
  NOR2_X1 U757 ( .A1(n714), .A2(n704), .ZN(G54) );
  NAND2_X1 U758 ( .A1(n710), .A2(G478), .ZN(n708) );
  XOR2_X1 U759 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n705) );
  NOR2_X1 U760 ( .A1(n714), .A2(n709), .ZN(G63) );
  NAND2_X1 U761 ( .A1(n710), .A2(G217), .ZN(n711) );
  XNOR2_X1 U762 ( .A(n712), .B(n711), .ZN(n713) );
  NOR2_X1 U763 ( .A1(n714), .A2(n713), .ZN(G66) );
  XNOR2_X1 U764 ( .A(n716), .B(n715), .ZN(n720) );
  XNOR2_X1 U765 ( .A(n717), .B(n720), .ZN(n719) );
  NAND2_X1 U766 ( .A1(n719), .A2(n718), .ZN(n724) );
  XNOR2_X1 U767 ( .A(G227), .B(n720), .ZN(n721) );
  NAND2_X1 U768 ( .A1(n721), .A2(G900), .ZN(n722) );
  NAND2_X1 U769 ( .A1(n722), .A2(G953), .ZN(n723) );
  NAND2_X1 U770 ( .A1(n724), .A2(n723), .ZN(G72) );
  XNOR2_X1 U771 ( .A(G131), .B(n725), .ZN(G33) );
  XNOR2_X1 U772 ( .A(G137), .B(n726), .ZN(G39) );
  XNOR2_X1 U773 ( .A(n727), .B(G122), .ZN(G24) );
  XNOR2_X1 U774 ( .A(G119), .B(n728), .ZN(G21) );
endmodule

