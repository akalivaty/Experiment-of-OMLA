//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 0 0 1 0 1 1 0 0 0 0 0 1 0 0 1 1 1 0 1 1 0 0 0 1 0 1 1 0 0 1 1 1 0 0 1 1 1 1 0 0 1 0 0 1 1 0 1 1 0 1 1 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:57 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1237,
    new_n1238, new_n1239, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  AOI22_X1  g0008(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n212));
  NAND4_X1  g0012(.A1(new_n209), .A2(new_n210), .A3(new_n211), .A4(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G20), .ZN(new_n214));
  AND2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(KEYINPUT1), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT64), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n214), .A2(G13), .ZN(new_n219));
  OAI211_X1 g0019(.A(new_n219), .B(G250), .C1(G257), .C2(G264), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT0), .ZN(new_n221));
  AND2_X1   g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(G20), .ZN(new_n223));
  OAI21_X1  g0023(.A(G50), .B1(G58), .B2(G68), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n221), .B1(new_n216), .B2(new_n215), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n218), .A2(new_n225), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT2), .B(G226), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(G264), .B(G270), .Z(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n230), .B(new_n233), .ZN(G358));
  XOR2_X1   g0034(.A(G87), .B(G97), .Z(new_n235));
  XOR2_X1   g0035(.A(G107), .B(G116), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G58), .B(G77), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G351));
  NAND2_X1  g0041(.A1(G20), .A2(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT8), .B(G58), .ZN(new_n243));
  NOR2_X1   g0043(.A1(G20), .A2(G33), .ZN(new_n244));
  INV_X1    g0044(.A(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(G20), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G33), .ZN(new_n247));
  XNOR2_X1  g0047(.A(KEYINPUT15), .B(G87), .ZN(new_n248));
  OAI221_X1 g0048(.A(new_n242), .B1(new_n243), .B2(new_n245), .C1(new_n247), .C2(new_n248), .ZN(new_n249));
  NAND4_X1  g0049(.A1(KEYINPUT66), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G1), .A2(G13), .ZN(new_n251));
  AND2_X1   g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT66), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n253), .B1(new_n214), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G77), .ZN(new_n257));
  INV_X1    g0057(.A(G13), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(G1), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G20), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n249), .A2(new_n256), .B1(new_n257), .B2(new_n261), .ZN(new_n262));
  AND3_X1   g0062(.A1(new_n252), .A2(new_n255), .A3(new_n260), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT69), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n264), .B1(new_n246), .B2(G1), .ZN(new_n265));
  INV_X1    g0065(.A(G1), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n266), .A2(KEYINPUT69), .A3(G20), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n263), .A2(G77), .A3(new_n268), .ZN(new_n269));
  AND2_X1   g0069(.A1(new_n262), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G169), .ZN(new_n271));
  XNOR2_X1  g0071(.A(KEYINPUT3), .B(G33), .ZN(new_n272));
  INV_X1    g0072(.A(G1698), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n272), .A2(G232), .A3(new_n273), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT70), .B(G107), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n272), .A2(G1698), .ZN(new_n276));
  INV_X1    g0076(.A(G238), .ZN(new_n277));
  OAI221_X1 g0077(.A(new_n274), .B1(new_n272), .B2(new_n275), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G33), .A2(G41), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n279), .A2(G1), .A3(G13), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G274), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n283), .B1(new_n222), .B2(new_n279), .ZN(new_n284));
  INV_X1    g0084(.A(G41), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(KEYINPUT65), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT65), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G41), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n284), .B(new_n266), .C1(new_n289), .C2(G45), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n266), .B1(G41), .B2(G45), .ZN(new_n291));
  AND2_X1   g0091(.A1(new_n280), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G244), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n282), .A2(new_n290), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n270), .B1(new_n271), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n295), .B1(G179), .B2(new_n294), .ZN(new_n296));
  AND3_X1   g0096(.A1(new_n255), .A2(new_n251), .A3(new_n250), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT68), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n247), .B(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G58), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n300), .A2(KEYINPUT67), .A3(KEYINPUT8), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT67), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n243), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n299), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  AOI22_X1  g0104(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n244), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n297), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n306), .B1(new_n202), .B2(new_n261), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n263), .A2(G50), .A3(new_n268), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n290), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n310), .B1(G226), .B2(new_n292), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n272), .A2(G222), .A3(new_n273), .ZN(new_n312));
  INV_X1    g0112(.A(G223), .ZN(new_n313));
  OAI221_X1 g0113(.A(new_n312), .B1(new_n257), .B2(new_n272), .C1(new_n276), .C2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n281), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n271), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n309), .B(new_n317), .C1(G179), .C2(new_n316), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n294), .A2(G200), .ZN(new_n319));
  INV_X1    g0119(.A(G190), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n319), .B(new_n270), .C1(new_n320), .C2(new_n294), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n296), .A2(new_n318), .A3(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n316), .A2(new_n320), .ZN(new_n323));
  INV_X1    g0123(.A(G200), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n324), .B1(new_n311), .B2(new_n315), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n309), .A2(KEYINPUT9), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT9), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n328), .B1(new_n307), .B2(new_n308), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n326), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(KEYINPUT10), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT10), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n326), .B(new_n332), .C1(new_n327), .C2(new_n329), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n322), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n280), .A2(G238), .A3(new_n291), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n290), .A2(new_n335), .ZN(new_n336));
  AND2_X1   g0136(.A1(KEYINPUT3), .A2(G33), .ZN(new_n337));
  NOR2_X1   g0137(.A1(KEYINPUT3), .A2(G33), .ZN(new_n338));
  OAI211_X1 g0138(.A(G226), .B(new_n273), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT71), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n272), .A2(KEYINPUT71), .A3(G226), .A4(new_n273), .ZN(new_n342));
  NAND2_X1  g0142(.A1(G33), .A2(G97), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n272), .A2(G232), .A3(G1698), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n341), .A2(new_n342), .A3(new_n343), .A4(new_n344), .ZN(new_n345));
  AOI211_X1 g0145(.A(KEYINPUT13), .B(new_n336), .C1(new_n281), .C2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT13), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n345), .A2(new_n281), .ZN(new_n348));
  INV_X1    g0148(.A(new_n336), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(G169), .B1(new_n346), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT14), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  OAI211_X1 g0153(.A(KEYINPUT14), .B(G169), .C1(new_n346), .C2(new_n350), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n348), .A2(new_n349), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(KEYINPUT72), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n336), .B1(new_n345), .B2(new_n281), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT72), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n357), .A2(KEYINPUT13), .A3(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G179), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n346), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n355), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(G68), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n261), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g0167(.A(new_n367), .B(KEYINPUT12), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n299), .A2(G77), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n244), .A2(G50), .B1(G20), .B2(new_n366), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n297), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n368), .B1(new_n371), .B2(KEYINPUT11), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(KEYINPUT11), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n263), .A2(G68), .A3(new_n268), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n365), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT16), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT7), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(new_n272), .B2(G20), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n337), .A2(new_n338), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n380), .A2(KEYINPUT7), .A3(new_n246), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n366), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n300), .A2(new_n366), .ZN(new_n383));
  OAI21_X1  g0183(.A(G20), .B1(new_n383), .B2(new_n201), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n244), .A2(G159), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n377), .B1(new_n382), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(KEYINPUT7), .B1(new_n380), .B2(new_n246), .ZN(new_n388));
  NOR4_X1   g0188(.A1(new_n337), .A2(new_n338), .A3(new_n378), .A4(G20), .ZN(new_n389));
  OAI21_X1  g0189(.A(G68), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n386), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n390), .A2(KEYINPUT16), .A3(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n387), .A2(new_n392), .A3(new_n256), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n303), .A2(KEYINPUT75), .A3(new_n268), .A4(new_n301), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n394), .A2(new_n263), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT75), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n303), .A2(new_n301), .ZN(new_n397));
  INV_X1    g0197(.A(new_n268), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n395), .A2(new_n399), .B1(new_n261), .B2(new_n397), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n280), .A2(G232), .A3(new_n291), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n290), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n313), .A2(new_n273), .ZN(new_n403));
  INV_X1    g0203(.A(G226), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(G1698), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n403), .B(new_n405), .C1(new_n337), .C2(new_n338), .ZN(new_n406));
  NAND2_X1  g0206(.A1(G33), .A2(G87), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n280), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n324), .B1(new_n402), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n406), .A2(new_n407), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n281), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n411), .A2(new_n320), .A3(new_n290), .A4(new_n401), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  XOR2_X1   g0213(.A(KEYINPUT76), .B(KEYINPUT17), .Z(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n393), .A2(new_n400), .A3(new_n413), .A4(new_n415), .ZN(new_n416));
  AND3_X1   g0216(.A1(new_n393), .A2(new_n400), .A3(new_n413), .ZN(new_n417));
  NOR2_X1   g0217(.A1(KEYINPUT76), .A2(KEYINPUT17), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n416), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n393), .A2(new_n400), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n271), .B1(new_n402), .B2(new_n408), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n411), .A2(new_n362), .A3(new_n290), .A4(new_n401), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT18), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n423), .B1(new_n393), .B2(new_n400), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT18), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n419), .A2(new_n426), .A3(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n334), .A2(new_n376), .A3(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(G200), .B1(new_n346), .B2(new_n350), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n375), .A2(new_n372), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n320), .B1(new_n358), .B2(new_n347), .ZN(new_n436));
  OAI21_X1  g0236(.A(KEYINPUT13), .B1(new_n358), .B2(new_n359), .ZN(new_n437));
  AOI211_X1 g0237(.A(KEYINPUT72), .B(new_n336), .C1(new_n281), .C2(new_n345), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT73), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT73), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n441), .B(new_n436), .C1(new_n437), .C2(new_n438), .ZN(new_n442));
  AOI211_X1 g0242(.A(KEYINPUT74), .B(new_n435), .C1(new_n440), .C2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT74), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n440), .A2(new_n442), .ZN(new_n445));
  AND2_X1   g0245(.A1(new_n433), .A2(new_n434), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n432), .A2(new_n448), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n246), .B(G87), .C1(new_n337), .C2(new_n338), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT22), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT22), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n272), .A2(new_n452), .A3(new_n246), .A4(G87), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n206), .A2(G20), .ZN(new_n455));
  INV_X1    g0255(.A(G116), .ZN(new_n456));
  OAI22_X1  g0256(.A1(KEYINPUT23), .A2(new_n455), .B1(new_n247), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n206), .A2(KEYINPUT70), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT70), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(G107), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n458), .A2(new_n460), .A3(G20), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n457), .B1(KEYINPUT23), .B2(new_n461), .ZN(new_n462));
  XOR2_X1   g0262(.A(KEYINPUT83), .B(KEYINPUT24), .Z(new_n463));
  AND3_X1   g0263(.A1(new_n454), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n463), .B1(new_n454), .B2(new_n462), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n256), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n266), .A2(G33), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n263), .A2(G107), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n259), .A2(G20), .A3(new_n206), .ZN(new_n469));
  XOR2_X1   g0269(.A(new_n469), .B(KEYINPUT25), .Z(new_n470));
  AND2_X1   g0270(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n466), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(G45), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n473), .A2(G1), .ZN(new_n474));
  XNOR2_X1  g0274(.A(KEYINPUT65), .B(G41), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n474), .B1(new_n475), .B2(KEYINPUT5), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT79), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT5), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n477), .B1(new_n478), .B2(G41), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n285), .A2(KEYINPUT79), .A3(KEYINPUT5), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  OAI211_X1 g0282(.A(G264), .B(new_n280), .C1(new_n476), .C2(new_n482), .ZN(new_n483));
  OAI211_X1 g0283(.A(G257), .B(G1698), .C1(new_n337), .C2(new_n338), .ZN(new_n484));
  OAI211_X1 g0284(.A(G250), .B(new_n273), .C1(new_n337), .C2(new_n338), .ZN(new_n485));
  NAND2_X1  g0285(.A1(G33), .A2(G294), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n281), .ZN(new_n488));
  INV_X1    g0288(.A(new_n474), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n489), .B1(new_n289), .B2(new_n478), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n490), .A2(new_n284), .A3(new_n481), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n483), .A2(new_n488), .A3(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n492), .A2(KEYINPUT84), .A3(G169), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n483), .A2(new_n488), .A3(new_n491), .A4(G179), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(KEYINPUT84), .B1(new_n492), .B2(G169), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n472), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT85), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n472), .B(KEYINPUT85), .C1(new_n495), .C2(new_n496), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n483), .A2(new_n488), .A3(new_n491), .A4(G190), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n492), .A2(G200), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n466), .A2(new_n471), .A3(new_n501), .A4(new_n502), .ZN(new_n503));
  AND3_X1   g0303(.A1(new_n499), .A2(new_n500), .A3(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n263), .A2(G116), .A3(new_n467), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n261), .A2(new_n456), .ZN(new_n506));
  AOI21_X1  g0306(.A(G20), .B1(G33), .B2(G283), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n254), .A2(G97), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n507), .A2(new_n508), .B1(G20), .B2(new_n456), .ZN(new_n509));
  AND3_X1   g0309(.A1(new_n256), .A2(KEYINPUT20), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(KEYINPUT20), .B1(new_n256), .B2(new_n509), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n505), .B(new_n506), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n380), .A2(G303), .ZN(new_n513));
  OAI211_X1 g0313(.A(G264), .B(G1698), .C1(new_n337), .C2(new_n338), .ZN(new_n514));
  OAI211_X1 g0314(.A(G257), .B(new_n273), .C1(new_n337), .C2(new_n338), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(KEYINPUT81), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT81), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n513), .A2(new_n518), .A3(new_n514), .A4(new_n515), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n517), .A2(new_n281), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n281), .B1(new_n490), .B2(new_n481), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n476), .A2(new_n482), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n521), .A2(G270), .B1(new_n522), .B2(new_n284), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n512), .A2(G179), .A3(new_n520), .A4(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n271), .B1(new_n523), .B2(new_n520), .ZN(new_n525));
  NOR2_X1   g0325(.A1(KEYINPUT82), .A2(KEYINPUT21), .ZN(new_n526));
  AND3_X1   g0326(.A1(new_n525), .A2(new_n526), .A3(new_n512), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n526), .B1(new_n525), .B2(new_n512), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n524), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n523), .A2(new_n520), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n512), .B1(new_n530), .B2(G200), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n523), .A2(new_n520), .A3(G190), .ZN(new_n532));
  AND2_X1   g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT80), .ZN(new_n535));
  OAI211_X1 g0335(.A(G244), .B(new_n273), .C1(new_n337), .C2(new_n338), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT4), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n272), .A2(KEYINPUT4), .A3(G244), .A4(new_n273), .ZN(new_n539));
  NAND2_X1  g0339(.A1(G33), .A2(G283), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n272), .A2(G250), .A3(G1698), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n538), .A2(new_n539), .A3(new_n540), .A4(new_n541), .ZN(new_n542));
  AND2_X1   g0342(.A1(new_n542), .A2(new_n281), .ZN(new_n543));
  OAI211_X1 g0343(.A(G257), .B(new_n280), .C1(new_n476), .C2(new_n482), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n491), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n535), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n544), .A2(new_n491), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n542), .A2(new_n281), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n547), .A2(KEYINPUT80), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(G190), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT6), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(KEYINPUT77), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT77), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(KEYINPUT6), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n206), .A2(G97), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(G97), .A2(G107), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n207), .A2(new_n553), .A3(new_n555), .A4(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n558), .A2(G20), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n244), .A2(G77), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n275), .B1(new_n379), .B2(new_n381), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n256), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n263), .A2(G97), .A3(new_n467), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n260), .A2(G97), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n565), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n548), .A2(KEYINPUT78), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT78), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n542), .A2(new_n571), .A3(new_n281), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n570), .A2(new_n547), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n569), .B1(new_n573), .B2(G200), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n551), .A2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(G250), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n473), .B2(G1), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n266), .A2(new_n283), .A3(G45), .ZN(new_n578));
  AND3_X1   g0378(.A1(new_n280), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  OAI211_X1 g0379(.A(G244), .B(G1698), .C1(new_n337), .C2(new_n338), .ZN(new_n580));
  OAI211_X1 g0380(.A(G238), .B(new_n273), .C1(new_n337), .C2(new_n338), .ZN(new_n581));
  NAND2_X1  g0381(.A1(G33), .A2(G116), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n579), .B1(new_n583), .B2(new_n281), .ZN(new_n584));
  OR2_X1    g0384(.A1(new_n584), .A2(new_n324), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n246), .B(G68), .C1(new_n337), .C2(new_n338), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT19), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(new_n247), .B2(new_n205), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(G87), .A2(G97), .ZN(new_n590));
  NAND3_X1  g0390(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n275), .A2(new_n590), .B1(new_n246), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n256), .B1(new_n589), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n261), .A2(new_n248), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n297), .A2(G87), .A3(new_n260), .A4(new_n467), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  AOI211_X1 g0396(.A(new_n320), .B(new_n579), .C1(new_n583), .C2(new_n281), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n583), .A2(new_n281), .ZN(new_n599));
  INV_X1    g0399(.A(new_n579), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n599), .A2(G179), .A3(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(new_n271), .B2(new_n584), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n263), .A2(new_n467), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n593), .B(new_n594), .C1(new_n603), .C2(new_n248), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n585), .A2(new_n598), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n542), .A2(new_n571), .A3(new_n281), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n571), .B1(new_n542), .B2(new_n281), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n545), .A2(G179), .ZN(new_n609));
  INV_X1    g0409(.A(new_n275), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n610), .B1(new_n388), .B2(new_n389), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n611), .A2(new_n562), .A3(new_n561), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n567), .B1(new_n612), .B2(new_n256), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n608), .A2(new_n609), .B1(new_n613), .B2(new_n566), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n546), .A2(new_n549), .A3(new_n271), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n575), .A2(new_n605), .A3(new_n616), .ZN(new_n617));
  AND4_X1   g0417(.A1(new_n449), .A2(new_n504), .A3(new_n534), .A4(new_n617), .ZN(G372));
  NAND2_X1  g0418(.A1(new_n426), .A2(new_n429), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n435), .B1(new_n440), .B2(new_n442), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n376), .B1(new_n620), .B2(new_n296), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n619), .B1(new_n621), .B2(new_n419), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n331), .A2(new_n333), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT90), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n331), .A2(KEYINPUT90), .A3(new_n333), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n318), .B1(new_n622), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n614), .A2(new_n605), .A3(KEYINPUT26), .A4(new_n615), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n602), .A2(new_n604), .ZN(new_n632));
  OR3_X1    g0432(.A1(new_n584), .A2(KEYINPUT86), .A3(new_n324), .ZN(new_n633));
  OAI21_X1  g0433(.A(KEYINPUT86), .B1(new_n584), .B2(new_n324), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n598), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n614), .A2(new_n632), .A3(new_n615), .A4(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT26), .ZN(new_n637));
  AOI22_X1  g0437(.A1(KEYINPUT89), .A2(new_n631), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OR2_X1    g0438(.A1(new_n631), .A2(KEYINPUT89), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n638), .A2(new_n639), .B1(new_n604), .B2(new_n602), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT88), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n497), .A2(KEYINPUT87), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT87), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n472), .B(new_n643), .C1(new_n495), .C2(new_n496), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n529), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n503), .A2(new_n632), .A3(new_n635), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n646), .A2(new_n575), .A3(new_n616), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n641), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n646), .A2(new_n575), .A3(new_n616), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n642), .A2(new_n644), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n649), .B(KEYINPUT88), .C1(new_n650), .C2(new_n529), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n640), .A2(new_n648), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n449), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n630), .A2(new_n653), .ZN(G369));
  INV_X1    g0454(.A(G330), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n259), .A2(new_n246), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(G213), .A3(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(G343), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n512), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n534), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n529), .A2(new_n512), .A3(new_n661), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n655), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  XNOR2_X1  g0465(.A(new_n665), .B(KEYINPUT91), .ZN(new_n666));
  INV_X1    g0466(.A(new_n661), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n497), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n472), .A2(new_n661), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n669), .B1(new_n504), .B2(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n666), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n504), .A2(new_n529), .A3(new_n667), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n650), .A2(new_n667), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n672), .A2(new_n675), .ZN(G399));
  INV_X1    g0476(.A(new_n219), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(new_n289), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n275), .A2(new_n456), .A3(new_n590), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n679), .A2(G1), .A3(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(new_n224), .B2(new_n679), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT28), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT29), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n652), .A2(new_n685), .A3(new_n667), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n499), .A2(new_n500), .ZN(new_n687));
  INV_X1    g0487(.A(new_n529), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n647), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n614), .A2(new_n605), .A3(new_n615), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT93), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(new_n691), .A3(new_n637), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n635), .A2(new_n632), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n693), .A2(KEYINPUT26), .A3(new_n615), .A4(new_n614), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n691), .B1(new_n690), .B2(new_n637), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n632), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n689), .B1(new_n697), .B2(KEYINPUT94), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT94), .ZN(new_n699));
  OAI211_X1 g0499(.A(new_n699), .B(new_n632), .C1(new_n695), .C2(new_n696), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n661), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n686), .B1(new_n701), .B2(new_n685), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n504), .A2(new_n617), .A3(new_n534), .A4(new_n667), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n483), .A2(new_n488), .ZN(new_n705));
  AOI211_X1 g0505(.A(new_n362), .B(new_n579), .C1(new_n583), .C2(new_n281), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n523), .A2(new_n705), .A3(new_n520), .A4(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n707), .B1(new_n546), .B2(new_n549), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(KEYINPUT30), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n584), .ZN(new_n711));
  AND3_X1   g0511(.A1(new_n492), .A2(new_n362), .A3(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n573), .A2(new_n712), .A3(new_n530), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n708), .B2(KEYINPUT30), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n661), .B1(new_n710), .B2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT31), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AND4_X1   g0517(.A1(new_n705), .A2(new_n523), .A3(new_n520), .A4(new_n706), .ZN(new_n718));
  AOI21_X1  g0518(.A(KEYINPUT30), .B1(new_n550), .B2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n713), .ZN(new_n720));
  OAI21_X1  g0520(.A(KEYINPUT92), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT92), .ZN(new_n722));
  OAI211_X1 g0522(.A(new_n722), .B(new_n713), .C1(new_n708), .C2(KEYINPUT30), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n721), .A2(new_n709), .A3(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n667), .A2(new_n716), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n704), .A2(new_n717), .A3(new_n726), .ZN(new_n727));
  AND2_X1   g0527(.A1(new_n727), .A2(G330), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n703), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n684), .B1(new_n731), .B2(G1), .ZN(G364));
  NOR2_X1   g0532(.A1(new_n258), .A2(G20), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n266), .B1(new_n733), .B2(G45), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n679), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n663), .A2(new_n655), .A3(new_n664), .ZN(new_n736));
  XNOR2_X1  g0536(.A(new_n736), .B(KEYINPUT95), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n666), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  XOR2_X1   g0538(.A(new_n738), .B(KEYINPUT96), .Z(new_n739));
  NOR2_X1   g0539(.A1(G13), .A2(G33), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(new_n246), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n741), .B(KEYINPUT98), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n663), .A2(new_n664), .A3(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n246), .A2(G179), .ZN(new_n745));
  NOR2_X1   g0545(.A1(G190), .A2(G200), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  AND2_X1   g0548(.A1(new_n748), .A2(G329), .ZN(new_n749));
  XOR2_X1   g0549(.A(KEYINPUT33), .B(G317), .Z(new_n750));
  NOR2_X1   g0550(.A1(new_n246), .A2(new_n362), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n324), .A2(G190), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n745), .A2(new_n752), .ZN(new_n754));
  INV_X1    g0554(.A(G283), .ZN(new_n755));
  OAI22_X1  g0555(.A1(new_n750), .A2(new_n753), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n751), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n757), .A2(new_n320), .A3(G200), .ZN(new_n758));
  AOI211_X1 g0558(.A(new_n749), .B(new_n756), .C1(G322), .C2(new_n758), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n320), .A2(G179), .A3(G200), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n246), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G294), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n320), .A2(new_n324), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n751), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n272), .B1(new_n766), .B2(G326), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n751), .A2(new_n746), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n764), .A2(new_n745), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI22_X1  g0571(.A1(G311), .A2(new_n769), .B1(new_n771), .B2(G303), .ZN(new_n772));
  AND4_X1   g0572(.A1(new_n759), .A2(new_n763), .A3(new_n767), .A4(new_n772), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n773), .A2(KEYINPUT100), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(KEYINPUT100), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n765), .A2(new_n202), .B1(new_n768), .B2(new_n257), .ZN(new_n776));
  INV_X1    g0576(.A(new_n753), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n380), .B(new_n776), .C1(G68), .C2(new_n777), .ZN(new_n778));
  XOR2_X1   g0578(.A(KEYINPUT99), .B(KEYINPUT32), .Z(new_n779));
  NAND3_X1  g0579(.A1(new_n748), .A2(G159), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n779), .B1(new_n748), .B2(G159), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n781), .B1(G97), .B2(new_n762), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n754), .A2(new_n206), .ZN(new_n783));
  INV_X1    g0583(.A(G87), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n770), .A2(new_n784), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n783), .B(new_n785), .C1(G58), .C2(new_n758), .ZN(new_n786));
  NAND4_X1  g0586(.A1(new_n778), .A2(new_n780), .A3(new_n782), .A4(new_n786), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n774), .A2(new_n775), .A3(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n251), .B1(G20), .B2(new_n271), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n743), .A2(new_n789), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n677), .A2(new_n380), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT97), .ZN(new_n793));
  INV_X1    g0593(.A(G355), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n793), .A2(new_n794), .B1(G116), .B2(new_n219), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n677), .A2(new_n272), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(G45), .B2(new_n224), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n797), .B1(G45), .B2(new_n240), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n791), .B1(new_n795), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n735), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n744), .A2(new_n790), .A3(new_n799), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n739), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(KEYINPUT101), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n802), .B(new_n803), .ZN(G396));
  NOR2_X1   g0604(.A1(new_n789), .A2(new_n740), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n735), .B1(new_n257), .B2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n789), .ZN(new_n807));
  INV_X1    g0607(.A(new_n754), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n272), .B1(new_n808), .B2(G87), .ZN(new_n809));
  INV_X1    g0609(.A(new_n758), .ZN(new_n810));
  INV_X1    g0610(.A(G294), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n809), .B1(new_n755), .B2(new_n753), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n766), .A2(G303), .B1(new_n748), .B2(G311), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n813), .B1(new_n206), .B2(new_n770), .C1(new_n456), .C2(new_n768), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n812), .B(new_n814), .C1(G97), .C2(new_n762), .ZN(new_n815));
  INV_X1    g0615(.A(G137), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n765), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(G143), .ZN(new_n818));
  INV_X1    g0618(.A(G159), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n810), .A2(new_n818), .B1(new_n768), .B2(new_n819), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n817), .B(new_n820), .C1(G150), .C2(new_n777), .ZN(new_n821));
  OR2_X1    g0621(.A1(new_n821), .A2(KEYINPUT34), .ZN(new_n822));
  AOI22_X1  g0622(.A1(G50), .A2(new_n771), .B1(new_n748), .B2(G132), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n380), .B1(new_n808), .B2(G68), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n823), .B(new_n824), .C1(new_n300), .C2(new_n761), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(new_n821), .B2(KEYINPUT34), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n815), .B1(new_n822), .B2(new_n826), .ZN(new_n827));
  OR2_X1    g0627(.A1(new_n296), .A2(new_n661), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n321), .B1(new_n270), .B2(new_n667), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(new_n296), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n740), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n806), .B1(new_n807), .B2(new_n827), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n652), .A2(new_n667), .ZN(new_n835));
  INV_X1    g0635(.A(new_n831), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n652), .A2(new_n667), .A3(new_n831), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n840), .A2(new_n728), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT102), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n735), .B1(new_n839), .B2(new_n729), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n841), .A2(new_n842), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n834), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(G384));
  NAND2_X1  g0648(.A1(new_n697), .A2(KEYINPUT94), .ZN(new_n849));
  INV_X1    g0649(.A(new_n689), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n849), .A2(new_n700), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n685), .B1(new_n851), .B2(new_n667), .ZN(new_n852));
  INV_X1    g0652(.A(new_n686), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n449), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n630), .ZN(new_n855));
  XOR2_X1   g0655(.A(new_n855), .B(KEYINPUT105), .Z(new_n856));
  AOI22_X1  g0656(.A1(new_n353), .A2(new_n354), .B1(new_n361), .B2(new_n363), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n857), .A2(new_n434), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n661), .B1(new_n375), .B2(new_n372), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NOR3_X1   g0660(.A1(new_n858), .A2(new_n620), .A3(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n857), .B1(new_n443), .B2(new_n447), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n861), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n863), .B1(new_n838), .B2(new_n828), .ZN(new_n864));
  INV_X1    g0664(.A(new_n659), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n420), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n430), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n393), .A2(new_n400), .A3(new_n413), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n425), .A2(new_n866), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(KEYINPUT37), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n417), .A2(new_n427), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT37), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n872), .A2(new_n873), .A3(new_n866), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n868), .A2(new_n875), .A3(KEYINPUT38), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT38), .B1(new_n868), .B2(new_n875), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n864), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT39), .ZN(new_n880));
  NOR3_X1   g0680(.A1(new_n877), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT104), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n868), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT103), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n870), .A2(KEYINPUT37), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n873), .B1(new_n872), .B2(new_n866), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n884), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n871), .A2(new_n874), .A3(KEYINPUT103), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n430), .A2(KEYINPUT104), .A3(new_n867), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n883), .A2(new_n887), .A3(new_n888), .A4(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT38), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n876), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n881), .B1(new_n893), .B2(new_n880), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n858), .A2(new_n667), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n619), .A2(new_n659), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n879), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n856), .B(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n441), .B1(new_n361), .B2(new_n436), .ZN(new_n901));
  INV_X1    g0701(.A(new_n442), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n446), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n376), .A2(new_n903), .A3(new_n859), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(KEYINPUT74), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n620), .A2(new_n444), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n365), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n904), .B1(new_n907), .B2(new_n859), .ZN(new_n908));
  OAI211_X1 g0708(.A(KEYINPUT31), .B(new_n661), .C1(new_n710), .C2(new_n714), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n704), .A2(new_n717), .A3(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n908), .A2(new_n831), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n877), .B1(new_n890), .B2(new_n891), .ZN(new_n912));
  OAI21_X1  g0712(.A(KEYINPUT40), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n878), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT40), .B1(new_n914), .B2(new_n876), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n915), .A2(new_n831), .A3(new_n908), .A4(new_n910), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n449), .A2(new_n910), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n917), .A2(new_n918), .ZN(new_n921));
  NOR3_X1   g0721(.A1(new_n920), .A2(new_n921), .A3(new_n655), .ZN(new_n922));
  OAI22_X1  g0722(.A1(new_n900), .A2(new_n922), .B1(new_n266), .B2(new_n733), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n923), .B1(new_n900), .B2(new_n922), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n223), .A2(new_n456), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n558), .A2(new_n560), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT35), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n928), .B1(new_n927), .B2(new_n926), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT36), .ZN(new_n930));
  OR3_X1    g0730(.A1(new_n383), .A2(new_n224), .A3(new_n257), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n202), .A2(G68), .ZN(new_n932));
  AOI211_X1 g0732(.A(new_n266), .B(G13), .C1(new_n931), .C2(new_n932), .ZN(new_n933));
  OR3_X1    g0733(.A1(new_n924), .A2(new_n930), .A3(new_n933), .ZN(G367));
  NAND2_X1  g0734(.A1(new_n569), .A2(new_n661), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n575), .A2(new_n616), .A3(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n614), .A2(new_n615), .A3(new_n661), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n673), .A2(new_n938), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n939), .B(KEYINPUT42), .Z(new_n940));
  OAI21_X1  g0740(.A(new_n616), .B1(new_n687), .B2(new_n936), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n940), .B1(new_n667), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n596), .A2(new_n661), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n693), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n632), .B2(new_n943), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT106), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n946), .A2(KEYINPUT43), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(KEYINPUT43), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n945), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n942), .A2(new_n949), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n950), .B(KEYINPUT107), .Z(new_n951));
  AND2_X1   g0751(.A1(new_n945), .A2(KEYINPUT43), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n951), .B1(new_n942), .B2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n672), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n955), .A2(new_n938), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n954), .B(new_n956), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n678), .B(KEYINPUT41), .Z(new_n958));
  INV_X1    g0758(.A(KEYINPUT111), .ZN(new_n959));
  OR3_X1    g0759(.A1(new_n675), .A2(KEYINPUT108), .A3(new_n938), .ZN(new_n960));
  OAI21_X1  g0760(.A(KEYINPUT108), .B1(new_n675), .B2(new_n938), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AND2_X1   g0762(.A1(new_n962), .A2(KEYINPUT45), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n962), .A2(KEYINPUT45), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n675), .A2(new_n938), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT110), .ZN(new_n967));
  XOR2_X1   g0767(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n967), .A2(new_n968), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n965), .A2(new_n955), .A3(new_n969), .A4(new_n970), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n970), .B(new_n969), .C1(new_n963), .C2(new_n964), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n672), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n671), .B1(new_n688), .B2(new_n661), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n673), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n666), .B(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n730), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n959), .B1(new_n974), .B2(new_n979), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n971), .A2(new_n973), .A3(KEYINPUT111), .A4(new_n978), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n958), .B1(new_n982), .B2(new_n731), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n734), .B(KEYINPUT112), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n957), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  NOR3_X1   g0786(.A1(new_n233), .A2(new_n677), .A3(new_n272), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n791), .B1(new_n219), .B2(new_n248), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n765), .A2(new_n818), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n770), .A2(new_n300), .B1(new_n754), .B2(new_n257), .ZN(new_n990));
  AOI211_X1 g0790(.A(new_n989), .B(new_n990), .C1(G150), .C2(new_n758), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n768), .A2(new_n202), .B1(new_n747), .B2(new_n816), .ZN(new_n992));
  AOI211_X1 g0792(.A(new_n380), .B(new_n992), .C1(G159), .C2(new_n777), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n991), .B(new_n993), .C1(new_n366), .C2(new_n761), .ZN(new_n994));
  INV_X1    g0794(.A(G317), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n753), .A2(new_n811), .B1(new_n747), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(G311), .B2(new_n766), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n272), .B1(new_n808), .B2(G97), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n758), .A2(G303), .B1(G283), .B2(new_n769), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n771), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT46), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n770), .B2(new_n456), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n1001), .B(new_n1003), .C1(new_n275), .C2(new_n761), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n994), .B1(new_n1000), .B2(new_n1004), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n1005), .B(KEYINPUT47), .Z(new_n1006));
  OAI221_X1 g0806(.A(new_n800), .B1(new_n987), .B2(new_n988), .C1(new_n1006), .C2(new_n807), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1007), .B(KEYINPUT113), .Z(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(new_n742), .B2(new_n945), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n986), .A2(new_n1009), .ZN(G387));
  NAND2_X1  g0810(.A1(new_n730), .A2(new_n977), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n979), .A2(new_n678), .A3(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n796), .B1(new_n230), .B2(new_n473), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n681), .B2(new_n793), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n243), .A2(G50), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT50), .ZN(new_n1016));
  AOI21_X1  g0816(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1016), .A2(new_n681), .A3(new_n1017), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n1014), .A2(new_n1018), .B1(new_n206), .B2(new_n677), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n791), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n800), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n758), .A2(G317), .B1(G303), .B2(new_n769), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(G322), .A2(new_n766), .B1(new_n777), .B2(G311), .ZN(new_n1023));
  AND2_X1   g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  AND2_X1   g0824(.A1(new_n1024), .A2(KEYINPUT48), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n1024), .A2(KEYINPUT48), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n761), .A2(new_n755), .B1(new_n770), .B2(new_n811), .ZN(new_n1027));
  NOR3_X1   g0827(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n1028), .A2(KEYINPUT49), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(KEYINPUT49), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n380), .B1(new_n754), .B2(new_n456), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(G326), .B2(new_n748), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1029), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(G159), .A2(new_n766), .B1(new_n769), .B2(G68), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n202), .B2(new_n810), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n761), .A2(new_n248), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n272), .B1(new_n754), .B2(new_n205), .ZN(new_n1037));
  NOR3_X1   g0837(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(G150), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n770), .A2(new_n257), .B1(new_n747), .B2(new_n1039), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT114), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1038), .B(new_n1041), .C1(new_n397), .C2(new_n753), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n807), .B1(new_n1033), .B2(new_n1042), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1021), .B(new_n1043), .C1(new_n671), .C2(new_n743), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n977), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1044), .B1(new_n1045), .B2(new_n985), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1012), .A2(new_n1046), .ZN(G393));
  AOI21_X1  g0847(.A(new_n679), .B1(new_n974), .B2(new_n979), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n982), .A2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n971), .A2(new_n973), .A3(new_n985), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n791), .B1(new_n205), .B2(new_n219), .ZN(new_n1051));
  AND2_X1   g0851(.A1(new_n237), .A2(new_n796), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n800), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n758), .A2(G159), .B1(new_n766), .B2(G150), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT51), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n272), .B1(new_n754), .B2(new_n784), .C1(new_n761), .C2(new_n257), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n202), .A2(new_n753), .B1(new_n770), .B2(new_n366), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n768), .A2(new_n243), .B1(new_n747), .B2(new_n818), .ZN(new_n1058));
  OR3_X1    g0858(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n758), .A2(G311), .B1(new_n766), .B2(G317), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT52), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n272), .B(new_n783), .C1(G116), .C2(new_n762), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(G283), .A2(new_n771), .B1(new_n777), .B2(G303), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(G294), .A2(new_n769), .B1(new_n748), .B2(G322), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n1055), .A2(new_n1059), .B1(new_n1061), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1053), .B1(new_n1066), .B2(new_n789), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n938), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1067), .B1(new_n1068), .B2(new_n742), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1050), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1049), .A2(new_n1071), .ZN(G390));
  XNOR2_X1  g0872(.A(new_n895), .B(KEYINPUT115), .ZN(new_n1073));
  AND2_X1   g0873(.A1(new_n893), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n828), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(new_n701), .B2(new_n830), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT116), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n908), .A2(new_n1077), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n904), .B(KEYINPUT116), .C1(new_n907), .C2(new_n859), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1074), .B1(new_n1076), .B2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n912), .A2(KEYINPUT39), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n864), .A2(new_n896), .B1(new_n1082), .B2(new_n881), .ZN(new_n1083));
  AND3_X1   g0883(.A1(new_n727), .A2(G330), .A3(new_n831), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(new_n908), .ZN(new_n1085));
  AND3_X1   g0885(.A1(new_n1081), .A2(new_n1083), .A3(new_n1085), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n908), .A2(G330), .A3(new_n831), .A4(new_n910), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n985), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n735), .B1(new_n397), .B2(new_n805), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(G50), .A2(new_n808), .B1(new_n748), .B2(G125), .ZN(new_n1092));
  INV_X1    g0892(.A(G128), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1092), .B1(new_n1093), .B2(new_n765), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT53), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n770), .A2(new_n1039), .ZN(new_n1096));
  INV_X1    g0896(.A(G132), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n272), .B1(new_n1095), .B2(new_n1096), .C1(new_n810), .C2(new_n1097), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n1094), .B(new_n1098), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(KEYINPUT54), .B(G143), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n816), .A2(new_n753), .B1(new_n768), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(G159), .B2(new_n762), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT118), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(G116), .A2(new_n758), .B1(new_n762), .B2(G77), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT119), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(G97), .A2(new_n769), .B1(new_n748), .B2(G294), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1106), .B1(new_n755), .B2(new_n765), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n753), .A2(new_n275), .B1(new_n754), .B2(new_n366), .ZN(new_n1108));
  NOR4_X1   g0908(.A1(new_n1107), .A2(new_n272), .A3(new_n785), .A4(new_n1108), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n1099), .A2(new_n1103), .B1(new_n1105), .B2(new_n1109), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n1091), .B1(new_n807), .B2(new_n1110), .C1(new_n894), .C2(new_n832), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1090), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n727), .A2(G330), .A3(new_n831), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n863), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1114), .A2(new_n1087), .B1(new_n828), .B2(new_n838), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n910), .A2(G330), .A3(new_n831), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n1080), .A2(new_n1116), .B1(new_n908), .B2(new_n1084), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1115), .B1(new_n1117), .B2(new_n1076), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n449), .A2(G330), .A3(new_n910), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n854), .A2(new_n630), .A3(new_n1119), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1087), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n838), .A2(new_n828), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n908), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n894), .B1(new_n1124), .B2(new_n895), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n893), .A2(new_n1073), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n851), .A2(new_n667), .A3(new_n830), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n828), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1080), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1126), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1122), .B1(new_n1125), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1081), .A2(new_n1083), .A3(new_n1085), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1121), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT117), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1121), .A2(new_n1131), .A3(KEYINPUT117), .A4(new_n1132), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1121), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n679), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1112), .B1(new_n1137), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(G378));
  NAND2_X1  g0942(.A1(new_n309), .A2(new_n865), .ZN(new_n1143));
  AND3_X1   g0943(.A1(new_n627), .A2(new_n318), .A3(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1143), .B1(new_n627), .B2(new_n318), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  OR3_X1    g0947(.A1(new_n1144), .A2(new_n1145), .A3(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1147), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1148), .A2(new_n740), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n766), .A2(G125), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n1151), .B1(new_n770), .B2(new_n1100), .C1(new_n810), .C2(new_n1093), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n1097), .A2(new_n753), .B1(new_n768), .B2(new_n816), .ZN(new_n1153));
  XOR2_X1   g0953(.A(new_n1153), .B(KEYINPUT122), .Z(new_n1154));
  AOI211_X1 g0954(.A(new_n1152), .B(new_n1154), .C1(G150), .C2(new_n762), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  OR2_X1    g0956(.A1(new_n1156), .A2(KEYINPUT59), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(KEYINPUT59), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n254), .B(new_n285), .C1(new_n754), .C2(new_n819), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(G124), .B2(new_n748), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1157), .A2(new_n1158), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n380), .A2(new_n475), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n754), .A2(new_n300), .B1(new_n747), .B2(new_n755), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n1162), .B(new_n1163), .C1(G77), .C2(new_n771), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT121), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n765), .A2(new_n456), .B1(new_n753), .B2(new_n205), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n810), .A2(new_n206), .B1(new_n248), .B2(new_n768), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n1166), .B(new_n1167), .C1(G68), .C2(new_n762), .ZN(new_n1168));
  AND2_X1   g0968(.A1(new_n1165), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(KEYINPUT58), .ZN(new_n1170));
  OR2_X1    g0970(.A1(new_n1169), .A2(KEYINPUT58), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1162), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1172));
  XOR2_X1   g0972(.A(new_n1172), .B(KEYINPUT120), .Z(new_n1173));
  NAND4_X1  g0973(.A1(new_n1161), .A2(new_n1170), .A3(new_n1171), .A4(new_n1173), .ZN(new_n1174));
  AND2_X1   g0974(.A1(new_n1174), .A2(new_n789), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n735), .B(new_n1175), .C1(new_n202), .C2(new_n805), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1150), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n655), .B1(new_n913), .B2(new_n916), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT123), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1178), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  AOI211_X1 g0981(.A(KEYINPUT123), .B(new_n655), .C1(new_n913), .C2(new_n916), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n917), .A2(G330), .ZN(new_n1184));
  NOR3_X1   g0984(.A1(new_n1184), .A2(new_n1178), .A3(KEYINPUT123), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n899), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1184), .A2(KEYINPUT123), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1187), .A2(new_n1188), .A3(new_n1178), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n899), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1186), .A2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1177), .B1(new_n1193), .B2(new_n984), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1119), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n629), .B(new_n1196), .C1(new_n702), .C2(new_n449), .ZN(new_n1197));
  AOI21_X1  g0997(.A(KEYINPUT117), .B1(new_n1089), .B2(new_n1121), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1136), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1197), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  AND2_X1   g1000(.A1(new_n1186), .A2(new_n1192), .ZN(new_n1201));
  AOI21_X1  g1001(.A(KEYINPUT57), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1120), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1186), .A2(new_n1192), .A3(KEYINPUT57), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n678), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1195), .B1(new_n1202), .B2(new_n1205), .ZN(G375));
  OAI22_X1  g1006(.A1(new_n810), .A2(new_n755), .B1(new_n765), .B2(new_n811), .ZN(new_n1207));
  INV_X1    g1007(.A(G303), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n770), .A2(new_n205), .B1(new_n747), .B2(new_n1208), .ZN(new_n1209));
  NOR3_X1   g1009(.A1(new_n1207), .A2(new_n1209), .A3(new_n1036), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n380), .B1(new_n754), .B2(new_n257), .ZN(new_n1211));
  XOR2_X1   g1011(.A(new_n1211), .B(KEYINPUT125), .Z(new_n1212));
  OAI22_X1  g1012(.A1(new_n456), .A2(new_n753), .B1(new_n768), .B2(new_n275), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT124), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1210), .A2(new_n1212), .A3(new_n1214), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n765), .A2(new_n1097), .B1(new_n753), .B2(new_n1100), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n380), .B(new_n1216), .C1(G58), .C2(new_n808), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n770), .A2(new_n819), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n768), .A2(new_n1039), .B1(new_n747), .B2(new_n1093), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n1218), .B(new_n1219), .C1(G137), .C2(new_n758), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1217), .B(new_n1220), .C1(new_n202), .C2(new_n761), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n807), .B1(new_n1215), .B2(new_n1221), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n735), .B(new_n1222), .C1(new_n366), .C2(new_n805), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(new_n1129), .B2(new_n832), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1224), .B1(new_n1118), .B2(new_n984), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1121), .A2(new_n958), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1225), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(G381));
  OR2_X1    g1029(.A1(G396), .A2(G393), .ZN(new_n1230));
  OR3_X1    g1030(.A1(G390), .A2(G384), .A3(new_n1230), .ZN(new_n1231));
  NOR3_X1   g1031(.A1(new_n1231), .A2(G387), .A3(G381), .ZN(new_n1232));
  INV_X1    g1032(.A(G375), .ZN(new_n1233));
  OR2_X1    g1033(.A1(new_n1233), .A2(KEYINPUT126), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(KEYINPUT126), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1232), .A2(new_n1141), .A3(new_n1234), .A4(new_n1235), .ZN(G407));
  NAND2_X1  g1036(.A1(new_n660), .A2(G213), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1234), .A2(new_n1141), .A3(new_n1235), .A4(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(G407), .A2(G213), .A3(new_n1239), .ZN(G409));
  NAND2_X1  g1040(.A1(new_n1238), .A2(G2897), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT60), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1079), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n862), .A2(new_n860), .ZN(new_n1245));
  AOI21_X1  g1045(.A(KEYINPUT116), .B1(new_n1245), .B2(new_n904), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1116), .B1(new_n1244), .B2(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1076), .A2(new_n1247), .A3(new_n1085), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1115), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1243), .B1(new_n1250), .B2(new_n1197), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1250), .A2(new_n1197), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n678), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  OAI21_X1  g1053(.A(KEYINPUT60), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1254), .A2(new_n1227), .ZN(new_n1255));
  OAI21_X1  g1055(.A(KEYINPUT127), .B1(new_n1253), .B2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n679), .B1(new_n1254), .B2(new_n1227), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT127), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1257), .A2(new_n1258), .A3(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1256), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1225), .ZN(new_n1262));
  AOI21_X1  g1062(.A(G384), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  AOI211_X1 g1063(.A(new_n847), .B(new_n1225), .C1(new_n1256), .C2(new_n1260), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1242), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  NOR3_X1   g1065(.A1(new_n1253), .A2(new_n1255), .A3(KEYINPUT127), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1258), .B1(new_n1257), .B2(new_n1259), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1262), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n847), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1261), .A2(G384), .A3(new_n1262), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1269), .A2(new_n1270), .A3(new_n1241), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1265), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  OAI211_X1 g1073(.A(G378), .B(new_n1195), .C1(new_n1202), .C2(new_n1205), .ZN(new_n1274));
  NOR3_X1   g1074(.A1(new_n1203), .A2(new_n958), .A3(new_n1193), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1141), .B1(new_n1275), .B2(new_n1194), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1274), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n1237), .ZN(new_n1278));
  AOI21_X1  g1078(.A(KEYINPUT61), .B1(new_n1273), .B2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT63), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1280), .B1(new_n1278), .B2(new_n1282), .ZN(new_n1283));
  AND2_X1   g1083(.A1(new_n1012), .A2(new_n1046), .ZN(new_n1284));
  XNOR2_X1  g1084(.A(G396), .B(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(G390), .A2(new_n1285), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(G396), .B(G393), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1287), .A2(new_n1049), .A3(new_n1071), .ZN(new_n1288));
  AND4_X1   g1088(.A1(new_n986), .A2(new_n1286), .A3(new_n1009), .A4(new_n1288), .ZN(new_n1289));
  AOI22_X1  g1089(.A1(new_n1286), .A2(new_n1288), .B1(new_n986), .B2(new_n1009), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1238), .B1(new_n1274), .B2(new_n1276), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1292), .A2(KEYINPUT63), .A3(new_n1281), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1279), .A2(new_n1283), .A3(new_n1291), .A4(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT62), .ZN(new_n1295));
  AND3_X1   g1095(.A1(new_n1292), .A2(new_n1295), .A3(new_n1281), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT61), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1297), .B1(new_n1292), .B2(new_n1272), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1295), .B1(new_n1292), .B2(new_n1281), .ZN(new_n1299));
  NOR3_X1   g1099(.A1(new_n1296), .A2(new_n1298), .A3(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1294), .B1(new_n1300), .B2(new_n1291), .ZN(G405));
  OR2_X1    g1101(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(G375), .A2(new_n1141), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(new_n1274), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n1281), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1282), .A2(new_n1303), .A3(new_n1274), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  XNOR2_X1  g1107(.A(new_n1302), .B(new_n1307), .ZN(G402));
endmodule


