//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 1 1 0 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 1 0 1 0 1 0 1 1 1 1 0 0 0 0 1 1 0 0 1 1 1 1 0 0 0 0 0 0 1 0 1 1 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:27 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n763, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G107), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G104), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT78), .ZN(new_n192));
  INV_X1    g006(.A(G104), .ZN(new_n193));
  OAI211_X1 g007(.A(new_n192), .B(KEYINPUT3), .C1(new_n193), .C2(G107), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n189), .A2(G104), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n192), .B1(new_n196), .B2(KEYINPUT3), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n191), .B1(new_n195), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT3), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n199), .A2(new_n189), .A3(G104), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT79), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT79), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n202), .A2(new_n199), .A3(new_n189), .A4(G104), .ZN(new_n203));
  AND2_X1   g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  OAI21_X1  g018(.A(G101), .B1(new_n198), .B2(new_n204), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT3), .B1(new_n193), .B2(G107), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT78), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(new_n194), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n201), .A2(new_n203), .ZN(new_n209));
  INV_X1    g023(.A(G101), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n208), .A2(new_n209), .A3(new_n210), .A4(new_n191), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n205), .A2(KEYINPUT4), .A3(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G119), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT66), .B1(new_n213), .B2(G116), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT66), .ZN(new_n215));
  INV_X1    g029(.A(G116), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n215), .A2(new_n216), .A3(G119), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n216), .A2(G119), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT67), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n219), .B1(new_n214), .B2(new_n217), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT67), .ZN(new_n225));
  XNOR2_X1  g039(.A(KEYINPUT2), .B(G113), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n223), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n221), .A2(new_n226), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  XOR2_X1   g044(.A(KEYINPUT80), .B(KEYINPUT4), .Z(new_n231));
  OAI211_X1 g045(.A(G101), .B(new_n231), .C1(new_n198), .C2(new_n204), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n212), .A2(new_n230), .A3(new_n232), .ZN(new_n233));
  AOI211_X1 g047(.A(new_n222), .B(new_n219), .C1(new_n217), .C2(new_n214), .ZN(new_n234));
  AOI21_X1  g048(.A(KEYINPUT67), .B1(new_n218), .B2(new_n220), .ZN(new_n235));
  OAI21_X1  g049(.A(KEYINPUT5), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(G113), .B1(new_n220), .B2(KEYINPUT5), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n191), .A2(new_n196), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G101), .ZN(new_n241));
  AND2_X1   g055(.A1(new_n211), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n239), .A2(new_n242), .A3(new_n229), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n233), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g058(.A(G110), .B(G122), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n233), .A2(new_n243), .A3(new_n245), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n247), .A2(KEYINPUT6), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G146), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G143), .ZN(new_n251));
  INV_X1    g065(.A(G143), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G146), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT1), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n251), .A2(new_n253), .A3(new_n254), .A4(G128), .ZN(new_n255));
  INV_X1    g069(.A(G128), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n256), .B1(new_n251), .B2(KEYINPUT1), .ZN(new_n257));
  XNOR2_X1  g071(.A(G143), .B(G146), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n255), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G125), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT0), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(new_n256), .ZN(new_n263));
  NAND2_X1  g077(.A1(KEYINPUT0), .A2(G128), .ZN(new_n264));
  AOI22_X1  g078(.A1(new_n251), .A2(new_n253), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n251), .A2(new_n253), .A3(new_n264), .ZN(new_n266));
  OAI21_X1  g080(.A(G125), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n261), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G953), .ZN(new_n269));
  AND2_X1   g083(.A1(new_n269), .A2(G224), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n269), .A2(G224), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n261), .A2(new_n272), .A3(new_n267), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n244), .A2(new_n275), .A3(new_n246), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n249), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n211), .A2(new_n241), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n223), .A2(new_n225), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n237), .B1(new_n279), .B2(KEYINPUT5), .ZN(new_n280));
  OAI211_X1 g094(.A(KEYINPUT83), .B(new_n278), .C1(new_n280), .C2(new_n228), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT83), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n228), .B1(new_n236), .B2(new_n238), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n282), .B1(new_n283), .B2(new_n242), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n237), .B1(new_n224), .B2(KEYINPUT5), .ZN(new_n285));
  OR3_X1    g099(.A1(new_n278), .A2(new_n228), .A3(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n281), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n245), .B(KEYINPUT8), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT7), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n272), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n271), .A2(new_n273), .A3(new_n291), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n261), .A2(new_n290), .A3(new_n267), .A4(new_n272), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n190), .B1(new_n207), .B2(new_n194), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n210), .B1(new_n295), .B2(new_n209), .ZN(new_n296));
  AOI22_X1  g110(.A1(new_n227), .A2(new_n229), .B1(new_n296), .B2(new_n231), .ZN(new_n297));
  AOI22_X1  g111(.A1(new_n297), .A2(new_n212), .B1(new_n283), .B2(new_n242), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n294), .B1(new_n298), .B2(new_n245), .ZN(new_n299));
  AOI21_X1  g113(.A(G902), .B1(new_n289), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n277), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(G210), .B1(G237), .B2(G902), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(KEYINPUT84), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n277), .A2(new_n300), .A3(new_n304), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n188), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT9), .B(G234), .ZN(new_n309));
  OAI21_X1  g123(.A(G221), .B1(new_n309), .B2(G902), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT82), .ZN(new_n312));
  INV_X1    g126(.A(new_n259), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n278), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n251), .A2(new_n253), .ZN(new_n315));
  OAI211_X1 g129(.A(KEYINPUT81), .B(KEYINPUT1), .C1(new_n252), .C2(G146), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G128), .ZN(new_n317));
  AOI21_X1  g131(.A(KEYINPUT81), .B1(new_n251), .B2(KEYINPUT1), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n315), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(new_n255), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(new_n211), .A3(new_n241), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n314), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(KEYINPUT65), .A2(G131), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G134), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G137), .ZN(new_n326));
  INV_X1    g140(.A(G137), .ZN(new_n327));
  AOI21_X1  g141(.A(KEYINPUT64), .B1(new_n327), .B2(G134), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT11), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n326), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT64), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n331), .B1(new_n325), .B2(G137), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n332), .A2(KEYINPUT11), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n324), .B1(new_n330), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n332), .A2(KEYINPUT11), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n327), .A2(G134), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n336), .A2(new_n331), .A3(new_n329), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n335), .A2(new_n337), .A3(new_n323), .A4(new_n326), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n334), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(KEYINPUT12), .B1(new_n322), .B2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT12), .ZN(new_n341));
  INV_X1    g155(.A(new_n339), .ZN(new_n342));
  AOI211_X1 g156(.A(new_n341), .B(new_n342), .C1(new_n314), .C2(new_n321), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n312), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(KEYINPUT68), .B1(new_n265), .B2(new_n266), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n263), .A2(new_n264), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n315), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n258), .A2(new_n264), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT68), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n345), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n211), .A2(KEYINPUT4), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n351), .B(new_n232), .C1(new_n352), .C2(new_n296), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT10), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n321), .A2(new_n354), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n211), .A2(KEYINPUT10), .A3(new_n259), .A4(new_n241), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n353), .A2(new_n342), .A3(new_n355), .A4(new_n356), .ZN(new_n357));
  XNOR2_X1  g171(.A(G110), .B(G140), .ZN(new_n358));
  INV_X1    g172(.A(G227), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n359), .A2(G953), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n358), .B(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  AND2_X1   g176(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  AND3_X1   g177(.A1(new_n320), .A2(new_n211), .A3(new_n241), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n259), .B1(new_n211), .B2(new_n241), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n339), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(new_n341), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n322), .A2(KEYINPUT12), .A3(new_n339), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n367), .A2(new_n368), .A3(KEYINPUT82), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n344), .A2(new_n363), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n353), .A2(new_n355), .A3(new_n356), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n339), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n357), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n361), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n370), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G469), .ZN(new_n376));
  INV_X1    g190(.A(G902), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n357), .B1(new_n340), .B2(new_n343), .ZN(new_n379));
  AOI22_X1  g193(.A1(new_n379), .A2(new_n361), .B1(new_n363), .B2(new_n372), .ZN(new_n380));
  OAI21_X1  g194(.A(G469), .B1(new_n380), .B2(G902), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n311), .B1(new_n378), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n308), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G237), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT70), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT70), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G237), .ZN(new_n387));
  AOI21_X1  g201(.A(G953), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n252), .A2(KEYINPUT85), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT85), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G143), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  AND3_X1   g206(.A1(new_n388), .A2(G214), .A3(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n391), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n394), .B1(new_n388), .B2(G214), .ZN(new_n395));
  OAI21_X1  g209(.A(G131), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(KEYINPUT88), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n386), .A2(G237), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n384), .A2(KEYINPUT70), .ZN(new_n399));
  OAI211_X1 g213(.A(G214), .B(new_n269), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n391), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n388), .A2(G214), .A3(new_n392), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT88), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n403), .A2(new_n404), .A3(G131), .ZN(new_n405));
  INV_X1    g219(.A(G131), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n401), .A2(new_n406), .A3(new_n402), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n397), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT75), .ZN(new_n409));
  INV_X1    g223(.A(G140), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(G125), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n260), .A2(G140), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT16), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n409), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(G125), .B(G140), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(KEYINPUT75), .A3(KEYINPUT16), .ZN(new_n417));
  INV_X1    g231(.A(new_n411), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n414), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n415), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n420), .A2(new_n250), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT89), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT19), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n416), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(KEYINPUT89), .A2(KEYINPUT19), .ZN(new_n425));
  MUX2_X1   g239(.A(new_n416), .B(new_n424), .S(new_n425), .Z(new_n426));
  AOI21_X1  g240(.A(new_n421), .B1(new_n426), .B2(new_n250), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n408), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(KEYINPUT18), .A2(G131), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n401), .A2(new_n429), .A3(new_n402), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT87), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n430), .B(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(KEYINPUT76), .B1(new_n413), .B2(G146), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT76), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n416), .A2(new_n434), .A3(new_n250), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT86), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n436), .B(new_n437), .C1(new_n250), .C2(new_n416), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n434), .B1(new_n416), .B2(new_n250), .ZN(new_n439));
  AND4_X1   g253(.A1(new_n434), .A2(new_n411), .A3(new_n412), .A4(new_n250), .ZN(new_n440));
  OAI22_X1  g254(.A1(new_n439), .A2(new_n440), .B1(new_n250), .B2(new_n416), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT86), .ZN(new_n442));
  INV_X1    g256(.A(new_n429), .ZN(new_n443));
  AOI22_X1  g257(.A1(new_n438), .A2(new_n442), .B1(new_n443), .B2(new_n403), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n432), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n428), .A2(new_n445), .ZN(new_n446));
  XNOR2_X1  g260(.A(G113), .B(G122), .ZN(new_n447));
  XNOR2_X1  g261(.A(KEYINPUT90), .B(G104), .ZN(new_n448));
  XOR2_X1   g262(.A(new_n447), .B(new_n448), .Z(new_n449));
  NAND2_X1  g263(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT17), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n397), .A2(new_n451), .A3(new_n405), .A4(new_n407), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n404), .B1(new_n403), .B2(G131), .ZN(new_n453));
  AOI211_X1 g267(.A(KEYINPUT88), .B(new_n406), .C1(new_n401), .C2(new_n402), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT17), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n416), .A2(KEYINPUT16), .ZN(new_n456));
  AOI22_X1  g270(.A1(new_n456), .A2(new_n409), .B1(new_n414), .B2(new_n418), .ZN(new_n457));
  AOI21_X1  g271(.A(G146), .B1(new_n457), .B2(new_n417), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(new_n421), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n452), .A2(new_n455), .A3(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n449), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(new_n461), .A3(new_n445), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n450), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(G475), .A2(G902), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(KEYINPUT20), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT20), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n463), .A2(new_n467), .A3(new_n464), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(G234), .A2(G237), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n470), .A2(G952), .A3(new_n269), .ZN(new_n471));
  XOR2_X1   g285(.A(new_n471), .B(KEYINPUT94), .Z(new_n472));
  AND3_X1   g286(.A1(new_n470), .A2(G902), .A3(G953), .ZN(new_n473));
  XNOR2_X1  g287(.A(KEYINPUT21), .B(G898), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AND2_X1   g289(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n256), .A2(G143), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT91), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT13), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n252), .A2(G128), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n479), .B(new_n480), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n482), .A2(new_n481), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n484), .A2(new_n478), .ZN(new_n485));
  OAI21_X1  g299(.A(KEYINPUT91), .B1(new_n479), .B2(new_n481), .ZN(new_n486));
  OAI211_X1 g300(.A(G134), .B(new_n483), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n216), .A2(G122), .ZN(new_n488));
  INV_X1    g302(.A(G122), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n489), .A2(G116), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n189), .ZN(new_n492));
  OAI21_X1  g306(.A(G107), .B1(new_n488), .B2(new_n490), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n478), .A2(new_n482), .ZN(new_n494));
  AOI22_X1  g308(.A1(new_n492), .A2(new_n493), .B1(new_n325), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n487), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(KEYINPUT92), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT92), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n487), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT93), .ZN(new_n500));
  INV_X1    g314(.A(new_n490), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n500), .B1(new_n501), .B2(KEYINPUT14), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n501), .B1(new_n488), .B2(KEYINPUT14), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NOR3_X1   g318(.A1(new_n501), .A2(new_n500), .A3(KEYINPUT14), .ZN(new_n505));
  OAI21_X1  g319(.A(G107), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n494), .A2(new_n325), .ZN(new_n507));
  OAI21_X1  g321(.A(G134), .B1(new_n478), .B2(new_n482), .ZN(new_n508));
  AOI22_X1  g322(.A1(new_n507), .A2(new_n508), .B1(new_n189), .B2(new_n491), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n497), .A2(new_n499), .A3(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(G217), .ZN(new_n512));
  NOR3_X1   g326(.A1(new_n309), .A2(new_n512), .A3(G953), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  AOI22_X1  g329(.A1(new_n496), .A2(KEYINPUT92), .B1(new_n506), .B2(new_n509), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n516), .A2(new_n499), .A3(new_n513), .ZN(new_n517));
  AOI21_X1  g331(.A(G902), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(G478), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n519), .A2(KEYINPUT15), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n518), .B(new_n520), .ZN(new_n521));
  AND3_X1   g335(.A1(new_n460), .A2(new_n461), .A3(new_n445), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n461), .B1(new_n460), .B2(new_n445), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n377), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(G475), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n469), .A2(new_n477), .A3(new_n521), .A4(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(KEYINPUT95), .B1(new_n383), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(G472), .A2(G902), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT31), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n351), .A2(new_n339), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n254), .B1(G143), .B2(new_n250), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n315), .B1(new_n532), .B2(new_n256), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n336), .A2(new_n326), .ZN(new_n534));
  AOI22_X1  g348(.A1(new_n533), .A2(new_n255), .B1(G131), .B2(new_n534), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n335), .A2(new_n337), .A3(new_n406), .A4(new_n326), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n531), .A2(KEYINPUT30), .A3(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT30), .ZN(new_n539));
  AOI22_X1  g353(.A1(new_n334), .A2(new_n338), .B1(new_n347), .B2(new_n348), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n534), .A2(G131), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n259), .A2(new_n536), .A3(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n539), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n538), .A2(new_n230), .A3(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT69), .ZN(new_n545));
  AND2_X1   g359(.A1(new_n227), .A2(new_n229), .ZN(new_n546));
  AOI22_X1  g360(.A1(new_n351), .A2(new_n339), .B1(new_n535), .B2(new_n536), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n544), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n538), .A2(new_n543), .A3(new_n545), .A4(new_n230), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n552));
  AND3_X1   g366(.A1(new_n388), .A2(G210), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n552), .B1(new_n388), .B2(G210), .ZN(new_n554));
  XNOR2_X1  g368(.A(KEYINPUT26), .B(G101), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  OR3_X1    g370(.A1(new_n553), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n556), .B1(new_n553), .B2(new_n554), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n530), .B1(new_n551), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n559), .ZN(new_n561));
  AOI211_X1 g375(.A(KEYINPUT31), .B(new_n561), .C1(new_n549), .C2(new_n550), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n547), .ZN(new_n564));
  OAI21_X1  g378(.A(KEYINPUT28), .B1(new_n564), .B2(new_n230), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT28), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n546), .A2(new_n547), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n230), .B1(new_n540), .B2(new_n542), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n561), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n529), .B1(new_n563), .B2(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(KEYINPUT72), .B1(new_n572), .B2(KEYINPUT32), .ZN(new_n573));
  INV_X1    g387(.A(G472), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT29), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n568), .A2(new_n575), .A3(new_n569), .ZN(new_n576));
  AOI22_X1  g390(.A1(new_n565), .A2(new_n567), .B1(new_n230), .B2(new_n564), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n576), .B(new_n559), .C1(new_n575), .C2(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n559), .B1(new_n549), .B2(new_n550), .ZN(new_n579));
  AOI21_X1  g393(.A(G902), .B1(new_n579), .B2(new_n575), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n574), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n581), .B1(new_n572), .B2(KEYINPUT32), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n551), .A2(new_n559), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(KEYINPUT31), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n551), .A2(new_n530), .A3(new_n559), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n584), .A2(new_n571), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n528), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT72), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT32), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n573), .A2(new_n582), .A3(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(G234), .ZN(new_n592));
  OAI21_X1  g406(.A(G217), .B1(new_n592), .B2(G902), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(KEYINPUT73), .ZN(new_n594));
  XNOR2_X1  g408(.A(KEYINPUT22), .B(G137), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n269), .A2(G221), .A3(G234), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n595), .B(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n213), .A2(G128), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n256), .A2(KEYINPUT23), .A3(G119), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n256), .A2(G119), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n599), .B(new_n600), .C1(new_n602), .C2(KEYINPUT23), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(G110), .ZN(new_n604));
  XOR2_X1   g418(.A(KEYINPUT24), .B(G110), .Z(new_n605));
  NAND2_X1  g419(.A1(new_n601), .A2(new_n599), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT74), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n601), .A2(new_n599), .A3(KEYINPUT74), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n605), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n436), .B1(new_n604), .B2(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n611), .A2(new_n421), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n603), .A2(G110), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n608), .A2(new_n609), .A3(new_n605), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n457), .A2(G146), .A3(new_n417), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n420), .A2(new_n250), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n598), .B1(new_n612), .B2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n615), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n620), .B1(new_n458), .B2(new_n421), .ZN(new_n621));
  OAI211_X1 g435(.A(new_n616), .B(new_n436), .C1(new_n604), .C2(new_n610), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n621), .A2(new_n622), .A3(new_n597), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n619), .A2(new_n623), .A3(new_n377), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT25), .ZN(new_n625));
  AND2_X1   g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n594), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AND2_X1   g442(.A1(new_n619), .A2(new_n623), .ZN(new_n629));
  AOI21_X1  g443(.A(G902), .B1(new_n592), .B2(G217), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT77), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n467), .B1(new_n463), .B2(new_n464), .ZN(new_n636));
  INV_X1    g450(.A(new_n464), .ZN(new_n637));
  AOI211_X1 g451(.A(KEYINPUT20), .B(new_n637), .C1(new_n450), .C2(new_n462), .ZN(new_n638));
  OAI211_X1 g452(.A(new_n525), .B(new_n521), .C1(new_n636), .C2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n639), .A2(new_n476), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT95), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n640), .A2(new_n641), .A3(new_n308), .A4(new_n382), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n527), .A2(new_n591), .A3(new_n635), .A4(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(KEYINPUT96), .B(G101), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G3));
  AOI211_X1 g459(.A(G469), .B(G902), .C1(new_n370), .C2(new_n374), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n379), .A2(new_n361), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n363), .A2(new_n372), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n647), .A2(G469), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(G469), .A2(G902), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n310), .B1(new_n646), .B2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n634), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(G902), .B1(new_n563), .B2(new_n571), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(new_n574), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n655), .A2(new_n572), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(new_n657), .B(KEYINPUT97), .Z(new_n658));
  NAND2_X1  g472(.A1(new_n377), .A2(G478), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n511), .A2(new_n514), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n513), .B1(new_n516), .B2(new_n499), .ZN(new_n661));
  OAI21_X1  g475(.A(KEYINPUT33), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT33), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n515), .A2(new_n663), .A3(new_n517), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n659), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(KEYINPUT98), .B1(new_n518), .B2(G478), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AOI211_X1 g481(.A(KEYINPUT98), .B(new_n659), .C1(new_n662), .C2(new_n664), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n525), .B1(new_n636), .B2(new_n638), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n188), .B1(new_n301), .B2(new_n302), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n277), .A2(new_n300), .A3(new_n303), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n671), .A2(new_n674), .A3(new_n476), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n658), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT34), .B(G104), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G6));
  INV_X1    g492(.A(new_n520), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n518), .B(new_n679), .ZN(new_n680));
  OAI211_X1 g494(.A(new_n525), .B(new_n680), .C1(new_n636), .C2(new_n638), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n674), .A2(new_n476), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n658), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT35), .B(G107), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G9));
  OR3_X1    g499(.A1(new_n612), .A2(new_n618), .A3(KEYINPUT99), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n598), .A2(KEYINPUT36), .ZN(new_n687));
  OAI21_X1  g501(.A(KEYINPUT99), .B1(new_n612), .B2(new_n618), .ZN(new_n688));
  AND3_X1   g502(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n687), .B1(new_n686), .B2(new_n688), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n630), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n628), .A2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n655), .A2(new_n572), .A3(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n527), .A2(new_n694), .A3(new_n642), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT37), .B(G110), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT100), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n695), .B(new_n697), .ZN(G12));
  NOR3_X1   g512(.A1(new_n652), .A2(new_n674), .A3(new_n693), .ZN(new_n699));
  XOR2_X1   g513(.A(new_n472), .B(KEYINPUT102), .Z(new_n700));
  INV_X1    g514(.A(G900), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n473), .A2(new_n701), .ZN(new_n702));
  XOR2_X1   g516(.A(new_n702), .B(KEYINPUT101), .Z(new_n703));
  NAND2_X1  g517(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n681), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n591), .A2(new_n699), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G128), .ZN(G30));
  XNOR2_X1  g522(.A(new_n704), .B(KEYINPUT39), .ZN(new_n709));
  AND2_X1   g523(.A1(new_n382), .A2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT40), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n307), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n304), .B1(new_n277), .B2(new_n300), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(KEYINPUT38), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n670), .A2(new_n693), .A3(new_n680), .A4(new_n187), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n712), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n710), .A2(new_n711), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n549), .A2(new_n559), .A3(new_n550), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n559), .B1(new_n546), .B2(new_n547), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n564), .A2(new_n230), .ZN(new_n722));
  AOI21_X1  g536(.A(G902), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n574), .B1(new_n720), .B2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(KEYINPUT103), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n725), .B1(KEYINPUT32), .B2(new_n572), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT104), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n726), .A2(new_n573), .A3(new_n727), .A4(new_n590), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n588), .B1(new_n587), .B2(new_n589), .ZN(new_n730));
  AOI211_X1 g544(.A(KEYINPUT72), .B(KEYINPUT32), .C1(new_n586), .C2(new_n528), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n727), .B1(new_n732), .B2(new_n726), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n718), .B(new_n719), .C1(new_n729), .C2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G143), .ZN(G45));
  NAND3_X1  g549(.A1(new_n669), .A2(new_n670), .A3(new_n704), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n591), .A2(new_n699), .A3(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G146), .ZN(G48));
  INV_X1    g553(.A(new_n375), .ZN(new_n740));
  OAI21_X1  g554(.A(G469), .B1(new_n740), .B2(G902), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n741), .A2(new_n310), .A3(new_n378), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n591), .A2(new_n675), .A3(new_n635), .A4(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(KEYINPUT41), .B(G113), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G15));
  NAND4_X1  g560(.A1(new_n591), .A2(new_n682), .A3(new_n635), .A4(new_n743), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G116), .ZN(G18));
  NOR3_X1   g562(.A1(new_n742), .A2(new_n674), .A3(new_n693), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n749), .A2(new_n591), .A3(new_n640), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G119), .ZN(G21));
  NAND4_X1  g565(.A1(new_n670), .A2(new_n672), .A3(new_n680), .A4(new_n673), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n752), .A2(new_n742), .A3(new_n476), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT105), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n754), .B1(new_n654), .B2(new_n574), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n586), .A2(new_n377), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n756), .A2(KEYINPUT105), .A3(G472), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n563), .B1(new_n559), .B2(new_n577), .ZN(new_n758));
  AOI22_X1  g572(.A1(new_n755), .A2(new_n757), .B1(new_n528), .B2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(new_n632), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n753), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G122), .ZN(G24));
  NAND3_X1  g576(.A1(new_n749), .A2(new_n759), .A3(new_n737), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G125), .ZN(G27));
  NAND3_X1  g578(.A1(new_n306), .A2(new_n187), .A3(new_n307), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n736), .A2(new_n652), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n587), .A2(new_n589), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n632), .B1(new_n582), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n766), .A2(new_n768), .A3(KEYINPUT42), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n766), .A2(new_n591), .A3(new_n635), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT42), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n770), .A2(KEYINPUT106), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g586(.A(KEYINPUT106), .B1(new_n770), .B2(new_n771), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n769), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G131), .ZN(G33));
  NAND2_X1  g589(.A1(new_n591), .A2(new_n635), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n652), .A2(new_n765), .ZN(new_n777));
  AOI22_X1  g591(.A1(new_n466), .A2(new_n468), .B1(G475), .B2(new_n524), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT107), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n778), .A2(new_n779), .A3(new_n680), .A4(new_n704), .ZN(new_n780));
  OAI21_X1  g594(.A(KEYINPUT107), .B1(new_n681), .B2(new_n705), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n777), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  OAI21_X1  g596(.A(KEYINPUT108), .B1(new_n776), .B2(new_n782), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n777), .A2(new_n780), .A3(new_n781), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT108), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n784), .A2(new_n785), .A3(new_n591), .A4(new_n635), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G134), .ZN(G36));
  INV_X1    g602(.A(KEYINPUT98), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n665), .A2(new_n789), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n790), .B1(new_n665), .B2(new_n666), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n670), .A2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT43), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g608(.A(KEYINPUT43), .B1(new_n670), .B2(new_n791), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n796), .A2(new_n656), .A3(new_n693), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(KEYINPUT44), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(KEYINPUT109), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n797), .A2(KEYINPUT44), .ZN(new_n800));
  INV_X1    g614(.A(new_n765), .ZN(new_n801));
  OR2_X1    g615(.A1(new_n380), .A2(KEYINPUT45), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n380), .A2(KEYINPUT45), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n802), .A2(G469), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT46), .B1(new_n804), .B2(new_n650), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n805), .A2(new_n646), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n804), .A2(KEYINPUT46), .A3(new_n650), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n311), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n808), .A2(new_n709), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n800), .A2(new_n801), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n799), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G137), .ZN(G39));
  NAND2_X1  g626(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n808), .A2(new_n813), .ZN(new_n814));
  XOR2_X1   g628(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n815));
  OAI21_X1  g629(.A(new_n814), .B1(new_n808), .B2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  NOR4_X1   g631(.A1(new_n591), .A2(new_n635), .A3(new_n736), .A4(new_n765), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(G140), .ZN(G42));
  NOR3_X1   g634(.A1(new_n632), .A2(new_n188), .A3(new_n311), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n716), .A2(new_n792), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n741), .A2(new_n378), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n822), .B1(KEYINPUT49), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n733), .A2(new_n729), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n823), .A2(KEYINPUT49), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(KEYINPUT111), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n824), .A2(new_n825), .A3(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT53), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n308), .A2(new_n477), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n671), .A2(new_n681), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n653), .A2(new_n831), .A3(new_n656), .A4(new_n832), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n643), .A2(new_n695), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n758), .A2(new_n528), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT105), .B1(new_n756), .B2(G472), .ZN(new_n836));
  AOI211_X1 g650(.A(new_n754), .B(new_n574), .C1(new_n586), .C2(new_n377), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n692), .B(new_n835), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n737), .A2(new_n777), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT112), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n573), .A2(new_n582), .A3(new_n590), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n639), .A2(new_n693), .A3(new_n705), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n777), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n841), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n591), .A2(KEYINPUT112), .A3(new_n843), .A4(new_n777), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n840), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n834), .A2(new_n787), .A3(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT113), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n829), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n692), .A2(new_n705), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n382), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n852), .A2(new_n752), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n853), .B1(new_n733), .B2(new_n729), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT52), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n591), .B(new_n699), .C1(new_n706), .C2(new_n737), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n854), .A2(new_n855), .A3(new_n763), .A4(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n763), .ZN(new_n858));
  INV_X1    g672(.A(new_n853), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n572), .A2(KEYINPUT32), .ZN(new_n860));
  INV_X1    g674(.A(new_n725), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n573), .A2(new_n590), .A3(new_n860), .A4(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(KEYINPUT104), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n859), .B1(new_n863), .B2(new_n728), .ZN(new_n864));
  OAI21_X1  g678(.A(KEYINPUT52), .B1(new_n858), .B2(new_n864), .ZN(new_n865));
  AND4_X1   g679(.A1(new_n744), .A2(new_n761), .A3(new_n747), .A4(new_n750), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n857), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n834), .A2(new_n787), .A3(new_n847), .A4(KEYINPUT113), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n850), .A2(new_n867), .A3(new_n774), .A4(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT54), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n774), .A2(new_n857), .A3(new_n866), .A4(new_n865), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n829), .B1(new_n871), .B2(new_n848), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n869), .A2(new_n870), .A3(new_n872), .ZN(new_n873));
  OR3_X1    g687(.A1(new_n871), .A2(new_n829), .A3(new_n848), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(new_n872), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n873), .B1(new_n875), .B2(KEYINPUT54), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n796), .A2(new_n700), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n743), .A2(KEYINPUT117), .A3(new_n801), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT117), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n879), .B1(new_n742), .B2(new_n765), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n877), .A2(new_n881), .A3(new_n768), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT121), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(KEYINPUT48), .ZN(new_n884));
  OR2_X1    g698(.A1(new_n883), .A2(KEYINPUT48), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n882), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  AOI211_X1 g700(.A(new_n634), .B(new_n472), .C1(new_n878), .C2(new_n880), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(new_n825), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n886), .B1(new_n888), .B2(new_n671), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n882), .A2(new_n884), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n877), .A2(new_n760), .A3(new_n759), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n891), .A2(new_n674), .A3(new_n742), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n269), .A2(G952), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT120), .ZN(new_n894));
  NOR4_X1   g708(.A1(new_n889), .A2(new_n890), .A3(new_n892), .A4(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT116), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n716), .A2(new_n188), .A3(new_n743), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n896), .B1(new_n891), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(KEYINPUT50), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT50), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n896), .B(new_n900), .C1(new_n891), .C2(new_n897), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n877), .A2(new_n881), .A3(new_n692), .A4(new_n759), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n887), .A2(new_n825), .A3(new_n778), .A4(new_n791), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT118), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n904), .A2(new_n905), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n902), .B(new_n903), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n741), .A2(new_n311), .A3(new_n378), .ZN(new_n909));
  INV_X1    g723(.A(new_n814), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n808), .A2(new_n815), .ZN(new_n911));
  OAI211_X1 g725(.A(KEYINPUT119), .B(new_n909), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n891), .A2(new_n765), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(KEYINPUT119), .B1(new_n816), .B2(new_n909), .ZN(new_n915));
  OAI21_X1  g729(.A(KEYINPUT51), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n895), .B1(new_n908), .B2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT51), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n909), .B(KEYINPUT115), .Z(new_n919));
  INV_X1    g733(.A(KEYINPUT114), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n919), .B1(new_n817), .B2(new_n920), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n816), .A2(KEYINPUT114), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n913), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OR2_X1    g737(.A1(new_n906), .A2(new_n907), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n923), .A2(new_n924), .A3(new_n902), .A4(new_n903), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n917), .B1(new_n918), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n876), .A2(KEYINPUT122), .A3(new_n926), .ZN(new_n927));
  OR2_X1    g741(.A1(G952), .A2(G953), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(KEYINPUT122), .B1(new_n876), .B2(new_n926), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n828), .B1(new_n929), .B2(new_n930), .ZN(G75));
  AOI21_X1  g745(.A(new_n377), .B1(new_n869), .B2(new_n872), .ZN(new_n932));
  AOI21_X1  g746(.A(KEYINPUT56), .B1(new_n932), .B2(G210), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n249), .A2(new_n276), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(new_n274), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT55), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n933), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n269), .A2(G952), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  OR3_X1    g755(.A1(new_n933), .A2(KEYINPUT123), .A3(new_n937), .ZN(new_n942));
  OAI21_X1  g756(.A(KEYINPUT123), .B1(new_n933), .B2(new_n937), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(G51));
  AOI211_X1 g758(.A(new_n377), .B(new_n804), .C1(new_n869), .C2(new_n872), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n650), .B(KEYINPUT57), .Z(new_n946));
  AOI21_X1  g760(.A(new_n870), .B1(new_n869), .B2(new_n872), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n946), .B1(new_n873), .B2(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n945), .B1(new_n948), .B2(new_n375), .ZN(new_n949));
  OAI21_X1  g763(.A(KEYINPUT124), .B1(new_n949), .B2(new_n939), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT124), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n869), .A2(new_n872), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(KEYINPUT54), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n869), .A2(new_n870), .A3(new_n872), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n740), .B1(new_n955), .B2(new_n946), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n951), .B(new_n940), .C1(new_n956), .C2(new_n945), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n950), .A2(new_n957), .ZN(G54));
  AND2_X1   g772(.A1(KEYINPUT58), .A2(G475), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n932), .A2(new_n463), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n463), .B1(new_n932), .B2(new_n959), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n960), .A2(new_n961), .A3(new_n939), .ZN(G60));
  NAND2_X1  g776(.A1(new_n662), .A2(new_n664), .ZN(new_n963));
  INV_X1    g777(.A(new_n876), .ZN(new_n964));
  NAND2_X1  g778(.A1(G478), .A2(G902), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT59), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n963), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n955), .A2(new_n963), .A3(new_n966), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n940), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n967), .A2(new_n969), .ZN(G63));
  XNOR2_X1  g784(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n971));
  NAND2_X1  g785(.A1(G217), .A2(G902), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n971), .B(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n973), .B1(new_n869), .B2(new_n872), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n974), .B1(new_n689), .B2(new_n690), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n975), .B(new_n940), .C1(new_n629), .C2(new_n974), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT61), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n976), .B(new_n977), .ZN(G66));
  AND2_X1   g792(.A1(new_n866), .A2(new_n834), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(G224), .A2(G953), .ZN(new_n981));
  OAI22_X1  g795(.A1(new_n980), .A2(G953), .B1(new_n474), .B2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(G898), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n934), .B1(new_n983), .B2(G953), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n982), .B(new_n984), .ZN(G69));
  AOI22_X1  g799(.A1(new_n799), .A2(new_n810), .B1(new_n817), .B2(new_n818), .ZN(new_n986));
  INV_X1    g800(.A(new_n776), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n987), .A2(new_n710), .A3(new_n801), .A4(new_n832), .ZN(new_n988));
  INV_X1    g802(.A(new_n858), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n734), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(KEYINPUT62), .ZN(new_n991));
  OR2_X1    g805(.A1(new_n990), .A2(KEYINPUT62), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n986), .A2(new_n988), .A3(new_n991), .A4(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(new_n269), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n538), .A2(new_n543), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(new_n426), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n269), .A2(G900), .ZN(new_n998));
  INV_X1    g812(.A(new_n752), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n809), .A2(new_n999), .A3(new_n768), .ZN(new_n1000));
  AND3_X1   g814(.A1(new_n1000), .A2(new_n787), .A3(new_n989), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n986), .A2(new_n774), .A3(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n998), .B1(new_n1002), .B2(new_n269), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n997), .B1(new_n1003), .B2(new_n996), .ZN(new_n1004));
  OAI21_X1  g818(.A(G953), .B1(new_n359), .B2(new_n701), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1005), .B(KEYINPUT126), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1004), .B(new_n1006), .ZN(G72));
  NAND2_X1  g821(.A1(G472), .A2(G902), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1008), .B(KEYINPUT63), .Z(new_n1009));
  OAI21_X1  g823(.A(new_n1009), .B1(new_n993), .B2(new_n980), .ZN(new_n1010));
  INV_X1    g824(.A(new_n720), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n939), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(new_n579), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n875), .A2(new_n1013), .A3(new_n720), .A4(new_n1009), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1009), .B1(new_n1002), .B2(new_n980), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1015), .A2(new_n579), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n1012), .A2(new_n1014), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT127), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND4_X1  g833(.A1(new_n1012), .A2(KEYINPUT127), .A3(new_n1014), .A4(new_n1016), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1019), .A2(new_n1020), .ZN(G57));
endmodule


