

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753;

  XNOR2_X1 U378 ( .A(n519), .B(n441), .ZN(n729) );
  XNOR2_X1 U379 ( .A(n425), .B(n424), .ZN(n519) );
  INV_X1 U380 ( .A(KEYINPUT3), .ZN(n439) );
  NAND2_X1 U381 ( .A1(n718), .A2(G475), .ZN(n645) );
  AND2_X2 U382 ( .A1(n372), .A2(n374), .ZN(n718) );
  AND2_X2 U383 ( .A1(n557), .A2(n676), .ZN(n533) );
  XNOR2_X1 U384 ( .A(n571), .B(n570), .ZN(n619) );
  NAND2_X2 U385 ( .A1(n544), .A2(n543), .ZN(n561) );
  XNOR2_X2 U386 ( .A(n527), .B(G472), .ZN(n681) );
  NOR2_X1 U387 ( .A1(n553), .A2(n552), .ZN(n661) );
  INV_X2 U388 ( .A(G953), .ZN(n741) );
  XNOR2_X1 U389 ( .A(n409), .B(n365), .ZN(n543) );
  NOR2_X2 U390 ( .A1(G953), .A2(G237), .ZN(n516) );
  INV_X1 U391 ( .A(KEYINPUT110), .ZN(n398) );
  XNOR2_X1 U392 ( .A(n396), .B(KEYINPUT119), .ZN(n748) );
  XNOR2_X1 U393 ( .A(n405), .B(n356), .ZN(n417) );
  NOR2_X1 U394 ( .A1(n705), .A2(n548), .ZN(n541) );
  XNOR2_X1 U395 ( .A(n399), .B(n398), .ZN(n607) );
  XNOR2_X1 U396 ( .A(n539), .B(n538), .ZN(n705) );
  XNOR2_X1 U397 ( .A(n358), .B(G478), .ZN(n550) );
  XNOR2_X1 U398 ( .A(n481), .B(G134), .ZN(n508) );
  XOR2_X1 U399 ( .A(KEYINPUT70), .B(G131), .Z(n509) );
  NOR2_X2 U400 ( .A1(n603), .A2(n620), .ZN(n694) );
  XNOR2_X1 U401 ( .A(n736), .B(G146), .ZN(n525) );
  XNOR2_X1 U402 ( .A(n442), .B(G146), .ZN(n467) );
  INV_X1 U403 ( .A(G125), .ZN(n442) );
  XOR2_X1 U404 ( .A(G137), .B(G140), .Z(n511) );
  XNOR2_X1 U405 ( .A(n508), .B(n509), .ZN(n736) );
  OR2_X1 U406 ( .A1(n713), .A2(G902), .ZN(n515) );
  NOR2_X1 U407 ( .A1(n611), .A2(n610), .ZN(n613) );
  INV_X1 U408 ( .A(KEYINPUT90), .ZN(n427) );
  XNOR2_X1 U409 ( .A(G113), .B(G104), .ZN(n384) );
  XNOR2_X1 U410 ( .A(G140), .B(KEYINPUT101), .ZN(n468) );
  XOR2_X1 U411 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n474) );
  XNOR2_X1 U412 ( .A(n467), .B(n387), .ZN(n498) );
  XNOR2_X1 U413 ( .A(n466), .B(KEYINPUT10), .ZN(n387) );
  AND2_X1 U414 ( .A1(n526), .A2(n630), .ZN(n527) );
  XNOR2_X1 U415 ( .A(G119), .B(G116), .ZN(n424) );
  XNOR2_X1 U416 ( .A(n439), .B(G113), .ZN(n425) );
  XOR2_X1 U417 ( .A(G137), .B(KEYINPUT5), .Z(n518) );
  XNOR2_X1 U418 ( .A(G119), .B(G128), .ZN(n499) );
  XOR2_X1 U419 ( .A(KEYINPUT71), .B(G110), .Z(n500) );
  XNOR2_X1 U420 ( .A(KEYINPUT96), .B(KEYINPUT78), .ZN(n502) );
  XOR2_X1 U421 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n503) );
  XNOR2_X1 U422 ( .A(n486), .B(n485), .ZN(n504) );
  XOR2_X1 U423 ( .A(KEYINPUT68), .B(KEYINPUT8), .Z(n486) );
  NAND2_X1 U424 ( .A1(n391), .A2(KEYINPUT36), .ZN(n390) );
  NAND2_X1 U425 ( .A1(n608), .A2(n395), .ZN(n393) );
  INV_X1 U426 ( .A(n608), .ZN(n391) );
  NAND2_X1 U427 ( .A1(n430), .A2(n357), .ZN(n465) );
  XNOR2_X1 U428 ( .A(n507), .B(KEYINPUT25), .ZN(n420) );
  OR2_X1 U429 ( .A1(n719), .A2(G902), .ZN(n421) );
  INV_X1 U430 ( .A(KEYINPUT64), .ZN(n373) );
  XNOR2_X1 U431 ( .A(n411), .B(n512), .ZN(n514) );
  XNOR2_X1 U432 ( .A(n359), .B(n513), .ZN(n411) );
  XOR2_X1 U433 ( .A(KEYINPUT12), .B(KEYINPUT102), .Z(n471) );
  XOR2_X1 U434 ( .A(KEYINPUT11), .B(KEYINPUT98), .Z(n469) );
  INV_X1 U435 ( .A(G237), .ZN(n451) );
  NOR2_X1 U436 ( .A1(n675), .A2(n576), .ZN(n606) );
  NAND2_X1 U437 ( .A1(n676), .A2(n360), .ZN(n576) );
  NOR2_X1 U438 ( .A1(n622), .A2(n621), .ZN(n627) );
  INV_X1 U439 ( .A(KEYINPUT48), .ZN(n612) );
  XNOR2_X1 U440 ( .A(n562), .B(KEYINPUT45), .ZN(n626) );
  XNOR2_X1 U441 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n444) );
  NAND2_X1 U442 ( .A1(n626), .A2(n627), .ZN(n667) );
  AND2_X1 U443 ( .A1(n606), .A2(n659), .ZN(n400) );
  OR2_X1 U444 ( .A1(n681), .A2(n435), .ZN(n419) );
  XNOR2_X1 U445 ( .A(n567), .B(KEYINPUT113), .ZN(n418) );
  NOR2_X1 U446 ( .A1(n676), .A2(n407), .ZN(n406) );
  NAND2_X1 U447 ( .A1(n408), .A2(n360), .ZN(n407) );
  INV_X1 U448 ( .A(KEYINPUT76), .ZN(n382) );
  XNOR2_X1 U449 ( .A(n446), .B(G107), .ZN(n728) );
  XOR2_X1 U450 ( .A(KEYINPUT105), .B(G122), .Z(n483) );
  XNOR2_X1 U451 ( .A(G116), .B(G107), .ZN(n482) );
  XNOR2_X1 U452 ( .A(KEYINPUT103), .B(KEYINPUT9), .ZN(n487) );
  XOR2_X1 U453 ( .A(KEYINPUT104), .B(KEYINPUT7), .Z(n488) );
  XNOR2_X1 U454 ( .A(n509), .B(n384), .ZN(n388) );
  XNOR2_X1 U455 ( .A(n728), .B(n521), .ZN(n512) );
  NAND2_X1 U456 ( .A1(G234), .A2(G237), .ZN(n460) );
  NAND2_X1 U457 ( .A1(n535), .A2(n412), .ZN(n539) );
  INV_X1 U458 ( .A(KEYINPUT91), .ZN(n536) );
  INV_X1 U459 ( .A(n681), .ZN(n577) );
  XNOR2_X1 U460 ( .A(n385), .B(KEYINPUT22), .ZN(n557) );
  NOR2_X1 U461 ( .A1(n548), .A2(n497), .ZN(n385) );
  XNOR2_X1 U462 ( .A(n524), .B(n525), .ZN(n630) );
  XNOR2_X1 U463 ( .A(n402), .B(n735), .ZN(n719) );
  AND2_X1 U464 ( .A1(n504), .A2(G221), .ZN(n403) );
  NAND2_X1 U465 ( .A1(n619), .A2(n603), .ZN(n405) );
  OR2_X1 U466 ( .A1(n614), .A2(n390), .ZN(n389) );
  NOR2_X1 U467 ( .A1(n587), .A2(n586), .ZN(n657) );
  XNOR2_X1 U468 ( .A(n603), .B(n401), .ZN(n659) );
  INV_X1 U469 ( .A(KEYINPUT109), .ZN(n401) );
  XNOR2_X1 U470 ( .A(n712), .B(n371), .ZN(n714) );
  XNOR2_X1 U471 ( .A(n713), .B(n711), .ZN(n371) );
  AND2_X1 U472 ( .A1(n709), .A2(n708), .ZN(n710) );
  XOR2_X1 U473 ( .A(n572), .B(KEYINPUT40), .Z(n356) );
  INV_X1 U474 ( .A(n675), .ZN(n408) );
  AND2_X1 U475 ( .A1(n432), .A2(n434), .ZN(n357) );
  OR2_X1 U476 ( .A1(G902), .A2(n715), .ZN(n358) );
  XOR2_X1 U477 ( .A(n511), .B(n510), .Z(n359) );
  XOR2_X1 U478 ( .A(KEYINPUT82), .B(n565), .Z(n360) );
  INV_X1 U479 ( .A(n689), .ZN(n435) );
  XOR2_X1 U480 ( .A(G143), .B(G122), .Z(n361) );
  XOR2_X1 U481 ( .A(n419), .B(n418), .Z(n362) );
  OR2_X1 U482 ( .A1(n561), .A2(KEYINPUT44), .ZN(n363) );
  AND2_X1 U483 ( .A1(n564), .A2(n464), .ZN(n364) );
  XOR2_X1 U484 ( .A(KEYINPUT80), .B(KEYINPUT35), .Z(n365) );
  XOR2_X1 U485 ( .A(n641), .B(n640), .Z(n366) );
  XOR2_X1 U486 ( .A(n644), .B(n643), .Z(n367) );
  XNOR2_X1 U487 ( .A(n630), .B(KEYINPUT62), .ZN(n368) );
  XNOR2_X1 U488 ( .A(n498), .B(n511), .ZN(n735) );
  XNOR2_X1 U489 ( .A(n634), .B(n633), .ZN(n722) );
  INV_X1 U490 ( .A(n722), .ZN(n380) );
  XOR2_X1 U491 ( .A(KEYINPUT88), .B(KEYINPUT56), .Z(n369) );
  XOR2_X1 U492 ( .A(KEYINPUT66), .B(KEYINPUT60), .Z(n370) );
  NAND2_X1 U493 ( .A1(n426), .A2(n363), .ZN(n562) );
  NOR2_X2 U494 ( .A1(n551), .A2(n550), .ZN(n603) );
  XNOR2_X1 U495 ( .A(n625), .B(n373), .ZN(n372) );
  INV_X1 U496 ( .A(n672), .ZN(n374) );
  XNOR2_X1 U497 ( .A(n375), .B(n369), .ZN(G51) );
  NAND2_X1 U498 ( .A1(n378), .A2(n380), .ZN(n375) );
  XNOR2_X1 U499 ( .A(n376), .B(n370), .ZN(G60) );
  NAND2_X1 U500 ( .A1(n379), .A2(n380), .ZN(n376) );
  XNOR2_X1 U501 ( .A(n377), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U502 ( .A1(n381), .A2(n380), .ZN(n377) );
  NAND2_X1 U503 ( .A1(n417), .A2(n585), .ZN(n416) );
  NOR2_X1 U504 ( .A1(n704), .A2(n587), .ZN(n584) );
  NAND2_X1 U505 ( .A1(n400), .A2(n605), .ZN(n399) );
  XNOR2_X1 U506 ( .A(n428), .B(n427), .ZN(n426) );
  XNOR2_X1 U507 ( .A(n642), .B(n366), .ZN(n378) );
  XNOR2_X1 U508 ( .A(n645), .B(n367), .ZN(n379) );
  XNOR2_X1 U509 ( .A(n631), .B(n368), .ZN(n381) );
  XNOR2_X1 U510 ( .A(n383), .B(n382), .ZN(n568) );
  NAND2_X1 U511 ( .A1(n406), .A2(n580), .ZN(n383) );
  NAND2_X1 U512 ( .A1(n429), .A2(n560), .ZN(n428) );
  NAND2_X1 U513 ( .A1(n386), .A2(n657), .ZN(n599) );
  NAND2_X1 U514 ( .A1(n595), .A2(n594), .ZN(n386) );
  AND2_X1 U515 ( .A1(n600), .A2(n438), .ZN(n601) );
  XNOR2_X1 U516 ( .A(n501), .B(n505), .ZN(n404) );
  XNOR2_X1 U517 ( .A(n404), .B(n403), .ZN(n402) );
  XNOR2_X1 U518 ( .A(n388), .B(n498), .ZN(n478) );
  NAND2_X1 U519 ( .A1(n392), .A2(n389), .ZN(n397) );
  AND2_X1 U520 ( .A1(n394), .A2(n393), .ZN(n392) );
  NAND2_X1 U521 ( .A1(n614), .A2(n395), .ZN(n394) );
  INV_X1 U522 ( .A(KEYINPUT36), .ZN(n395) );
  NAND2_X1 U523 ( .A1(n397), .A2(n535), .ZN(n396) );
  INV_X1 U524 ( .A(n417), .ZN(n750) );
  NAND2_X1 U525 ( .A1(n678), .A2(n580), .ZN(n566) );
  NOR2_X1 U526 ( .A1(n676), .A2(n675), .ZN(n678) );
  XNOR2_X2 U527 ( .A(n421), .B(n420), .ZN(n676) );
  INV_X1 U528 ( .A(n543), .ZN(n753) );
  NAND2_X1 U529 ( .A1(n410), .A2(n597), .ZN(n409) );
  XNOR2_X1 U530 ( .A(n541), .B(n540), .ZN(n410) );
  NOR2_X1 U531 ( .A1(n604), .A2(n413), .ZN(n412) );
  NAND2_X1 U532 ( .A1(n535), .A2(n678), .ZN(n414) );
  INV_X1 U533 ( .A(n678), .ZN(n413) );
  NOR2_X1 U534 ( .A1(n414), .A2(n681), .ZN(n685) );
  XNOR2_X2 U535 ( .A(n580), .B(KEYINPUT1), .ZN(n535) );
  XNOR2_X1 U536 ( .A(n416), .B(n415), .ZN(n602) );
  INV_X1 U537 ( .A(KEYINPUT46), .ZN(n415) );
  XNOR2_X1 U538 ( .A(n729), .B(n422), .ZN(n448) );
  XNOR2_X1 U539 ( .A(n445), .B(n423), .ZN(n422) );
  XNOR2_X1 U540 ( .A(n467), .B(n481), .ZN(n423) );
  NAND2_X1 U541 ( .A1(n561), .A2(KEYINPUT44), .ZN(n429) );
  OR2_X2 U542 ( .A1(n616), .A2(n431), .ZN(n436) );
  XNOR2_X2 U543 ( .A(n455), .B(n454), .ZN(n616) );
  NAND2_X1 U544 ( .A1(n357), .A2(n436), .ZN(n586) );
  AND2_X2 U545 ( .A1(n436), .A2(n364), .ZN(n430) );
  INV_X1 U546 ( .A(n459), .ZN(n431) );
  NAND2_X1 U547 ( .A1(n616), .A2(n433), .ZN(n432) );
  NOR2_X1 U548 ( .A1(n459), .A2(n435), .ZN(n433) );
  NAND2_X1 U549 ( .A1(n435), .A2(n459), .ZN(n434) );
  XNOR2_X1 U550 ( .A(n569), .B(KEYINPUT75), .ZN(n596) );
  AND2_X2 U551 ( .A1(n638), .A2(n636), .ZN(n544) );
  XNOR2_X2 U552 ( .A(n530), .B(n529), .ZN(n638) );
  XNOR2_X2 U553 ( .A(n534), .B(KEYINPUT32), .ZN(n636) );
  BUF_X1 U554 ( .A(n627), .Z(n739) );
  BUF_X1 U555 ( .A(n626), .Z(n723) );
  NAND2_X1 U556 ( .A1(n602), .A2(n601), .ZN(n611) );
  NOR2_X2 U557 ( .A1(n629), .A2(n628), .ZN(n672) );
  OR2_X1 U558 ( .A1(G953), .A2(n706), .ZN(n437) );
  AND2_X1 U559 ( .A1(n599), .A2(n639), .ZN(n438) );
  INV_X1 U560 ( .A(n751), .ZN(n585) );
  INV_X1 U561 ( .A(n604), .ZN(n605) );
  INV_X1 U562 ( .A(KEYINPUT89), .ZN(n609) );
  INV_X1 U563 ( .A(n521), .ZN(n522) );
  XNOR2_X1 U564 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U565 ( .A(n523), .B(n522), .ZN(n524) );
  NAND2_X1 U566 ( .A1(n596), .A2(n690), .ZN(n571) );
  NOR2_X1 U567 ( .A1(n707), .A2(n437), .ZN(n708) );
  XNOR2_X1 U568 ( .A(KEYINPUT16), .B(G122), .ZN(n440) );
  XNOR2_X1 U569 ( .A(n440), .B(KEYINPUT74), .ZN(n441) );
  XNOR2_X2 U570 ( .A(G143), .B(G128), .ZN(n481) );
  NAND2_X1 U571 ( .A1(n741), .A2(G224), .ZN(n443) );
  XNOR2_X1 U572 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U573 ( .A(G110), .B(G104), .Z(n446) );
  XNOR2_X1 U574 ( .A(G101), .B(KEYINPUT67), .ZN(n447) );
  XNOR2_X1 U575 ( .A(n447), .B(KEYINPUT4), .ZN(n521) );
  XNOR2_X1 U576 ( .A(n448), .B(n512), .ZN(n641) );
  XNOR2_X1 U577 ( .A(G902), .B(KEYINPUT93), .ZN(n450) );
  INV_X1 U578 ( .A(KEYINPUT15), .ZN(n449) );
  XNOR2_X1 U579 ( .A(n450), .B(n449), .ZN(n493) );
  INV_X1 U580 ( .A(n493), .ZN(n623) );
  OR2_X2 U581 ( .A1(n641), .A2(n623), .ZN(n455) );
  INV_X1 U582 ( .A(G902), .ZN(n526) );
  NAND2_X1 U583 ( .A1(n526), .A2(n451), .ZN(n456) );
  NAND2_X1 U584 ( .A1(n456), .A2(G210), .ZN(n453) );
  INV_X1 U585 ( .A(KEYINPUT94), .ZN(n452) );
  XNOR2_X1 U586 ( .A(n453), .B(n452), .ZN(n454) );
  NAND2_X1 U587 ( .A1(n456), .A2(G214), .ZN(n689) );
  XNOR2_X1 U588 ( .A(KEYINPUT77), .B(KEYINPUT19), .ZN(n458) );
  INV_X1 U589 ( .A(KEYINPUT65), .ZN(n457) );
  XNOR2_X1 U590 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U591 ( .A(n460), .B(KEYINPUT14), .ZN(n701) );
  INV_X1 U592 ( .A(G952), .ZN(n632) );
  NAND2_X1 U593 ( .A1(n741), .A2(n632), .ZN(n462) );
  NAND2_X1 U594 ( .A1(G953), .A2(n526), .ZN(n461) );
  AND2_X1 U595 ( .A1(n462), .A2(n461), .ZN(n463) );
  AND2_X1 U596 ( .A1(n701), .A2(n463), .ZN(n564) );
  NAND2_X1 U597 ( .A1(G953), .A2(G898), .ZN(n464) );
  XNOR2_X2 U598 ( .A(n465), .B(KEYINPUT0), .ZN(n548) );
  INV_X1 U599 ( .A(KEYINPUT69), .ZN(n466) );
  XNOR2_X1 U600 ( .A(n469), .B(n468), .ZN(n473) );
  NAND2_X1 U601 ( .A1(G214), .A2(n516), .ZN(n470) );
  XNOR2_X1 U602 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U603 ( .A(n473), .B(n472), .ZN(n476) );
  XNOR2_X1 U604 ( .A(n474), .B(n361), .ZN(n475) );
  XNOR2_X1 U605 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U606 ( .A(n478), .B(n477), .ZN(n644) );
  NAND2_X1 U607 ( .A1(n644), .A2(n526), .ZN(n480) );
  XNOR2_X1 U608 ( .A(KEYINPUT13), .B(G475), .ZN(n479) );
  XNOR2_X1 U609 ( .A(n480), .B(n479), .ZN(n551) );
  XNOR2_X1 U610 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U611 ( .A(n508), .B(n484), .ZN(n492) );
  NAND2_X1 U612 ( .A1(G234), .A2(n741), .ZN(n485) );
  NAND2_X1 U613 ( .A1(G217), .A2(n504), .ZN(n490) );
  XNOR2_X1 U614 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U615 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U616 ( .A(n491), .B(n492), .ZN(n715) );
  INV_X1 U617 ( .A(n550), .ZN(n552) );
  AND2_X1 U618 ( .A1(n551), .A2(n552), .ZN(n573) );
  NAND2_X1 U619 ( .A1(G234), .A2(n493), .ZN(n494) );
  XNOR2_X1 U620 ( .A(KEYINPUT20), .B(n494), .ZN(n506) );
  AND2_X1 U621 ( .A1(n506), .A2(G221), .ZN(n496) );
  INV_X1 U622 ( .A(KEYINPUT21), .ZN(n495) );
  XNOR2_X1 U623 ( .A(n496), .B(n495), .ZN(n675) );
  NAND2_X1 U624 ( .A1(n573), .A2(n408), .ZN(n497) );
  XNOR2_X1 U625 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U626 ( .A(n503), .B(n502), .ZN(n505) );
  NAND2_X1 U627 ( .A1(G217), .A2(n506), .ZN(n507) );
  XNOR2_X1 U628 ( .A(KEYINPUT95), .B(KEYINPUT79), .ZN(n513) );
  NAND2_X1 U629 ( .A1(G227), .A2(n741), .ZN(n510) );
  XNOR2_X1 U630 ( .A(n514), .B(n525), .ZN(n713) );
  XNOR2_X2 U631 ( .A(n515), .B(G469), .ZN(n580) );
  NAND2_X1 U632 ( .A1(n516), .A2(G210), .ZN(n517) );
  XNOR2_X1 U633 ( .A(n518), .B(n517), .ZN(n520) );
  XNOR2_X1 U634 ( .A(n519), .B(n520), .ZN(n523) );
  NOR2_X1 U635 ( .A1(n535), .A2(n577), .ZN(n528) );
  NAND2_X1 U636 ( .A1(n533), .A2(n528), .ZN(n530) );
  INV_X1 U637 ( .A(KEYINPUT107), .ZN(n529) );
  INV_X1 U638 ( .A(KEYINPUT6), .ZN(n531) );
  XNOR2_X1 U639 ( .A(n681), .B(n531), .ZN(n604) );
  AND2_X1 U640 ( .A1(n535), .A2(n604), .ZN(n532) );
  NAND2_X1 U641 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U642 ( .A(KEYINPUT33), .B(KEYINPUT72), .Z(n537) );
  XOR2_X1 U643 ( .A(KEYINPUT34), .B(KEYINPUT81), .Z(n540) );
  INV_X1 U644 ( .A(n551), .ZN(n553) );
  NAND2_X1 U645 ( .A1(n553), .A2(n550), .ZN(n542) );
  XOR2_X1 U646 ( .A(KEYINPUT108), .B(n542), .Z(n597) );
  INV_X1 U647 ( .A(n548), .ZN(n545) );
  NAND2_X1 U648 ( .A1(n685), .A2(n545), .ZN(n547) );
  XOR2_X1 U649 ( .A(KEYINPUT31), .B(KEYINPUT97), .Z(n546) );
  XNOR2_X1 U650 ( .A(n547), .B(n546), .ZN(n662) );
  OR2_X1 U651 ( .A1(n566), .A2(n577), .ZN(n549) );
  NOR2_X1 U652 ( .A1(n549), .A2(n548), .ZN(n651) );
  NOR2_X1 U653 ( .A1(n662), .A2(n651), .ZN(n555) );
  XNOR2_X1 U654 ( .A(KEYINPUT106), .B(n661), .ZN(n620) );
  XNOR2_X1 U655 ( .A(KEYINPUT86), .B(n694), .ZN(n554) );
  NOR2_X1 U656 ( .A1(n555), .A2(n554), .ZN(n559) );
  INV_X1 U657 ( .A(n676), .ZN(n575) );
  NAND2_X1 U658 ( .A1(n604), .A2(n575), .ZN(n556) );
  NOR2_X1 U659 ( .A1(n535), .A2(n556), .ZN(n558) );
  AND2_X1 U660 ( .A1(n558), .A2(n557), .ZN(n646) );
  NOR2_X1 U661 ( .A1(n559), .A2(n646), .ZN(n560) );
  NAND2_X1 U662 ( .A1(G953), .A2(G900), .ZN(n563) );
  NAND2_X1 U663 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U664 ( .A(KEYINPUT30), .B(KEYINPUT112), .Z(n567) );
  NAND2_X1 U665 ( .A1(n568), .A2(n362), .ZN(n569) );
  XOR2_X1 U666 ( .A(KEYINPUT38), .B(n616), .Z(n690) );
  XOR2_X1 U667 ( .A(KEYINPUT73), .B(KEYINPUT39), .Z(n570) );
  XNOR2_X1 U668 ( .A(KEYINPUT117), .B(KEYINPUT116), .ZN(n572) );
  INV_X1 U669 ( .A(n573), .ZN(n692) );
  NAND2_X1 U670 ( .A1(n690), .A2(n689), .ZN(n693) );
  NOR2_X1 U671 ( .A1(n692), .A2(n693), .ZN(n574) );
  XNOR2_X1 U672 ( .A(KEYINPUT41), .B(n574), .ZN(n704) );
  XOR2_X1 U673 ( .A(KEYINPUT115), .B(KEYINPUT28), .Z(n579) );
  AND2_X1 U674 ( .A1(n577), .A2(n606), .ZN(n578) );
  XNOR2_X1 U675 ( .A(n579), .B(n578), .ZN(n582) );
  XNOR2_X1 U676 ( .A(n580), .B(KEYINPUT114), .ZN(n581) );
  NAND2_X1 U677 ( .A1(n582), .A2(n581), .ZN(n587) );
  XNOR2_X1 U678 ( .A(KEYINPUT118), .B(KEYINPUT42), .ZN(n583) );
  XNOR2_X1 U679 ( .A(n584), .B(n583), .ZN(n751) );
  INV_X1 U680 ( .A(KEYINPUT47), .ZN(n590) );
  NOR2_X1 U681 ( .A1(n657), .A2(KEYINPUT85), .ZN(n588) );
  NOR2_X1 U682 ( .A1(n694), .A2(n588), .ZN(n589) );
  NOR2_X1 U683 ( .A1(n590), .A2(n589), .ZN(n592) );
  INV_X1 U684 ( .A(KEYINPUT85), .ZN(n594) );
  NOR2_X1 U685 ( .A1(KEYINPUT47), .A2(n594), .ZN(n591) );
  NOR2_X1 U686 ( .A1(n592), .A2(n591), .ZN(n600) );
  XOR2_X1 U687 ( .A(KEYINPUT86), .B(n694), .Z(n593) );
  NAND2_X1 U688 ( .A1(n593), .A2(n590), .ZN(n595) );
  AND2_X1 U689 ( .A1(n597), .A2(n596), .ZN(n598) );
  NAND2_X1 U690 ( .A1(n391), .A2(n598), .ZN(n639) );
  NAND2_X1 U691 ( .A1(n607), .A2(n689), .ZN(n614) );
  INV_X1 U692 ( .A(n616), .ZN(n608) );
  XNOR2_X1 U693 ( .A(n748), .B(n609), .ZN(n610) );
  XNOR2_X1 U694 ( .A(n613), .B(n612), .ZN(n622) );
  NOR2_X1 U695 ( .A1(n535), .A2(n614), .ZN(n615) );
  XNOR2_X1 U696 ( .A(n615), .B(KEYINPUT43), .ZN(n617) );
  NOR2_X1 U697 ( .A1(n617), .A2(n391), .ZN(n618) );
  XNOR2_X1 U698 ( .A(n618), .B(KEYINPUT111), .ZN(n752) );
  NAND2_X1 U699 ( .A1(n619), .A2(n620), .ZN(n664) );
  NAND2_X1 U700 ( .A1(n752), .A2(n664), .ZN(n621) );
  INV_X1 U701 ( .A(KEYINPUT2), .ZN(n668) );
  NAND2_X1 U702 ( .A1(n667), .A2(n668), .ZN(n624) );
  NAND2_X1 U703 ( .A1(n624), .A2(n623), .ZN(n625) );
  INV_X1 U704 ( .A(n723), .ZN(n629) );
  NAND2_X1 U705 ( .A1(n739), .A2(KEYINPUT2), .ZN(n628) );
  NAND2_X1 U706 ( .A1(n718), .A2(G472), .ZN(n631) );
  NAND2_X1 U707 ( .A1(n632), .A2(G953), .ZN(n634) );
  INV_X1 U708 ( .A(KEYINPUT92), .ZN(n633) );
  XOR2_X1 U709 ( .A(G119), .B(KEYINPUT127), .Z(n635) );
  XNOR2_X1 U710 ( .A(n636), .B(n635), .ZN(G21) );
  XNOR2_X1 U711 ( .A(G110), .B(KEYINPUT122), .ZN(n637) );
  XNOR2_X1 U712 ( .A(n638), .B(n637), .ZN(G12) );
  XNOR2_X1 U713 ( .A(n639), .B(G143), .ZN(G45) );
  NAND2_X1 U714 ( .A1(n718), .A2(G210), .ZN(n642) );
  XOR2_X1 U715 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n640) );
  XOR2_X1 U716 ( .A(KEYINPUT125), .B(KEYINPUT59), .Z(n643) );
  XOR2_X1 U717 ( .A(G101), .B(n646), .Z(G3) );
  NAND2_X1 U718 ( .A1(n651), .A2(n659), .ZN(n647) );
  XNOR2_X1 U719 ( .A(n647), .B(G104), .ZN(G6) );
  XOR2_X1 U720 ( .A(KEYINPUT27), .B(KEYINPUT121), .Z(n649) );
  XNOR2_X1 U721 ( .A(G107), .B(KEYINPUT26), .ZN(n648) );
  XNOR2_X1 U722 ( .A(n649), .B(n648), .ZN(n650) );
  XOR2_X1 U723 ( .A(KEYINPUT120), .B(n650), .Z(n653) );
  NAND2_X1 U724 ( .A1(n651), .A2(n661), .ZN(n652) );
  XNOR2_X1 U725 ( .A(n653), .B(n652), .ZN(G9) );
  XOR2_X1 U726 ( .A(KEYINPUT123), .B(KEYINPUT29), .Z(n655) );
  NAND2_X1 U727 ( .A1(n657), .A2(n661), .ZN(n654) );
  XNOR2_X1 U728 ( .A(n655), .B(n654), .ZN(n656) );
  XOR2_X1 U729 ( .A(G128), .B(n656), .Z(G30) );
  NAND2_X1 U730 ( .A1(n657), .A2(n659), .ZN(n658) );
  XNOR2_X1 U731 ( .A(n658), .B(G146), .ZN(G48) );
  NAND2_X1 U732 ( .A1(n662), .A2(n659), .ZN(n660) );
  XNOR2_X1 U733 ( .A(n660), .B(G113), .ZN(G15) );
  NAND2_X1 U734 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U735 ( .A(n663), .B(G116), .ZN(G18) );
  XNOR2_X1 U736 ( .A(G134), .B(n664), .ZN(G36) );
  INV_X1 U737 ( .A(KEYINPUT84), .ZN(n665) );
  NOR2_X1 U738 ( .A1(KEYINPUT2), .A2(n665), .ZN(n666) );
  AND2_X1 U739 ( .A1(n667), .A2(n666), .ZN(n670) );
  NOR2_X1 U740 ( .A1(KEYINPUT84), .A2(n668), .ZN(n669) );
  NOR2_X1 U741 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U742 ( .A(n671), .B(KEYINPUT83), .ZN(n673) );
  NOR2_X1 U743 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U744 ( .A(n674), .B(KEYINPUT87), .ZN(n709) );
  NAND2_X1 U745 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U746 ( .A(n677), .B(KEYINPUT49), .ZN(n683) );
  NOR2_X1 U747 ( .A1(n678), .A2(n535), .ZN(n679) );
  XOR2_X1 U748 ( .A(KEYINPUT50), .B(n679), .Z(n680) );
  NAND2_X1 U749 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U750 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U751 ( .A1(n685), .A2(n684), .ZN(n686) );
  XOR2_X1 U752 ( .A(n686), .B(KEYINPUT124), .Z(n687) );
  XNOR2_X1 U753 ( .A(KEYINPUT51), .B(n687), .ZN(n688) );
  NOR2_X1 U754 ( .A1(n704), .A2(n688), .ZN(n699) );
  NOR2_X1 U755 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U756 ( .A1(n692), .A2(n691), .ZN(n696) );
  NOR2_X1 U757 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U758 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U759 ( .A1(n705), .A2(n697), .ZN(n698) );
  NOR2_X1 U760 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U761 ( .A(KEYINPUT52), .B(n700), .ZN(n703) );
  NAND2_X1 U762 ( .A1(n701), .A2(G952), .ZN(n702) );
  NOR2_X1 U763 ( .A1(n703), .A2(n702), .ZN(n707) );
  NOR2_X1 U764 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U765 ( .A(KEYINPUT53), .B(n710), .ZN(G75) );
  NAND2_X1 U766 ( .A1(n718), .A2(G469), .ZN(n712) );
  XOR2_X1 U767 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n711) );
  NOR2_X1 U768 ( .A1(n714), .A2(n722), .ZN(G54) );
  NAND2_X1 U769 ( .A1(n718), .A2(G478), .ZN(n716) );
  XNOR2_X1 U770 ( .A(n715), .B(n716), .ZN(n717) );
  NOR2_X1 U771 ( .A1(n722), .A2(n717), .ZN(G63) );
  NAND2_X1 U772 ( .A1(n718), .A2(G217), .ZN(n720) );
  XNOR2_X1 U773 ( .A(n719), .B(n720), .ZN(n721) );
  NOR2_X1 U774 ( .A1(n722), .A2(n721), .ZN(G66) );
  NAND2_X1 U775 ( .A1(n723), .A2(n741), .ZN(n727) );
  NAND2_X1 U776 ( .A1(G953), .A2(G224), .ZN(n724) );
  XNOR2_X1 U777 ( .A(KEYINPUT61), .B(n724), .ZN(n725) );
  NAND2_X1 U778 ( .A1(n725), .A2(G898), .ZN(n726) );
  NAND2_X1 U779 ( .A1(n727), .A2(n726), .ZN(n734) );
  XNOR2_X1 U780 ( .A(n728), .B(G101), .ZN(n730) );
  XNOR2_X1 U781 ( .A(n729), .B(n730), .ZN(n732) );
  NOR2_X1 U782 ( .A1(G898), .A2(n741), .ZN(n731) );
  NOR2_X1 U783 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U784 ( .A(n734), .B(n733), .ZN(G69) );
  XNOR2_X1 U785 ( .A(n735), .B(KEYINPUT4), .ZN(n737) );
  XOR2_X1 U786 ( .A(n737), .B(n736), .Z(n743) );
  INV_X1 U787 ( .A(n743), .ZN(n738) );
  XOR2_X1 U788 ( .A(n738), .B(KEYINPUT126), .Z(n740) );
  XNOR2_X1 U789 ( .A(n740), .B(n739), .ZN(n742) );
  NAND2_X1 U790 ( .A1(n742), .A2(n741), .ZN(n747) );
  XOR2_X1 U791 ( .A(G227), .B(n743), .Z(n744) );
  NAND2_X1 U792 ( .A1(n744), .A2(G900), .ZN(n745) );
  NAND2_X1 U793 ( .A1(n745), .A2(G953), .ZN(n746) );
  NAND2_X1 U794 ( .A1(n747), .A2(n746), .ZN(G72) );
  XNOR2_X1 U795 ( .A(n748), .B(G125), .ZN(n749) );
  XNOR2_X1 U796 ( .A(n749), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U797 ( .A(n750), .B(G131), .Z(G33) );
  XOR2_X1 U798 ( .A(G137), .B(n751), .Z(G39) );
  XNOR2_X1 U799 ( .A(G140), .B(n752), .ZN(G42) );
  XOR2_X1 U800 ( .A(G122), .B(n753), .Z(G24) );
endmodule

