//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 0 0 1 0 1 0 1 0 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 1 1 0 0 1 0 0 1 0 1 0 0 0 1 1 1 1 0 0 1 1 1 0 0 1 0 0 0 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n839, new_n840, new_n841, new_n842,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n981,
    new_n982, new_n983;
  INV_X1    g000(.A(G227gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G169gat), .ZN(new_n206));
  INV_X1    g005(.A(G176gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n206), .A2(new_n207), .A3(KEYINPUT23), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT23), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n209), .B1(G169gat), .B2(G176gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT65), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  AOI21_X1  g012(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n208), .B(new_n210), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT24), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n216), .A2(G183gat), .A3(G190gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(G183gat), .A2(G190gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT24), .ZN(new_n219));
  NOR2_X1   g018(.A1(G183gat), .A2(G190gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n217), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT25), .B1(new_n215), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT64), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n223), .A2(G176gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n207), .A2(KEYINPUT64), .ZN(new_n225));
  OAI211_X1 g024(.A(KEYINPUT23), .B(new_n206), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n211), .B(new_n212), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT25), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n226), .A2(new_n227), .A3(new_n228), .A4(new_n210), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n222), .B1(new_n229), .B2(new_n221), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT26), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n232), .A2(new_n206), .A3(new_n207), .ZN(new_n233));
  OAI21_X1  g032(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n233), .B(new_n234), .C1(new_n213), .C2(new_n214), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(new_n218), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT66), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT27), .B(G183gat), .ZN(new_n238));
  INV_X1    g037(.A(G190gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  OR2_X1    g039(.A1(new_n240), .A2(KEYINPUT28), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n235), .A2(new_n242), .A3(new_n218), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n240), .A2(KEYINPUT28), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n237), .A2(new_n241), .A3(new_n243), .A4(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n231), .A2(new_n245), .ZN(new_n246));
  XOR2_X1   g045(.A(G127gat), .B(G134gat), .Z(new_n247));
  NOR2_X1   g046(.A1(new_n247), .A2(KEYINPUT1), .ZN(new_n248));
  INV_X1    g047(.A(G113gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(G120gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(KEYINPUT67), .B(G120gat), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n250), .B1(new_n251), .B2(new_n249), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n248), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G113gat), .B(G120gat), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n247), .B1(KEYINPUT1), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n246), .A2(new_n256), .ZN(new_n257));
  AND2_X1   g056(.A1(new_n253), .A2(new_n255), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n231), .A2(new_n245), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n205), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(KEYINPUT68), .B1(new_n260), .B2(KEYINPUT33), .ZN(new_n261));
  INV_X1    g060(.A(new_n259), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n258), .B1(new_n231), .B2(new_n245), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n204), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT68), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT33), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  XOR2_X1   g066(.A(G15gat), .B(G43gat), .Z(new_n268));
  XNOR2_X1  g067(.A(G71gat), .B(G99gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n264), .A2(KEYINPUT32), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n261), .A2(new_n267), .A3(new_n270), .A4(new_n271), .ZN(new_n272));
  NOR3_X1   g071(.A1(new_n262), .A2(new_n204), .A3(new_n263), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n273), .B(KEYINPUT34), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n270), .A2(KEYINPUT33), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n264), .A2(KEYINPUT32), .A3(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n272), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n278));
  OR2_X1    g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n272), .A2(new_n276), .ZN(new_n280));
  INV_X1    g079(.A(new_n274), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(new_n277), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n279), .B1(new_n283), .B2(KEYINPUT69), .ZN(new_n284));
  XNOR2_X1  g083(.A(G1gat), .B(G29gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n285), .B(G85gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT0), .B(G57gat), .ZN(new_n287));
  XOR2_X1   g086(.A(new_n286), .B(new_n287), .Z(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  XOR2_X1   g088(.A(G141gat), .B(G148gat), .Z(new_n290));
  INV_X1    g089(.A(G155gat), .ZN(new_n291));
  INV_X1    g090(.A(G162gat), .ZN(new_n292));
  OAI21_X1  g091(.A(KEYINPUT2), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G155gat), .B(G162gat), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n290), .A2(new_n293), .A3(new_n295), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n299), .A2(KEYINPUT3), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(KEYINPUT3), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n300), .B1(KEYINPUT72), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT72), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n299), .A2(new_n303), .A3(KEYINPUT3), .ZN(new_n304));
  AND2_X1   g103(.A1(new_n304), .A2(new_n256), .ZN(new_n305));
  AND2_X1   g104(.A1(new_n297), .A2(new_n298), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n258), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT4), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n256), .A2(new_n299), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT4), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI22_X1  g110(.A1(new_n302), .A2(new_n305), .B1(new_n308), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(G225gat), .A2(G233gat), .ZN(new_n313));
  XOR2_X1   g112(.A(KEYINPUT74), .B(KEYINPUT5), .Z(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n312), .A2(new_n313), .A3(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n256), .A2(new_n299), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n307), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n313), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(new_n314), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT73), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n311), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n309), .A2(KEYINPUT73), .A3(new_n310), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n324), .A2(new_n308), .A3(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n320), .B1(new_n302), .B2(new_n305), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n322), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n289), .B1(new_n317), .B2(new_n328), .ZN(new_n329));
  AND2_X1   g128(.A1(new_n326), .A2(new_n327), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n288), .B(new_n316), .C1(new_n330), .C2(new_n322), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT6), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n329), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  OAI211_X1 g132(.A(KEYINPUT6), .B(new_n289), .C1(new_n317), .C2(new_n328), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT71), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT70), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n246), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n231), .A2(new_n245), .A3(KEYINPUT70), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT29), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(G226gat), .A2(G233gat), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n336), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n246), .A2(new_n342), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT29), .ZN(new_n345));
  AND3_X1   g144(.A1(new_n231), .A2(new_n245), .A3(KEYINPUT70), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT70), .B1(new_n231), .B2(new_n245), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n348), .A2(KEYINPUT71), .A3(new_n341), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n343), .A2(new_n344), .A3(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(G197gat), .B(G204gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(KEYINPUT22), .ZN(new_n352));
  NAND2_X1  g151(.A1(G211gat), .A2(G218gat), .ZN(new_n353));
  INV_X1    g152(.A(G211gat), .ZN(new_n354));
  INV_X1    g153(.A(G218gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n352), .A2(new_n353), .A3(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT22), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n353), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(new_n351), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n350), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n338), .A2(new_n342), .A3(new_n339), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n246), .A2(new_n345), .A3(new_n341), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n362), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n363), .A2(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(G8gat), .B(G36gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(G64gat), .B(G92gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n369), .B(new_n370), .ZN(new_n371));
  NOR3_X1   g170(.A1(new_n368), .A2(KEYINPUT30), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n366), .B1(new_n350), .B2(new_n362), .ZN(new_n373));
  INV_X1    g172(.A(new_n371), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT30), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  AOI211_X1 g174(.A(new_n366), .B(new_n371), .C1(new_n350), .C2(new_n362), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n284), .B(new_n335), .C1(new_n372), .C2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(G228gat), .A2(G233gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n357), .B(KEYINPUT76), .ZN(new_n380));
  INV_X1    g179(.A(new_n360), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n345), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT3), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n306), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n362), .B1(new_n300), .B2(KEYINPUT29), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n379), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n361), .A2(KEYINPUT77), .A3(new_n345), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(new_n383), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT77), .B1(new_n361), .B2(new_n345), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n299), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(new_n385), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n387), .B1(new_n379), .B2(new_n392), .ZN(new_n393));
  OR2_X1    g192(.A1(new_n393), .A2(G22gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT78), .ZN(new_n395));
  XNOR2_X1  g194(.A(G78gat), .B(G106gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n396), .B(KEYINPUT31), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n397), .B(G50gat), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n393), .A2(G22gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n394), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n395), .A2(new_n394), .A3(new_n400), .A4(new_n398), .ZN(new_n403));
  AND2_X1   g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  OR3_X1    g203(.A1(new_n378), .A2(KEYINPUT35), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n402), .A2(new_n403), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n406), .A2(new_n277), .A3(new_n282), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT75), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n377), .A2(new_n372), .ZN(new_n409));
  INV_X1    g208(.A(new_n335), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n368), .A2(new_n371), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n373), .A2(new_n374), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n412), .A2(KEYINPUT30), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n375), .A2(new_n376), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n416), .A2(KEYINPUT75), .A3(new_n335), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n407), .B1(new_n411), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT35), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n405), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT83), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT37), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n363), .A2(new_n422), .A3(new_n367), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n361), .B1(new_n364), .B2(new_n365), .ZN(new_n424));
  AOI211_X1 g223(.A(new_n422), .B(new_n424), .C1(new_n350), .C2(new_n361), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT82), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n371), .B(new_n423), .C1(new_n425), .C2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT38), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n350), .A2(new_n361), .ZN(new_n429));
  INV_X1    g228(.A(new_n424), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n429), .A2(KEYINPUT37), .A3(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n428), .B1(new_n431), .B2(KEYINPUT82), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n421), .B1(new_n427), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(KEYINPUT38), .B1(new_n425), .B2(new_n426), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n374), .B1(new_n373), .B2(new_n422), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n431), .A2(KEYINPUT82), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n434), .A2(KEYINPUT83), .A3(new_n435), .A4(new_n436), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n335), .A2(new_n376), .ZN(new_n438));
  INV_X1    g237(.A(new_n435), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n373), .A2(new_n422), .ZN(new_n440));
  OAI21_X1  g239(.A(KEYINPUT38), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n433), .A2(new_n437), .A3(new_n438), .A4(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT79), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n443), .B1(new_n312), .B2(new_n313), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NOR3_X1   g244(.A1(new_n312), .A2(new_n443), .A3(new_n313), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT39), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n319), .A2(new_n320), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n448), .B1(new_n449), .B2(KEYINPUT81), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n447), .B(new_n450), .C1(KEYINPUT81), .C2(new_n449), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT80), .ZN(new_n452));
  AND2_X1   g251(.A1(new_n302), .A2(new_n305), .ZN(new_n453));
  AND2_X1   g252(.A1(new_n308), .A2(new_n311), .ZN(new_n454));
  OAI211_X1 g253(.A(KEYINPUT79), .B(new_n320), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT39), .B1(new_n455), .B2(new_n444), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n452), .B1(new_n457), .B2(new_n288), .ZN(new_n458));
  NOR3_X1   g257(.A1(new_n456), .A2(KEYINPUT80), .A3(new_n289), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n451), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT40), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  OAI211_X1 g261(.A(KEYINPUT40), .B(new_n451), .C1(new_n458), .C2(new_n459), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n409), .A2(new_n329), .A3(new_n462), .A4(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n442), .A2(new_n464), .A3(new_n406), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n411), .A2(new_n404), .A3(new_n417), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT36), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n284), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n283), .A2(KEYINPUT36), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n465), .A2(new_n466), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n420), .A2(new_n472), .ZN(new_n473));
  AND2_X1   g272(.A1(G71gat), .A2(G78gat), .ZN(new_n474));
  NOR2_X1   g273(.A1(G71gat), .A2(G78gat), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  XNOR2_X1  g275(.A(G57gat), .B(G64gat), .ZN(new_n477));
  AOI21_X1  g276(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(G64gat), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(G57gat), .ZN(new_n481));
  INV_X1    g280(.A(G57gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(G64gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(G71gat), .B(G78gat), .ZN(new_n485));
  INV_X1    g284(.A(new_n478), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n479), .A2(new_n487), .A3(KEYINPUT89), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT89), .B1(new_n479), .B2(new_n487), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT21), .ZN(new_n491));
  XNOR2_X1  g290(.A(G15gat), .B(G22gat), .ZN(new_n492));
  INV_X1    g291(.A(G1gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT16), .ZN(new_n494));
  AND2_X1   g293(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n492), .A2(G1gat), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n497), .B(G8gat), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT90), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n491), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n499), .B1(new_n491), .B2(new_n498), .ZN(new_n502));
  OAI21_X1  g301(.A(KEYINPUT88), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n491), .A2(new_n498), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT90), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT88), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n505), .A2(new_n506), .A3(new_n500), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT19), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n479), .A2(new_n487), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n511), .A2(KEYINPUT21), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n503), .A2(new_n507), .A3(KEYINPUT19), .ZN(new_n514));
  AND3_X1   g313(.A1(new_n510), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n513), .B1(new_n510), .B2(new_n514), .ZN(new_n516));
  XOR2_X1   g315(.A(G183gat), .B(G211gat), .Z(new_n517));
  NAND2_X1  g316(.A1(G231gat), .A2(G233gat), .ZN(new_n518));
  XOR2_X1   g317(.A(new_n517), .B(new_n518), .Z(new_n519));
  XOR2_X1   g318(.A(G127gat), .B(G155gat), .Z(new_n520));
  XNOR2_X1  g319(.A(new_n520), .B(KEYINPUT20), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n519), .B(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  OR3_X1    g322(.A1(new_n515), .A2(new_n516), .A3(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n523), .B1(new_n515), .B2(new_n516), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(G99gat), .A2(G106gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT8), .ZN(new_n528));
  NAND2_X1  g327(.A1(G85gat), .A2(G92gat), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT7), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(G85gat), .ZN(new_n532));
  INV_X1    g331(.A(G92gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n528), .A2(new_n531), .A3(new_n534), .A4(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(G99gat), .ZN(new_n537));
  INV_X1    g336(.A(G106gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AND2_X1   g338(.A1(new_n539), .A2(new_n527), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n536), .A2(new_n540), .ZN(new_n541));
  AND3_X1   g340(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n542));
  AOI21_X1  g341(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n539), .A2(new_n527), .ZN(new_n545));
  AOI22_X1  g344(.A1(KEYINPUT8), .A2(new_n527), .B1(new_n532), .B2(new_n533), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n541), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT85), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT86), .ZN(new_n550));
  XNOR2_X1  g349(.A(G43gat), .B(G50gat), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n550), .B1(new_n551), .B2(KEYINPUT15), .ZN(new_n552));
  INV_X1    g351(.A(G29gat), .ZN(new_n553));
  INV_X1    g352(.A(G36gat), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n553), .A2(new_n554), .A3(KEYINPUT14), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT14), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n556), .B1(G29gat), .B2(G36gat), .ZN(new_n557));
  OAI211_X1 g356(.A(new_n555), .B(new_n557), .C1(new_n553), .C2(new_n554), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n549), .B1(new_n552), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n551), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT15), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n559), .B(new_n562), .C1(new_n549), .C2(new_n558), .ZN(new_n563));
  OAI221_X1 g362(.A(new_n549), .B1(new_n560), .B2(new_n561), .C1(new_n552), .C2(new_n558), .ZN(new_n564));
  AND3_X1   g363(.A1(new_n563), .A2(KEYINPUT17), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(KEYINPUT17), .B1(new_n563), .B2(new_n564), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n548), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n563), .A2(new_n564), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n567), .B(new_n568), .C1(new_n548), .C2(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(G134gat), .B(G162gat), .Z(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT91), .ZN(new_n572));
  XOR2_X1   g371(.A(new_n570), .B(new_n572), .Z(new_n573));
  XOR2_X1   g372(.A(G190gat), .B(G218gat), .Z(new_n574));
  AOI21_X1  g373(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n573), .B(new_n576), .Z(new_n577));
  NAND2_X1  g376(.A1(new_n526), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G176gat), .B(G204gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(G148gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(KEYINPUT96), .B(G120gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(KEYINPUT97), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT10), .ZN(new_n585));
  NOR4_X1   g384(.A1(new_n488), .A2(new_n489), .A3(new_n548), .A4(new_n585), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n536), .A2(new_n540), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n545), .B1(new_n544), .B2(new_n546), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT92), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n539), .A2(new_n590), .A3(new_n527), .ZN(new_n591));
  AND3_X1   g390(.A1(new_n479), .A2(new_n487), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n479), .A2(new_n487), .A3(new_n591), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n548), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n593), .A2(new_n585), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT93), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT93), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n593), .A2(new_n598), .A3(new_n585), .A4(new_n595), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n586), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G230gat), .A2(G233gat), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n593), .A2(new_n595), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(new_n602), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n584), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT94), .ZN(new_n608));
  NOR3_X1   g407(.A1(new_n600), .A2(new_n608), .A3(new_n602), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n608), .B1(new_n600), .B2(new_n602), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n583), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  XOR2_X1   g411(.A(new_n606), .B(KEYINPUT95), .Z(new_n613));
  AOI21_X1  g412(.A(new_n607), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n498), .B1(new_n565), .B2(new_n566), .ZN(new_n616));
  NAND2_X1  g415(.A1(G229gat), .A2(G233gat), .ZN(new_n617));
  INV_X1    g416(.A(G8gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n497), .B(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n619), .A2(new_n564), .A3(new_n563), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n616), .A2(new_n617), .A3(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT18), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n569), .A2(new_n498), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n624), .A2(new_n620), .A3(KEYINPUT87), .ZN(new_n625));
  OR3_X1    g424(.A1(new_n569), .A2(new_n498), .A3(KEYINPUT87), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n617), .B(KEYINPUT13), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n625), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n616), .A2(KEYINPUT18), .A3(new_n617), .A4(new_n620), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n623), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G169gat), .B(G197gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G113gat), .B(G141gat), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n634), .B(new_n635), .Z(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT12), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n631), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n623), .A2(new_n637), .A3(new_n629), .A4(new_n630), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n615), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n473), .A2(new_n579), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(KEYINPUT98), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n578), .B1(new_n420), .B2(new_n472), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT98), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n646), .A2(new_n647), .A3(new_n643), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(new_n410), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(G1gat), .ZN(G1324gat));
  INV_X1    g450(.A(KEYINPUT99), .ZN(new_n652));
  XNOR2_X1  g451(.A(KEYINPUT16), .B(G8gat), .ZN(new_n653));
  AOI211_X1 g452(.A(new_n416), .B(new_n653), .C1(new_n645), .C2(new_n648), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n652), .B1(new_n654), .B2(KEYINPUT42), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT42), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n649), .A2(new_n409), .ZN(new_n657));
  OAI211_X1 g456(.A(KEYINPUT99), .B(new_n656), .C1(new_n657), .C2(new_n653), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(G8gat), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n654), .A2(KEYINPUT42), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n655), .A2(new_n658), .A3(new_n659), .A4(new_n660), .ZN(G1325gat));
  AOI21_X1  g460(.A(G15gat), .B1(new_n649), .B2(new_n284), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n471), .B1(new_n645), .B2(new_n648), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n662), .B1(G15gat), .B2(new_n663), .ZN(G1326gat));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n404), .ZN(new_n665));
  XNOR2_X1  g464(.A(KEYINPUT43), .B(G22gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(G1327gat));
  XNOR2_X1  g466(.A(new_n573), .B(new_n576), .ZN(new_n668));
  AND3_X1   g467(.A1(new_n465), .A2(new_n466), .A3(new_n471), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n378), .A2(KEYINPUT35), .A3(new_n404), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n404), .A2(new_n283), .ZN(new_n671));
  AOI21_X1  g470(.A(KEYINPUT75), .B1(new_n416), .B2(new_n335), .ZN(new_n672));
  AOI211_X1 g471(.A(new_n408), .B(new_n410), .C1(new_n414), .C2(new_n415), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n671), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n670), .B1(new_n674), .B2(KEYINPUT35), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n668), .B1(new_n669), .B2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n526), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(new_n643), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n679), .A2(new_n553), .A3(new_n410), .ZN(new_n680));
  XOR2_X1   g479(.A(KEYINPUT100), .B(KEYINPUT45), .Z(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n577), .B1(new_n420), .B2(new_n472), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n678), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(G29gat), .B1(new_n687), .B2(new_n335), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n682), .A2(new_n688), .ZN(G1328gat));
  NAND3_X1  g488(.A1(new_n679), .A2(new_n554), .A3(new_n409), .ZN(new_n690));
  XOR2_X1   g489(.A(new_n690), .B(KEYINPUT46), .Z(new_n691));
  OAI21_X1  g490(.A(G36gat), .B1(new_n687), .B2(new_n416), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(G1329gat));
  INV_X1    g492(.A(KEYINPUT102), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n685), .A2(new_n694), .A3(new_n470), .A4(new_n686), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n676), .A2(new_n684), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n473), .A2(KEYINPUT44), .A3(new_n668), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n696), .A2(new_n470), .A3(new_n697), .A4(new_n686), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(KEYINPUT102), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n695), .A2(new_n699), .A3(G43gat), .ZN(new_n700));
  INV_X1    g499(.A(G43gat), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n679), .A2(new_n701), .A3(new_n284), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n702), .A2(KEYINPUT47), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n698), .A2(G43gat), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(new_n702), .ZN(new_n706));
  XOR2_X1   g505(.A(KEYINPUT101), .B(KEYINPUT47), .Z(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n704), .A2(new_n708), .ZN(G1330gat));
  AND2_X1   g508(.A1(new_n404), .A2(G50gat), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n696), .A2(new_n697), .A3(new_n686), .A4(new_n710), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n676), .A2(new_n406), .A3(new_n678), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n711), .B1(G50gat), .B2(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT48), .ZN(G1331gat));
  NAND4_X1  g513(.A1(new_n473), .A2(new_n579), .A3(new_n642), .A4(new_n615), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT103), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n646), .A2(KEYINPUT103), .A3(new_n642), .A4(new_n615), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n719), .A2(new_n335), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(new_n482), .ZN(G1332gat));
  INV_X1    g520(.A(new_n719), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT49), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n409), .B1(new_n723), .B2(new_n480), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT104), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n722), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n723), .A2(new_n480), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(G1333gat));
  NAND3_X1  g527(.A1(new_n717), .A2(new_n284), .A3(new_n718), .ZN(new_n729));
  INV_X1    g528(.A(G71gat), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n717), .A2(G71gat), .A3(new_n470), .A4(new_n718), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(KEYINPUT50), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT50), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n731), .A2(new_n735), .A3(new_n732), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n736), .ZN(G1334gat));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n404), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(G78gat), .ZN(G1335gat));
  INV_X1    g538(.A(KEYINPUT105), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT51), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n677), .A2(new_n642), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n741), .B1(new_n676), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n526), .A2(new_n641), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n683), .A2(KEYINPUT51), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n614), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(G85gat), .B1(new_n746), .B2(new_n410), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n696), .A2(new_n697), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n744), .A2(new_n615), .ZN(new_n749));
  NOR4_X1   g548(.A1(new_n748), .A2(new_n532), .A3(new_n335), .A4(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n740), .B1(new_n747), .B2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(new_n749), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n685), .A2(G85gat), .A3(new_n410), .A4(new_n752), .ZN(new_n753));
  AOI211_X1 g552(.A(new_n335), .B(new_n614), .C1(new_n743), .C2(new_n745), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n753), .B(KEYINPUT105), .C1(new_n754), .C2(G85gat), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n751), .A2(new_n755), .ZN(G1336gat));
  INV_X1    g555(.A(KEYINPUT106), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n696), .A2(new_n409), .A3(new_n697), .A4(new_n752), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(G92gat), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n416), .A2(G92gat), .ZN(new_n760));
  AND4_X1   g559(.A1(KEYINPUT51), .A2(new_n473), .A3(new_n668), .A4(new_n744), .ZN(new_n761));
  AOI21_X1  g560(.A(KEYINPUT51), .B1(new_n683), .B2(new_n744), .ZN(new_n762));
  OAI211_X1 g561(.A(new_n615), .B(new_n760), .C1(new_n761), .C2(new_n762), .ZN(new_n763));
  AOI211_X1 g562(.A(new_n757), .B(KEYINPUT52), .C1(new_n759), .C2(new_n763), .ZN(new_n764));
  OR2_X1    g563(.A1(new_n757), .A2(KEYINPUT52), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n757), .A2(KEYINPUT52), .ZN(new_n766));
  AND4_X1   g565(.A1(new_n765), .A2(new_n759), .A3(new_n766), .A4(new_n763), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n764), .A2(new_n767), .ZN(G1337gat));
  NAND3_X1  g567(.A1(new_n746), .A2(new_n537), .A3(new_n284), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n748), .A2(new_n471), .A3(new_n749), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n769), .B1(new_n537), .B2(new_n770), .ZN(G1338gat));
  NOR2_X1   g570(.A1(new_n761), .A2(new_n762), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n404), .A2(new_n538), .A3(new_n615), .ZN(new_n774));
  XOR2_X1   g573(.A(new_n774), .B(KEYINPUT107), .Z(new_n775));
  NAND4_X1  g574(.A1(new_n696), .A2(new_n404), .A3(new_n697), .A4(new_n752), .ZN(new_n776));
  AOI22_X1  g575(.A1(new_n773), .A2(new_n775), .B1(new_n776), .B2(G106gat), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT53), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n778), .B1(new_n772), .B2(new_n774), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n776), .A2(G106gat), .ZN(new_n780));
  OAI22_X1  g579(.A1(new_n777), .A2(new_n778), .B1(new_n779), .B2(new_n780), .ZN(G1339gat));
  NAND2_X1  g580(.A1(new_n416), .A2(new_n410), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT110), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT54), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n785), .B1(new_n600), .B2(new_n602), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n597), .A2(new_n599), .ZN(new_n787));
  INV_X1    g586(.A(new_n586), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(KEYINPUT94), .B1(new_n789), .B2(new_n601), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n786), .B1(new_n790), .B2(new_n609), .ZN(new_n791));
  INV_X1    g590(.A(new_n583), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n792), .B1(new_n603), .B2(new_n785), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n791), .A2(KEYINPUT55), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(KEYINPUT108), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT108), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n791), .A2(new_n796), .A3(KEYINPUT55), .A4(new_n793), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n612), .A2(new_n613), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n791), .A2(new_n793), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n798), .A2(new_n641), .A3(new_n800), .A4(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT109), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n625), .A2(new_n626), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n805), .B1(new_n806), .B2(new_n627), .ZN(new_n807));
  AOI211_X1 g606(.A(KEYINPUT109), .B(new_n628), .C1(new_n625), .C2(new_n626), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n617), .B1(new_n616), .B2(new_n620), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n807), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(new_n636), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n640), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n812), .A2(new_n614), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n668), .B1(new_n804), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n799), .B1(new_n795), .B2(new_n797), .ZN(new_n816));
  INV_X1    g615(.A(new_n812), .ZN(new_n817));
  AND4_X1   g616(.A1(new_n668), .A2(new_n816), .A3(new_n817), .A4(new_n803), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n677), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  AND4_X1   g618(.A1(new_n526), .A2(new_n577), .A3(new_n642), .A4(new_n614), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n784), .B1(new_n822), .B2(new_n406), .ZN(new_n823));
  AOI211_X1 g622(.A(KEYINPUT110), .B(new_n404), .C1(new_n819), .C2(new_n821), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n284), .B(new_n783), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(G113gat), .B1(new_n825), .B2(new_n642), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n335), .B1(new_n819), .B2(new_n821), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n671), .ZN(new_n828));
  OR2_X1    g627(.A1(new_n828), .A2(KEYINPUT111), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(KEYINPUT111), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n829), .A2(new_n416), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n641), .A2(new_n249), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n826), .B1(new_n831), .B2(new_n832), .ZN(G1340gat));
  OAI21_X1  g632(.A(G120gat), .B1(new_n825), .B2(new_n614), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n614), .A2(new_n251), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n834), .B1(new_n831), .B2(new_n836), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n837), .B(KEYINPUT112), .ZN(G1341gat));
  INV_X1    g637(.A(G127gat), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n825), .A2(new_n839), .A3(new_n677), .ZN(new_n840));
  INV_X1    g639(.A(new_n831), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n526), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n840), .B1(new_n839), .B2(new_n842), .ZN(G1342gat));
  INV_X1    g642(.A(G134gat), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n829), .A2(new_n844), .A3(new_n416), .A4(new_n830), .ZN(new_n845));
  OAI21_X1  g644(.A(KEYINPUT56), .B1(new_n845), .B2(new_n577), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT113), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OR3_X1    g647(.A1(new_n845), .A2(KEYINPUT56), .A3(new_n577), .ZN(new_n849));
  OAI211_X1 g648(.A(KEYINPUT113), .B(KEYINPUT56), .C1(new_n845), .C2(new_n577), .ZN(new_n850));
  OAI21_X1  g649(.A(G134gat), .B1(new_n825), .B2(new_n577), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n848), .A2(new_n849), .A3(new_n850), .A4(new_n851), .ZN(G1343gat));
  INV_X1    g651(.A(KEYINPUT57), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n804), .A2(new_n814), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(new_n577), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n816), .A2(new_n668), .A3(new_n817), .A4(new_n803), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n526), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n853), .B(new_n404), .C1(new_n857), .C2(new_n820), .ZN(new_n858));
  XNOR2_X1  g657(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n859));
  AOI22_X1  g658(.A1(new_n801), .A2(new_n859), .B1(new_n639), .B2(new_n640), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n813), .B1(new_n816), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n856), .B1(new_n861), .B2(new_n668), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n820), .B1(new_n862), .B2(new_n677), .ZN(new_n863));
  OAI21_X1  g662(.A(KEYINPUT57), .B1(new_n863), .B2(new_n406), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n470), .A2(new_n782), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n858), .A2(new_n864), .A3(new_n641), .A4(new_n865), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n866), .A2(G141gat), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n470), .A2(new_n406), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n827), .A2(new_n868), .ZN(new_n869));
  NOR4_X1   g668(.A1(new_n869), .A2(G141gat), .A3(new_n409), .A4(new_n642), .ZN(new_n870));
  OAI21_X1  g669(.A(KEYINPUT58), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(KEYINPUT58), .B1(new_n866), .B2(G141gat), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT116), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT115), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n869), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n642), .A2(G141gat), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n827), .A2(KEYINPUT115), .A3(new_n868), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n875), .A2(new_n416), .A3(new_n876), .A4(new_n877), .ZN(new_n878));
  AND3_X1   g677(.A1(new_n872), .A2(new_n873), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n873), .B1(new_n872), .B2(new_n878), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n871), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT117), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  OAI211_X1 g682(.A(KEYINPUT117), .B(new_n871), .C1(new_n879), .C2(new_n880), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(G1344gat));
  INV_X1    g684(.A(KEYINPUT59), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n822), .A2(KEYINPUT57), .A3(new_n404), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n853), .B1(new_n863), .B2(new_n406), .ZN(new_n889));
  INV_X1    g688(.A(new_n889), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n615), .B(new_n865), .C1(new_n888), .C2(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n886), .B1(new_n891), .B2(G148gat), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n858), .A2(new_n864), .A3(new_n865), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n886), .B1(new_n893), .B2(new_n614), .ZN(new_n894));
  INV_X1    g693(.A(G148gat), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n875), .A2(new_n877), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n416), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n615), .A2(new_n895), .ZN(new_n899));
  OAI22_X1  g698(.A1(new_n892), .A2(new_n896), .B1(new_n898), .B2(new_n899), .ZN(G1345gat));
  NOR3_X1   g699(.A1(new_n893), .A2(new_n291), .A3(new_n677), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n897), .A2(new_n416), .A3(new_n526), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n901), .B1(new_n902), .B2(new_n291), .ZN(G1346gat));
  OAI21_X1  g702(.A(G162gat), .B1(new_n893), .B2(new_n577), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n668), .A2(new_n292), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n904), .B1(new_n898), .B2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT118), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n906), .B(new_n907), .ZN(G1347gat));
  INV_X1    g707(.A(KEYINPUT119), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n909), .B1(new_n822), .B2(new_n335), .ZN(new_n910));
  AOI211_X1 g709(.A(KEYINPUT119), .B(new_n410), .C1(new_n819), .C2(new_n821), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n409), .B(new_n671), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n913), .A2(new_n206), .A3(new_n641), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n409), .A2(new_n335), .A3(new_n284), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(KEYINPUT120), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n916), .B1(new_n823), .B2(new_n824), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT121), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI211_X1 g718(.A(KEYINPUT121), .B(new_n916), .C1(new_n823), .C2(new_n824), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n921), .A2(new_n641), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n914), .B1(new_n922), .B2(new_n206), .ZN(G1348gat));
  AOI21_X1  g722(.A(G176gat), .B1(new_n913), .B2(new_n615), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n614), .A2(new_n224), .A3(new_n225), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n924), .B1(new_n921), .B2(new_n925), .ZN(G1349gat));
  NAND3_X1  g725(.A1(new_n919), .A2(new_n526), .A3(new_n920), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(G183gat), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT122), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n526), .A2(new_n238), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n929), .B1(new_n913), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n928), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(KEYINPUT60), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT60), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n928), .A2(new_n934), .A3(new_n931), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n933), .A2(new_n935), .ZN(G1350gat));
  NAND3_X1  g735(.A1(new_n913), .A2(new_n239), .A3(new_n668), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT123), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n919), .A2(new_n668), .A3(new_n920), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n939), .A2(KEYINPUT61), .A3(G190gat), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(G190gat), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT61), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n938), .A2(new_n940), .A3(new_n943), .ZN(G1351gat));
  NAND2_X1  g743(.A1(new_n409), .A2(new_n335), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n470), .A2(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n947), .B1(new_n887), .B2(new_n889), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  OAI21_X1  g748(.A(G197gat), .B1(new_n949), .B2(new_n642), .ZN(new_n950));
  OAI211_X1 g749(.A(new_n409), .B(new_n868), .C1(new_n910), .C2(new_n911), .ZN(new_n951));
  OR2_X1    g750(.A1(new_n642), .A2(G197gat), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(G1352gat));
  INV_X1    g752(.A(new_n868), .ZN(new_n954));
  INV_X1    g753(.A(new_n910), .ZN(new_n955));
  INV_X1    g754(.A(new_n911), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  XOR2_X1   g756(.A(KEYINPUT124), .B(G204gat), .Z(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  NAND4_X1  g758(.A1(new_n957), .A2(new_n409), .A3(new_n615), .A4(new_n959), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(KEYINPUT62), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n615), .B1(new_n890), .B2(new_n888), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n958), .B1(new_n962), .B2(new_n947), .ZN(new_n963));
  INV_X1    g762(.A(new_n951), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT62), .ZN(new_n965));
  NAND4_X1  g764(.A1(new_n964), .A2(new_n965), .A3(new_n615), .A4(new_n959), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n961), .A2(new_n963), .A3(new_n966), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT125), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND4_X1  g768(.A1(new_n961), .A2(KEYINPUT125), .A3(new_n963), .A4(new_n966), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(G1353gat));
  NAND3_X1  g770(.A1(new_n964), .A2(new_n354), .A3(new_n526), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n948), .A2(new_n526), .ZN(new_n973));
  AND3_X1   g772(.A1(new_n973), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n974));
  AOI21_X1  g773(.A(KEYINPUT63), .B1(new_n973), .B2(G211gat), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n972), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n976), .A2(KEYINPUT126), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT126), .ZN(new_n978));
  OAI211_X1 g777(.A(new_n978), .B(new_n972), .C1(new_n974), .C2(new_n975), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n977), .A2(new_n979), .ZN(G1354gat));
  OAI21_X1  g779(.A(new_n355), .B1(new_n951), .B2(new_n577), .ZN(new_n981));
  XNOR2_X1  g780(.A(new_n981), .B(KEYINPUT127), .ZN(new_n982));
  NOR3_X1   g781(.A1(new_n949), .A2(new_n355), .A3(new_n577), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n982), .A2(new_n983), .ZN(G1355gat));
endmodule


