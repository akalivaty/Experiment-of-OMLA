//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 1 1 0 0 0 0 1 0 1 1 1 1 0 0 0 0 1 1 1 0 1 1 0 0 0 0 0 0 0 0 1 0 0 1 0 0 1 1 0 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:55 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n692, new_n693,
    new_n694, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984;
  INV_X1    g000(.A(KEYINPUT68), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT66), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  AOI22_X1  g003(.A1(new_n188), .A2(KEYINPUT11), .B1(new_n189), .B2(G137), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT11), .ZN(new_n191));
  INV_X1    g005(.A(G137), .ZN(new_n192));
  AND4_X1   g006(.A1(KEYINPUT66), .A2(new_n191), .A3(new_n192), .A4(G134), .ZN(new_n193));
  AOI22_X1  g007(.A1(KEYINPUT66), .A2(new_n191), .B1(new_n192), .B2(G134), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n190), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G131), .ZN(new_n196));
  INV_X1    g010(.A(G131), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n197), .B(new_n190), .C1(new_n193), .C2(new_n194), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  XOR2_X1   g013(.A(KEYINPUT0), .B(G128), .Z(new_n200));
  AND2_X1   g014(.A1(KEYINPUT65), .A2(G146), .ZN(new_n201));
  NOR2_X1   g015(.A1(KEYINPUT65), .A2(G146), .ZN(new_n202));
  NOR3_X1   g016(.A1(new_n201), .A2(new_n202), .A3(G143), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(G146), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n200), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(G143), .B1(new_n201), .B2(new_n202), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(G143), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n207), .A2(KEYINPUT0), .A3(G128), .A4(new_n210), .ZN(new_n211));
  AND2_X1   g025(.A1(new_n206), .A2(new_n211), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n189), .A2(G137), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(KEYINPUT67), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT67), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n215), .B1(new_n192), .B2(G134), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n214), .B(G131), .C1(new_n213), .C2(new_n216), .ZN(new_n217));
  AND2_X1   g031(.A1(new_n198), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT1), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n207), .A2(new_n219), .A3(G128), .A4(new_n210), .ZN(new_n220));
  INV_X1    g034(.A(G128), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n221), .B1(new_n207), .B2(KEYINPUT1), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n201), .A2(new_n202), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n205), .B1(new_n223), .B2(new_n204), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n220), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  AOI22_X1  g039(.A1(new_n199), .A2(new_n212), .B1(new_n218), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n187), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  XOR2_X1   g042(.A(G116), .B(G119), .Z(new_n229));
  XNOR2_X1  g043(.A(KEYINPUT2), .B(G113), .ZN(new_n230));
  XNOR2_X1  g044(.A(new_n229), .B(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n227), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n206), .A2(new_n211), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n233), .B1(new_n196), .B2(new_n198), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n198), .A2(new_n217), .ZN(new_n235));
  OR2_X1    g049(.A1(KEYINPUT65), .A2(G146), .ZN(new_n236));
  NAND2_X1  g050(.A1(KEYINPUT65), .A2(G146), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n204), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(G128), .B1(new_n238), .B2(new_n219), .ZN(new_n239));
  INV_X1    g053(.A(new_n205), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n236), .A2(new_n237), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n240), .B1(new_n241), .B2(G143), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n235), .B1(new_n243), .B2(new_n220), .ZN(new_n244));
  OAI211_X1 g058(.A(KEYINPUT68), .B(new_n232), .C1(new_n234), .C2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n226), .A2(KEYINPUT30), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n228), .A2(new_n231), .A3(new_n245), .A4(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n231), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n226), .A2(new_n248), .ZN(new_n249));
  AND2_X1   g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT31), .ZN(new_n251));
  XOR2_X1   g065(.A(KEYINPUT26), .B(G101), .Z(new_n252));
  NOR2_X1   g066(.A1(G237), .A2(G953), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G210), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n252), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n255), .B(new_n256), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n250), .A2(KEYINPUT70), .A3(new_n251), .A4(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n247), .A2(new_n249), .A3(new_n257), .ZN(new_n259));
  NOR3_X1   g073(.A1(new_n234), .A2(new_n244), .A3(new_n231), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n199), .A2(new_n212), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n218), .A2(new_n225), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n248), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(KEYINPUT28), .B1(new_n260), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT28), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n249), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n257), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n259), .B1(new_n267), .B2(KEYINPUT31), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n269), .B1(new_n259), .B2(KEYINPUT31), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n258), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(G472), .ZN(new_n272));
  INV_X1    g086(.A(G902), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT32), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n271), .A2(KEYINPUT32), .A3(new_n272), .A4(new_n273), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n264), .A2(new_n257), .A3(new_n266), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT29), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n280), .B(KEYINPUT71), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n247), .A2(new_n249), .ZN(new_n282));
  INV_X1    g096(.A(new_n257), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n284), .A2(new_n279), .A3(new_n278), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n273), .ZN(new_n286));
  OAI21_X1  g100(.A(G472), .B1(new_n281), .B2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n276), .A2(new_n277), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G217), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n289), .B1(G234), .B2(new_n273), .ZN(new_n290));
  OAI21_X1  g104(.A(KEYINPUT23), .B1(new_n221), .B2(G119), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n221), .A2(G119), .ZN(new_n292));
  MUX2_X1   g106(.A(KEYINPUT23), .B(new_n291), .S(new_n292), .Z(new_n293));
  XNOR2_X1  g107(.A(G119), .B(G128), .ZN(new_n294));
  XOR2_X1   g108(.A(KEYINPUT24), .B(G110), .Z(new_n295));
  OAI22_X1  g109(.A1(new_n293), .A2(G110), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT16), .ZN(new_n297));
  INV_X1    g111(.A(G140), .ZN(new_n298));
  OAI21_X1  g112(.A(KEYINPUT72), .B1(new_n298), .B2(G125), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(G125), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G125), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n302), .A2(G140), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(KEYINPUT72), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n297), .B1(new_n301), .B2(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n303), .A2(KEYINPUT16), .ZN(new_n306));
  OAI21_X1  g120(.A(G146), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n302), .A2(G140), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n241), .A2(new_n300), .A3(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n296), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n306), .ZN(new_n311));
  AND3_X1   g125(.A1(new_n298), .A2(KEYINPUT72), .A3(G125), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n312), .B1(new_n300), .B2(new_n299), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n208), .B(new_n311), .C1(new_n313), .C2(new_n297), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n307), .A2(new_n314), .ZN(new_n315));
  AOI22_X1  g129(.A1(new_n293), .A2(G110), .B1(new_n294), .B2(new_n295), .ZN(new_n316));
  AND3_X1   g130(.A1(new_n315), .A2(KEYINPUT73), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(KEYINPUT73), .B1(new_n315), .B2(new_n316), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n310), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT74), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OAI211_X1 g135(.A(KEYINPUT74), .B(new_n310), .C1(new_n317), .C2(new_n318), .ZN(new_n322));
  XNOR2_X1  g136(.A(KEYINPUT22), .B(G137), .ZN(new_n323));
  INV_X1    g137(.A(G953), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n324), .A2(G221), .A3(G234), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n323), .B(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n321), .A2(new_n322), .A3(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n319), .A2(new_n320), .A3(new_n326), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AND3_X1   g144(.A1(new_n330), .A2(KEYINPUT25), .A3(new_n273), .ZN(new_n331));
  AOI21_X1  g145(.A(KEYINPUT25), .B1(new_n330), .B2(new_n273), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n290), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n290), .A2(G902), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n330), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  AND2_X1   g151(.A1(new_n288), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT81), .ZN(new_n339));
  XNOR2_X1  g153(.A(KEYINPUT78), .B(KEYINPUT10), .ZN(new_n340));
  OAI21_X1  g154(.A(G128), .B1(new_n205), .B2(new_n219), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n341), .B1(new_n238), .B2(new_n209), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n342), .A2(new_n220), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT77), .ZN(new_n344));
  INV_X1    g158(.A(G104), .ZN(new_n345));
  AOI22_X1  g159(.A1(new_n344), .A2(KEYINPUT3), .B1(new_n345), .B2(G107), .ZN(new_n346));
  OAI22_X1  g160(.A1(new_n344), .A2(KEYINPUT3), .B1(new_n345), .B2(G107), .ZN(new_n347));
  INV_X1    g161(.A(G101), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT3), .ZN(new_n349));
  INV_X1    g163(.A(G107), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n349), .A2(new_n350), .A3(KEYINPUT77), .A4(G104), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n346), .A2(new_n347), .A3(new_n348), .A4(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n350), .A2(G104), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n345), .A2(G107), .ZN(new_n354));
  OAI21_X1  g168(.A(G101), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n340), .B1(new_n343), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(KEYINPUT79), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT79), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n352), .A2(new_n359), .A3(new_n355), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n358), .A2(new_n225), .A3(KEYINPUT10), .A4(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n346), .A2(new_n347), .A3(new_n351), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(G101), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n363), .A2(KEYINPUT4), .A3(new_n352), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT4), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n362), .A2(new_n365), .A3(G101), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n212), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n357), .A2(new_n361), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n199), .ZN(new_n369));
  INV_X1    g183(.A(new_n199), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n357), .A2(new_n361), .A3(new_n367), .A4(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  XNOR2_X1  g186(.A(G110), .B(G140), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n373), .B(KEYINPUT76), .ZN(new_n374));
  AND2_X1   g188(.A1(new_n324), .A2(G227), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n374), .B(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n372), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n356), .B1(new_n220), .B2(new_n342), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n358), .A2(new_n360), .ZN(new_n380));
  INV_X1    g194(.A(new_n225), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n379), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(KEYINPUT12), .B1(new_n382), .B2(new_n370), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT12), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n225), .B1(new_n358), .B2(new_n360), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n384), .B(new_n199), .C1(new_n385), .C2(new_n379), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n383), .A2(new_n371), .A3(new_n386), .A4(new_n376), .ZN(new_n387));
  AOI21_X1  g201(.A(G902), .B1(new_n378), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G469), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n339), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n383), .A2(new_n371), .A3(new_n386), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n377), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n369), .A2(new_n371), .A3(new_n376), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(KEYINPUT80), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT80), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n392), .A2(new_n396), .A3(new_n393), .ZN(new_n397));
  AOI21_X1  g211(.A(G902), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n390), .B1(new_n398), .B2(new_n389), .ZN(new_n399));
  INV_X1    g213(.A(new_n397), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n396), .B1(new_n392), .B2(new_n393), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n273), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n402), .A2(new_n339), .A3(G469), .ZN(new_n403));
  INV_X1    g217(.A(G952), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n404), .A2(G953), .ZN(new_n405));
  INV_X1    g219(.A(G234), .ZN(new_n406));
  INV_X1    g220(.A(G237), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n405), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  OAI211_X1 g223(.A(G902), .B(G953), .C1(new_n406), .C2(new_n407), .ZN(new_n410));
  XOR2_X1   g224(.A(new_n410), .B(KEYINPUT92), .Z(new_n411));
  XNOR2_X1  g225(.A(KEYINPUT21), .B(G898), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n409), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  XOR2_X1   g228(.A(KEYINPUT9), .B(G234), .Z(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(G221), .B1(new_n416), .B2(G902), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n417), .B(KEYINPUT75), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n399), .A2(new_n403), .A3(new_n414), .A4(new_n419), .ZN(new_n420));
  NOR2_X1   g234(.A1(G475), .A2(G902), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n301), .A2(new_n304), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(G146), .ZN(new_n423));
  NAND2_X1  g237(.A1(KEYINPUT18), .A2(G131), .ZN(new_n424));
  AND4_X1   g238(.A1(G143), .A2(new_n407), .A3(new_n324), .A4(G214), .ZN(new_n425));
  AOI21_X1  g239(.A(G143), .B1(new_n253), .B2(G214), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n424), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n407), .A2(new_n324), .A3(G214), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n204), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n253), .A2(G143), .A3(G214), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n429), .A2(KEYINPUT18), .A3(G131), .A4(new_n430), .ZN(new_n431));
  AOI22_X1  g245(.A1(new_n423), .A2(new_n309), .B1(new_n427), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT19), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n434), .B1(new_n301), .B2(new_n304), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n300), .A2(new_n308), .A3(new_n434), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NOR3_X1   g251(.A1(new_n435), .A2(new_n223), .A3(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT86), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n307), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(G131), .B1(new_n425), .B2(new_n426), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n429), .A2(new_n197), .A3(new_n430), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n241), .B(new_n436), .C1(new_n313), .C2(new_n434), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n443), .B1(new_n444), .B2(KEYINPUT86), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n433), .B1(new_n440), .B2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT87), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(G113), .B(G122), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n449), .B(new_n345), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n433), .B(KEYINPUT87), .C1(new_n440), .C2(new_n445), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n448), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT89), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n315), .A2(KEYINPUT88), .ZN(new_n455));
  MUX2_X1   g269(.A(new_n443), .B(new_n441), .S(KEYINPUT17), .Z(new_n456));
  INV_X1    g270(.A(KEYINPUT88), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n307), .A2(new_n314), .A3(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n455), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n459), .A2(new_n450), .A3(new_n433), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n453), .A2(new_n454), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n454), .B1(new_n453), .B2(new_n460), .ZN(new_n462));
  OAI211_X1 g276(.A(KEYINPUT20), .B(new_n421), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n441), .A2(new_n442), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n464), .B1(new_n438), .B2(new_n439), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n311), .B1(new_n313), .B2(new_n297), .ZN(new_n466));
  AOI22_X1  g280(.A1(new_n444), .A2(KEYINPUT86), .B1(new_n466), .B2(G146), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n432), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n451), .B1(new_n468), .B2(KEYINPUT87), .ZN(new_n469));
  INV_X1    g283(.A(new_n452), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n460), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(new_n421), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT20), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(G475), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n459), .A2(new_n433), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(new_n451), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(new_n460), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n475), .B1(new_n478), .B2(new_n273), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n463), .A2(new_n474), .A3(new_n480), .ZN(new_n481));
  XOR2_X1   g295(.A(G116), .B(G122), .Z(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(G107), .ZN(new_n483));
  XNOR2_X1  g297(.A(G116), .B(G122), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n350), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT13), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n487), .A2(new_n204), .A3(G128), .ZN(new_n488));
  XOR2_X1   g302(.A(G128), .B(G143), .Z(new_n489));
  OAI211_X1 g303(.A(G134), .B(new_n488), .C1(new_n489), .C2(new_n487), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT90), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g307(.A(G128), .B(G143), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(KEYINPUT90), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n493), .A2(new_n189), .A3(new_n495), .ZN(new_n496));
  OR2_X1    g310(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(G116), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n498), .A2(KEYINPUT14), .A3(G122), .ZN(new_n499));
  OAI211_X1 g313(.A(G107), .B(new_n499), .C1(new_n482), .C2(KEYINPUT14), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n189), .B1(new_n493), .B2(new_n495), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n485), .B(new_n500), .C1(new_n496), .C2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n415), .A2(G217), .A3(new_n324), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n504), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n497), .A2(new_n502), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(G478), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n509), .A2(KEYINPUT15), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n508), .A2(KEYINPUT91), .A3(new_n273), .A4(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n508), .A2(KEYINPUT91), .A3(new_n273), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n507), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n506), .B1(new_n497), .B2(new_n502), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n273), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT91), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n510), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n512), .B1(new_n514), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n481), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n229), .A2(new_n230), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT5), .ZN(new_n524));
  INV_X1    g338(.A(G119), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n525), .A3(G116), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n526), .B(KEYINPUT82), .ZN(new_n527));
  INV_X1    g341(.A(G113), .ZN(new_n528));
  XNOR2_X1  g342(.A(G116), .B(G119), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n528), .B1(new_n529), .B2(KEYINPUT5), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n523), .B1(new_n527), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n358), .A2(new_n531), .A3(new_n360), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n364), .A2(new_n231), .A3(new_n366), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  XOR2_X1   g348(.A(G110), .B(G122), .Z(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n535), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n532), .A2(new_n533), .A3(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n536), .A2(KEYINPUT6), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n233), .A2(G125), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n302), .B(new_n220), .C1(new_n222), .C2(new_n224), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n324), .A2(G224), .ZN(new_n543));
  XOR2_X1   g357(.A(new_n543), .B(KEYINPUT83), .Z(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n542), .B(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT6), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n534), .A2(new_n547), .A3(new_n535), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n539), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n544), .A2(KEYINPUT7), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n541), .B(KEYINPUT84), .ZN(new_n551));
  INV_X1    g365(.A(new_n540), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  OR2_X1    g367(.A1(new_n542), .A2(new_n550), .ZN(new_n554));
  XOR2_X1   g368(.A(new_n535), .B(KEYINPUT8), .Z(new_n555));
  INV_X1    g369(.A(new_n532), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n531), .B1(new_n352), .B2(new_n355), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n553), .A2(new_n554), .A3(new_n558), .A4(new_n538), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n549), .A2(new_n273), .A3(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(G210), .B1(G237), .B2(G902), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n549), .A2(new_n559), .A3(new_n273), .A4(new_n561), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(G214), .B1(G237), .B2(G902), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT85), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n565), .A2(KEYINPUT85), .A3(new_n566), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NOR3_X1   g385(.A1(new_n420), .A2(new_n522), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n338), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(G101), .ZN(G3));
  NAND2_X1  g388(.A1(new_n271), .A2(new_n273), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(G472), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n576), .A2(new_n274), .A3(new_n333), .A4(new_n335), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n577), .A2(new_n420), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT33), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n508), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n505), .A2(KEYINPUT33), .A3(new_n507), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT94), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n582), .A2(new_n583), .A3(G478), .A4(new_n273), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n517), .A2(new_n509), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n580), .A2(new_n581), .A3(G478), .A4(new_n273), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(KEYINPUT94), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n584), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  AND3_X1   g402(.A1(new_n481), .A2(new_n588), .A3(KEYINPUT95), .ZN(new_n589));
  AOI21_X1  g403(.A(KEYINPUT95), .B1(new_n481), .B2(new_n588), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT93), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n563), .A2(new_n592), .A3(new_n564), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n560), .A2(KEYINPUT93), .A3(new_n562), .ZN(new_n594));
  AND3_X1   g408(.A1(new_n593), .A2(new_n566), .A3(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n578), .A2(new_n591), .A3(new_n595), .ZN(new_n596));
  XOR2_X1   g410(.A(KEYINPUT34), .B(G104), .Z(new_n597));
  XNOR2_X1  g411(.A(new_n596), .B(new_n597), .ZN(G6));
  NAND2_X1  g412(.A1(new_n463), .A2(new_n480), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n471), .A2(KEYINPUT89), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n453), .A2(new_n454), .A3(new_n460), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(KEYINPUT20), .B1(new_n602), .B2(new_n421), .ZN(new_n603));
  INV_X1    g417(.A(new_n520), .ZN(new_n604));
  NOR3_X1   g418(.A1(new_n599), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n578), .A2(new_n595), .A3(new_n605), .ZN(new_n606));
  XOR2_X1   g420(.A(KEYINPUT35), .B(G107), .Z(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(G9));
  NOR2_X1   g422(.A1(new_n327), .A2(KEYINPUT36), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n319), .B(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n334), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n333), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n612), .A2(new_n576), .A3(new_n274), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT96), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n274), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n272), .B1(new_n271), .B2(new_n273), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n618), .A2(KEYINPUT96), .A3(new_n612), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n572), .A2(new_n615), .A3(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(KEYINPUT97), .B(KEYINPUT37), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(G110), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n620), .B(new_n622), .ZN(G12));
  AND3_X1   g437(.A1(new_n399), .A2(new_n403), .A3(new_n419), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n624), .A2(new_n288), .A3(new_n612), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT98), .ZN(new_n626));
  INV_X1    g440(.A(G900), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n409), .B1(new_n411), .B2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n605), .A2(new_n626), .A3(new_n595), .A4(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n421), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n631), .B1(new_n600), .B2(new_n601), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n479), .B1(new_n632), .B2(KEYINPUT20), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n421), .B1(new_n461), .B2(new_n462), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n473), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n633), .A2(new_n520), .A3(new_n635), .A4(new_n629), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n593), .A2(new_n566), .A3(new_n594), .ZN(new_n637));
  OAI21_X1  g451(.A(KEYINPUT98), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n630), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n625), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(G128), .ZN(G30));
  OAI21_X1  g455(.A(new_n283), .B1(new_n260), .B2(new_n263), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n259), .A2(G472), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(G472), .A2(G902), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(KEYINPUT99), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n276), .A2(new_n277), .A3(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n612), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n565), .B(KEYINPUT38), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n566), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n481), .A2(new_n520), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(new_n628), .B(KEYINPUT39), .Z(new_n655));
  NAND2_X1  g469(.A1(new_n624), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n657), .A2(KEYINPUT40), .ZN(new_n658));
  AND3_X1   g472(.A1(new_n624), .A2(KEYINPUT40), .A3(new_n655), .ZN(new_n659));
  OAI211_X1 g473(.A(new_n649), .B(new_n654), .C1(new_n658), .C2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G143), .ZN(G45));
  NAND3_X1  g475(.A1(new_n624), .A2(new_n288), .A3(new_n612), .ZN(new_n662));
  AND3_X1   g476(.A1(new_n481), .A2(new_n588), .A3(new_n629), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n663), .A2(KEYINPUT100), .A3(new_n595), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT100), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n481), .A2(new_n588), .A3(new_n629), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n665), .B1(new_n666), .B2(new_n637), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n662), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(new_n208), .ZN(G48));
  INV_X1    g484(.A(KEYINPUT101), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n671), .B1(new_n388), .B2(new_n389), .ZN(new_n672));
  INV_X1    g486(.A(new_n387), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n376), .B1(new_n369), .B2(new_n371), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n273), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(G469), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n675), .A2(new_n671), .A3(G469), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n418), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  AND3_X1   g493(.A1(new_n679), .A2(new_n595), .A3(new_n414), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n591), .A2(new_n680), .A3(new_n288), .A4(new_n337), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT41), .B(G113), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G15));
  NAND2_X1  g497(.A1(new_n677), .A2(new_n678), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n419), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n637), .ZN(new_n686));
  NOR4_X1   g500(.A1(new_n599), .A2(new_n603), .A3(new_n604), .A4(new_n413), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n686), .A2(new_n288), .A3(new_n337), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G116), .ZN(G18));
  NAND4_X1  g503(.A1(new_n680), .A2(new_n288), .A3(new_n521), .A4(new_n612), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G119), .ZN(G21));
  NOR3_X1   g505(.A1(new_n653), .A2(new_n637), .A3(new_n413), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n692), .A2(new_n618), .A3(new_n337), .A4(new_n679), .ZN(new_n693));
  XOR2_X1   g507(.A(KEYINPUT102), .B(G122), .Z(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G24));
  NOR4_X1   g509(.A1(new_n613), .A2(new_n637), .A3(new_n685), .A4(new_n666), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(new_n302), .ZN(G27));
  NAND2_X1  g511(.A1(new_n388), .A2(new_n389), .ZN(new_n698));
  NAND2_X1  g512(.A1(G469), .A2(G902), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(KEYINPUT103), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT104), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n393), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n369), .A2(KEYINPUT104), .A3(new_n371), .A4(new_n376), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n392), .A2(new_n703), .A3(G469), .A4(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n698), .A2(new_n701), .A3(new_n705), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n418), .A2(new_n652), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n706), .A2(new_n563), .A3(new_n564), .A4(new_n707), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n666), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n288), .A2(new_n337), .A3(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT42), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n288), .A2(new_n709), .A3(KEYINPUT42), .A4(new_n337), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G131), .ZN(G33));
  INV_X1    g529(.A(KEYINPUT105), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n636), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n288), .A2(new_n337), .A3(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n636), .A2(new_n716), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n720), .A2(new_n708), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  XOR2_X1   g536(.A(KEYINPUT106), .B(G134), .Z(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G36));
  INV_X1    g538(.A(KEYINPUT45), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n725), .B1(new_n400), .B2(new_n401), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n392), .A2(new_n703), .A3(KEYINPUT45), .A4(new_n704), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n726), .A2(G469), .A3(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n728), .A2(KEYINPUT46), .A3(new_n701), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT107), .ZN(new_n730));
  OR2_X1    g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT46), .ZN(new_n732));
  INV_X1    g546(.A(new_n728), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n732), .B1(new_n733), .B2(new_n700), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n729), .A2(new_n730), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n731), .A2(new_n698), .A3(new_n734), .A4(new_n735), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n736), .A2(new_n419), .A3(new_n655), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n565), .A2(new_n652), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n633), .A2(new_n588), .A3(new_n474), .ZN(new_n740));
  OR2_X1    g554(.A1(new_n740), .A2(KEYINPUT43), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(KEYINPUT43), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n743), .A2(new_n618), .A3(new_n648), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n739), .B1(new_n744), .B2(KEYINPUT44), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n737), .B(new_n745), .C1(KEYINPUT44), .C2(new_n744), .ZN(new_n746));
  XNOR2_X1  g560(.A(KEYINPUT108), .B(G137), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G39));
  NAND2_X1  g562(.A1(new_n736), .A2(new_n419), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n749), .A2(KEYINPUT47), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n749), .A2(KEYINPUT47), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n750), .A2(new_n751), .A3(new_n666), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n288), .A2(new_n337), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n752), .A2(new_n738), .A3(new_n753), .ZN(new_n754));
  XOR2_X1   g568(.A(KEYINPUT109), .B(G140), .Z(new_n755));
  XNOR2_X1  g569(.A(new_n754), .B(new_n755), .ZN(G42));
  AND3_X1   g570(.A1(new_n741), .A2(new_n409), .A3(new_n742), .ZN(new_n757));
  INV_X1    g571(.A(new_n577), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n650), .A2(new_n566), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n757), .A2(new_n758), .A3(new_n679), .A4(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT117), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n762), .A2(KEYINPUT50), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT50), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n764), .B1(new_n760), .B2(new_n761), .ZN(new_n765));
  OR2_X1    g579(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT118), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n685), .A2(new_n408), .A3(new_n739), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n768), .A2(new_n742), .A3(new_n741), .ZN(new_n769));
  INV_X1    g583(.A(new_n613), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n647), .A2(new_n336), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n481), .A2(new_n588), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(new_n768), .A3(new_n773), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n766), .A2(new_n767), .A3(new_n771), .A4(new_n774), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n771), .B(new_n774), .C1(new_n763), .C2(new_n765), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(KEYINPUT118), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n684), .A2(new_n418), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n778), .B1(new_n750), .B2(new_n751), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n743), .A2(new_n408), .A3(new_n577), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n779), .A2(new_n738), .A3(new_n780), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n775), .A2(new_n777), .A3(KEYINPUT51), .A4(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n776), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n781), .ZN(new_n784));
  XNOR2_X1  g598(.A(KEYINPUT116), .B(KEYINPUT51), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n780), .A2(new_n686), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n772), .A2(new_n591), .A3(new_n768), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n787), .A2(new_n405), .A3(new_n788), .ZN(new_n789));
  XOR2_X1   g603(.A(new_n789), .B(KEYINPUT119), .Z(new_n790));
  AND3_X1   g604(.A1(new_n782), .A2(new_n786), .A3(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT114), .ZN(new_n793));
  NOR4_X1   g607(.A1(new_n653), .A2(new_n637), .A3(new_n418), .A4(new_n628), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n649), .A2(new_n793), .A3(new_n706), .A4(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n794), .A2(new_n648), .A3(new_n647), .A4(new_n706), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(KEYINPUT114), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n696), .ZN(new_n799));
  AOI21_X1  g613(.A(KEYINPUT100), .B1(new_n663), .B2(new_n595), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n666), .A2(new_n665), .A3(new_n637), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n625), .B1(new_n802), .B2(new_n639), .ZN(new_n803));
  AND4_X1   g617(.A1(new_n792), .A2(new_n798), .A3(new_n799), .A4(new_n803), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n630), .A2(new_n638), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n662), .B1(new_n805), .B2(new_n668), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n806), .A2(new_n696), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n792), .B1(new_n807), .B2(new_n798), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n804), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n571), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT110), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n633), .A2(new_n811), .A3(new_n474), .A4(new_n520), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n481), .A2(new_n588), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n463), .A2(new_n474), .A3(new_n480), .A4(new_n520), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(KEYINPUT110), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n812), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n578), .A2(new_n810), .A3(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n620), .A2(new_n573), .A3(new_n817), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n712), .A2(new_n713), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n681), .A2(new_n690), .A3(new_n688), .A4(new_n693), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n770), .A2(new_n709), .ZN(new_n822));
  INV_X1    g636(.A(new_n721), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n822), .B1(new_n823), .B2(new_n718), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n633), .A2(new_n604), .A3(new_n635), .ZN(new_n825));
  OAI21_X1  g639(.A(KEYINPUT111), .B1(new_n825), .B2(new_n628), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n599), .A2(new_n603), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT111), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n827), .A2(new_n828), .A3(new_n604), .A4(new_n629), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n826), .A2(new_n738), .A3(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(KEYINPUT112), .B1(new_n662), .B2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n830), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT112), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n832), .A2(new_n625), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n824), .B1(new_n831), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT113), .B1(new_n821), .B2(new_n835), .ZN(new_n836));
  AND4_X1   g650(.A1(new_n681), .A2(new_n690), .A3(new_n688), .A4(new_n693), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n812), .A2(new_n813), .A3(new_n815), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n838), .A2(new_n420), .A3(new_n577), .ZN(new_n839));
  AOI22_X1  g653(.A1(new_n839), .A2(new_n810), .B1(new_n338), .B2(new_n572), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n837), .A2(new_n840), .A3(new_n620), .A4(new_n714), .ZN(new_n841));
  AOI22_X1  g655(.A1(new_n719), .A2(new_n721), .B1(new_n770), .B2(new_n709), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n833), .B1(new_n832), .B2(new_n625), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n662), .A2(new_n830), .A3(KEYINPUT112), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n842), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT113), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n841), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n809), .B1(new_n836), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT53), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n846), .B1(new_n841), .B2(new_n845), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n818), .A2(new_n820), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n851), .A2(new_n835), .A3(KEYINPUT113), .A4(new_n714), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT53), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n796), .B(new_n793), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n803), .A2(new_n799), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT52), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n807), .A2(new_n792), .A3(new_n798), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n857), .A2(KEYINPUT115), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT115), .B1(new_n857), .B2(new_n858), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n853), .B(new_n854), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n849), .A2(KEYINPUT54), .A3(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n821), .A2(KEYINPUT53), .A3(new_n835), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n864), .B1(new_n859), .B2(new_n860), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT54), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n857), .A2(new_n858), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n867), .B1(new_n850), .B2(new_n852), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n865), .B(new_n866), .C1(KEYINPUT53), .C2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n769), .A2(new_n338), .ZN(new_n870));
  XOR2_X1   g684(.A(new_n870), .B(KEYINPUT48), .Z(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n791), .A2(new_n862), .A3(new_n869), .A4(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT120), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n404), .A2(new_n324), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n862), .A2(new_n869), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n878), .A2(KEYINPUT120), .A3(new_n791), .A4(new_n872), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n875), .A2(new_n876), .A3(new_n879), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n684), .B(KEYINPUT49), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n650), .A2(new_n740), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n772), .A2(new_n707), .A3(new_n881), .A4(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n880), .A2(new_n883), .ZN(G75));
  AOI21_X1  g698(.A(KEYINPUT53), .B1(new_n853), .B2(new_n809), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT115), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n886), .B1(new_n804), .B2(new_n808), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n857), .A2(new_n858), .A3(KEYINPUT115), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n863), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OAI211_X1 g703(.A(G210), .B(G902), .C1(new_n885), .C2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT121), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n891), .A2(KEYINPUT56), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(KEYINPUT55), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT55), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n890), .A2(new_n895), .A3(new_n892), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n539), .A2(new_n548), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(new_n546), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n324), .A2(G952), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n899), .B1(new_n894), .B2(new_n896), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(G51));
  OAI21_X1  g718(.A(KEYINPUT54), .B1(new_n885), .B2(new_n889), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(new_n869), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n701), .A2(KEYINPUT57), .ZN(new_n907));
  OR2_X1    g721(.A1(new_n701), .A2(KEYINPUT57), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n909), .B1(new_n674), .B2(new_n673), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n848), .A2(new_n854), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n273), .B1(new_n911), .B2(new_n865), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n733), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n902), .B1(new_n910), .B2(new_n913), .ZN(G54));
  NAND3_X1  g728(.A1(new_n912), .A2(KEYINPUT58), .A3(G475), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n915), .B(new_n602), .Z(new_n916));
  NOR2_X1   g730(.A1(new_n916), .A2(new_n902), .ZN(G60));
  NAND2_X1  g731(.A1(G478), .A2(G902), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n918), .B(KEYINPUT59), .Z(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n877), .A2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT123), .ZN(new_n922));
  INV_X1    g736(.A(new_n582), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n919), .B1(new_n862), .B2(new_n869), .ZN(new_n925));
  OAI21_X1  g739(.A(KEYINPUT123), .B1(new_n925), .B2(new_n582), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n866), .B1(new_n911), .B2(new_n865), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n885), .A2(new_n889), .A3(KEYINPUT54), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n582), .B(new_n920), .C1(new_n928), .C2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT122), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n906), .A2(KEYINPUT122), .A3(new_n582), .A4(new_n920), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n902), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n927), .A2(new_n934), .A3(new_n935), .ZN(G63));
  NAND2_X1  g750(.A1(new_n911), .A2(new_n865), .ZN(new_n937));
  NAND2_X1  g751(.A1(G217), .A2(G902), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT60), .Z(new_n939));
  NAND3_X1  g753(.A1(new_n937), .A2(new_n610), .A3(new_n939), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n937), .A2(new_n939), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n935), .B(new_n940), .C1(new_n941), .C2(new_n330), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT124), .ZN(new_n943));
  AOI21_X1  g757(.A(KEYINPUT61), .B1(new_n940), .B2(new_n943), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n942), .B(new_n944), .ZN(G66));
  INV_X1    g759(.A(G224), .ZN(new_n946));
  OAI21_X1  g760(.A(G953), .B1(new_n412), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n947), .B1(new_n851), .B2(G953), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n898), .B1(G898), .B2(new_n324), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n948), .B(new_n949), .ZN(G69));
  NAND3_X1  g764(.A1(new_n228), .A2(new_n246), .A3(new_n245), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT125), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n435), .A2(new_n437), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n952), .B(new_n953), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n754), .A2(new_n746), .ZN(new_n955));
  INV_X1    g769(.A(new_n338), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n956), .A2(new_n637), .A3(new_n653), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n856), .B1(new_n737), .B2(new_n957), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n955), .A2(new_n714), .A3(new_n722), .A4(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n954), .B1(new_n959), .B2(G953), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n627), .A2(new_n324), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n660), .A2(new_n807), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT62), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n962), .B(new_n963), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n657), .A2(new_n338), .A3(new_n738), .A4(new_n816), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n964), .A2(new_n746), .A3(new_n754), .A4(new_n965), .ZN(new_n966));
  AND2_X1   g780(.A1(new_n966), .A2(new_n324), .ZN(new_n967));
  OAI22_X1  g781(.A1(new_n960), .A2(new_n961), .B1(new_n967), .B2(new_n954), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n324), .B1(G227), .B2(G900), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n968), .B(new_n969), .ZN(G72));
  XNOR2_X1  g784(.A(new_n644), .B(KEYINPUT63), .ZN(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(new_n851), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n972), .B1(new_n959), .B2(new_n973), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n250), .B(KEYINPUT126), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n974), .A2(new_n283), .A3(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n972), .B1(new_n966), .B2(new_n973), .ZN(new_n977));
  INV_X1    g791(.A(new_n975), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n977), .A2(new_n257), .A3(new_n978), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n979), .A2(KEYINPUT127), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n979), .A2(KEYINPUT127), .ZN(new_n981));
  OAI211_X1 g795(.A(new_n976), .B(new_n935), .C1(new_n980), .C2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n849), .A2(new_n861), .ZN(new_n983));
  AOI211_X1 g797(.A(new_n971), .B(new_n983), .C1(new_n259), .C2(new_n284), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n982), .A2(new_n984), .ZN(G57));
endmodule


