

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U552 ( .A1(G8), .A2(n733), .ZN(n785) );
  INV_X2 U553 ( .A(n728), .ZN(n733) );
  NOR2_X4 U554 ( .A1(n798), .A2(n800), .ZN(n728) );
  XNOR2_X1 U555 ( .A(n540), .B(n539), .ZN(n639) );
  NOR2_X1 U556 ( .A1(G2105), .A2(G2104), .ZN(n540) );
  NAND2_X1 U557 ( .A1(n639), .A2(G137), .ZN(n545) );
  XNOR2_X1 U558 ( .A(n548), .B(n547), .ZN(n549) );
  INV_X2 U559 ( .A(G2105), .ZN(n536) );
  XNOR2_X1 U560 ( .A(n553), .B(KEYINPUT65), .ZN(n697) );
  BUF_X1 U561 ( .A(n697), .Z(G160) );
  OR2_X1 U562 ( .A1(n785), .A2(n784), .ZN(n520) );
  NOR2_X1 U563 ( .A1(n785), .A2(n764), .ZN(n521) );
  AND2_X1 U564 ( .A1(n928), .A2(n836), .ZN(n522) );
  NOR2_X1 U565 ( .A1(n706), .A2(n705), .ZN(n708) );
  INV_X1 U566 ( .A(KEYINPUT29), .ZN(n726) );
  XNOR2_X1 U567 ( .A(n727), .B(n726), .ZN(n732) );
  AND2_X1 U568 ( .A1(n765), .A2(n521), .ZN(n766) );
  XOR2_X1 U569 ( .A(G1981), .B(G305), .Z(n932) );
  OR2_X1 U570 ( .A1(G164), .A2(G1384), .ZN(n798) );
  INV_X1 U571 ( .A(KEYINPUT104), .ZN(n780) );
  XNOR2_X1 U572 ( .A(KEYINPUT66), .B(KEYINPUT23), .ZN(n547) );
  INV_X1 U573 ( .A(KEYINPUT17), .ZN(n539) );
  BUF_X1 U574 ( .A(n639), .Z(n892) );
  AND2_X2 U575 ( .A1(n536), .A2(G2104), .ZN(n893) );
  NOR2_X1 U576 ( .A1(G651), .A2(n657), .ZN(n663) );
  NOR2_X2 U577 ( .A1(n606), .A2(n605), .ZN(n923) );
  NOR2_X1 U578 ( .A1(n543), .A2(n542), .ZN(G164) );
  INV_X1 U579 ( .A(G651), .ZN(n526) );
  NOR2_X1 U580 ( .A1(G543), .A2(n526), .ZN(n523) );
  XOR2_X2 U581 ( .A(KEYINPUT1), .B(n523), .Z(n662) );
  NAND2_X1 U582 ( .A1(G61), .A2(n662), .ZN(n525) );
  NOR2_X2 U583 ( .A1(G651), .A2(G543), .ZN(n669) );
  NAND2_X1 U584 ( .A1(G86), .A2(n669), .ZN(n524) );
  NAND2_X1 U585 ( .A1(n525), .A2(n524), .ZN(n529) );
  XOR2_X1 U586 ( .A(KEYINPUT0), .B(G543), .Z(n657) );
  NOR2_X2 U587 ( .A1(n657), .A2(n526), .ZN(n660) );
  NAND2_X1 U588 ( .A1(n660), .A2(G73), .ZN(n527) );
  XOR2_X1 U589 ( .A(KEYINPUT2), .B(n527), .Z(n528) );
  NOR2_X1 U590 ( .A1(n529), .A2(n528), .ZN(n531) );
  NAND2_X1 U591 ( .A1(n663), .A2(G48), .ZN(n530) );
  NAND2_X1 U592 ( .A1(n531), .A2(n530), .ZN(G305) );
  NOR2_X4 U593 ( .A1(G2104), .A2(n536), .ZN(n896) );
  NAND2_X1 U594 ( .A1(G126), .A2(n896), .ZN(n533) );
  AND2_X2 U595 ( .A1(G2105), .A2(G2104), .ZN(n898) );
  NAND2_X1 U596 ( .A1(G114), .A2(n898), .ZN(n532) );
  NAND2_X1 U597 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U598 ( .A(KEYINPUT88), .B(n534), .ZN(n535) );
  INV_X1 U599 ( .A(n535), .ZN(n538) );
  NAND2_X1 U600 ( .A1(n893), .A2(G102), .ZN(n537) );
  NAND2_X1 U601 ( .A1(n538), .A2(n537), .ZN(n543) );
  NAND2_X1 U602 ( .A1(G138), .A2(n639), .ZN(n541) );
  XNOR2_X1 U603 ( .A(KEYINPUT89), .B(n541), .ZN(n542) );
  NAND2_X1 U604 ( .A1(G113), .A2(n898), .ZN(n544) );
  NAND2_X1 U605 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U606 ( .A(n546), .B(KEYINPUT67), .ZN(n552) );
  AND2_X1 U607 ( .A1(G125), .A2(n896), .ZN(n550) );
  NAND2_X1 U608 ( .A1(G101), .A2(n893), .ZN(n548) );
  NOR2_X1 U609 ( .A1(n550), .A2(n549), .ZN(n551) );
  NAND2_X1 U610 ( .A1(n552), .A2(n551), .ZN(n553) );
  NAND2_X1 U611 ( .A1(G85), .A2(n669), .ZN(n555) );
  NAND2_X1 U612 ( .A1(G72), .A2(n660), .ZN(n554) );
  NAND2_X1 U613 ( .A1(n555), .A2(n554), .ZN(n559) );
  NAND2_X1 U614 ( .A1(G60), .A2(n662), .ZN(n557) );
  NAND2_X1 U615 ( .A1(G47), .A2(n663), .ZN(n556) );
  NAND2_X1 U616 ( .A1(n557), .A2(n556), .ZN(n558) );
  OR2_X1 U617 ( .A1(n559), .A2(n558), .ZN(G290) );
  XNOR2_X1 U618 ( .A(G2451), .B(G2446), .ZN(n569) );
  XOR2_X1 U619 ( .A(G2430), .B(G2443), .Z(n561) );
  XNOR2_X1 U620 ( .A(G2454), .B(G2435), .ZN(n560) );
  XNOR2_X1 U621 ( .A(n561), .B(n560), .ZN(n565) );
  XOR2_X1 U622 ( .A(G2438), .B(KEYINPUT108), .Z(n563) );
  XNOR2_X1 U623 ( .A(G1348), .B(G1341), .ZN(n562) );
  XNOR2_X1 U624 ( .A(n563), .B(n562), .ZN(n564) );
  XOR2_X1 U625 ( .A(n565), .B(n564), .Z(n567) );
  XNOR2_X1 U626 ( .A(KEYINPUT109), .B(G2427), .ZN(n566) );
  XNOR2_X1 U627 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U628 ( .A(n569), .B(n568), .ZN(n570) );
  AND2_X1 U629 ( .A1(n570), .A2(G14), .ZN(G401) );
  AND2_X1 U630 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U631 ( .A(G57), .ZN(G237) );
  NAND2_X1 U632 ( .A1(G64), .A2(n662), .ZN(n572) );
  NAND2_X1 U633 ( .A1(G52), .A2(n663), .ZN(n571) );
  NAND2_X1 U634 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U635 ( .A(KEYINPUT68), .B(n573), .ZN(n579) );
  NAND2_X1 U636 ( .A1(G90), .A2(n669), .ZN(n575) );
  NAND2_X1 U637 ( .A1(G77), .A2(n660), .ZN(n574) );
  NAND2_X1 U638 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U639 ( .A(KEYINPUT69), .B(n576), .ZN(n577) );
  XNOR2_X1 U640 ( .A(KEYINPUT9), .B(n577), .ZN(n578) );
  NOR2_X1 U641 ( .A1(n579), .A2(n578), .ZN(G171) );
  NAND2_X1 U642 ( .A1(n669), .A2(G89), .ZN(n580) );
  XOR2_X1 U643 ( .A(KEYINPUT4), .B(n580), .Z(n583) );
  NAND2_X1 U644 ( .A1(n660), .A2(G76), .ZN(n581) );
  XOR2_X1 U645 ( .A(KEYINPUT78), .B(n581), .Z(n582) );
  NOR2_X1 U646 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U647 ( .A(KEYINPUT79), .B(n584), .ZN(n585) );
  XNOR2_X1 U648 ( .A(n585), .B(KEYINPUT5), .ZN(n590) );
  NAND2_X1 U649 ( .A1(G63), .A2(n662), .ZN(n587) );
  NAND2_X1 U650 ( .A1(G51), .A2(n663), .ZN(n586) );
  NAND2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U652 ( .A(KEYINPUT6), .B(n588), .Z(n589) );
  NAND2_X1 U653 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U654 ( .A(KEYINPUT7), .B(n591), .ZN(G168) );
  XOR2_X1 U655 ( .A(G168), .B(KEYINPUT8), .Z(n592) );
  XNOR2_X1 U656 ( .A(KEYINPUT80), .B(n592), .ZN(G286) );
  NAND2_X1 U657 ( .A1(G7), .A2(G661), .ZN(n593) );
  XNOR2_X1 U658 ( .A(n593), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U659 ( .A(G223), .B(KEYINPUT71), .ZN(n842) );
  NAND2_X1 U660 ( .A1(n842), .A2(G567), .ZN(n594) );
  XOR2_X1 U661 ( .A(KEYINPUT11), .B(n594), .Z(G234) );
  NAND2_X1 U662 ( .A1(n663), .A2(G43), .ZN(n595) );
  XOR2_X1 U663 ( .A(KEYINPUT74), .B(n595), .Z(n606) );
  XOR2_X1 U664 ( .A(KEYINPUT72), .B(KEYINPUT14), .Z(n597) );
  NAND2_X1 U665 ( .A1(G56), .A2(n662), .ZN(n596) );
  XNOR2_X1 U666 ( .A(n597), .B(n596), .ZN(n603) );
  NAND2_X1 U667 ( .A1(n669), .A2(G81), .ZN(n598) );
  XNOR2_X1 U668 ( .A(n598), .B(KEYINPUT12), .ZN(n600) );
  NAND2_X1 U669 ( .A1(G68), .A2(n660), .ZN(n599) );
  NAND2_X1 U670 ( .A1(n600), .A2(n599), .ZN(n601) );
  XOR2_X1 U671 ( .A(KEYINPUT13), .B(n601), .Z(n602) );
  NOR2_X1 U672 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U673 ( .A(n604), .B(KEYINPUT73), .ZN(n605) );
  NAND2_X1 U674 ( .A1(G860), .A2(n923), .ZN(n607) );
  XOR2_X1 U675 ( .A(KEYINPUT75), .B(n607), .Z(G153) );
  NAND2_X1 U676 ( .A1(G868), .A2(G171), .ZN(n617) );
  NAND2_X1 U677 ( .A1(G54), .A2(n663), .ZN(n614) );
  NAND2_X1 U678 ( .A1(G66), .A2(n662), .ZN(n609) );
  NAND2_X1 U679 ( .A1(G92), .A2(n669), .ZN(n608) );
  NAND2_X1 U680 ( .A1(n609), .A2(n608), .ZN(n612) );
  NAND2_X1 U681 ( .A1(n660), .A2(G79), .ZN(n610) );
  XOR2_X1 U682 ( .A(KEYINPUT76), .B(n610), .Z(n611) );
  NOR2_X1 U683 ( .A1(n612), .A2(n611), .ZN(n613) );
  NAND2_X1 U684 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U685 ( .A(n615), .B(KEYINPUT15), .ZN(n937) );
  INV_X1 U686 ( .A(G868), .ZN(n632) );
  NAND2_X1 U687 ( .A1(n937), .A2(n632), .ZN(n616) );
  NAND2_X1 U688 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U689 ( .A(n618), .B(KEYINPUT77), .ZN(G284) );
  NAND2_X1 U690 ( .A1(G91), .A2(n669), .ZN(n620) );
  NAND2_X1 U691 ( .A1(G78), .A2(n660), .ZN(n619) );
  NAND2_X1 U692 ( .A1(n620), .A2(n619), .ZN(n621) );
  XOR2_X1 U693 ( .A(KEYINPUT70), .B(n621), .Z(n625) );
  NAND2_X1 U694 ( .A1(G65), .A2(n662), .ZN(n623) );
  NAND2_X1 U695 ( .A1(G53), .A2(n663), .ZN(n622) );
  AND2_X1 U696 ( .A1(n623), .A2(n622), .ZN(n624) );
  NAND2_X1 U697 ( .A1(n625), .A2(n624), .ZN(G299) );
  NAND2_X1 U698 ( .A1(G868), .A2(G286), .ZN(n627) );
  NAND2_X1 U699 ( .A1(G299), .A2(n632), .ZN(n626) );
  NAND2_X1 U700 ( .A1(n627), .A2(n626), .ZN(G297) );
  INV_X1 U701 ( .A(G860), .ZN(n628) );
  NAND2_X1 U702 ( .A1(n628), .A2(G559), .ZN(n629) );
  NAND2_X1 U703 ( .A1(n629), .A2(n937), .ZN(n630) );
  XNOR2_X1 U704 ( .A(n630), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U705 ( .A1(n937), .A2(G868), .ZN(n631) );
  NOR2_X1 U706 ( .A1(G559), .A2(n631), .ZN(n634) );
  AND2_X1 U707 ( .A1(n632), .A2(n923), .ZN(n633) );
  NOR2_X1 U708 ( .A1(n634), .A2(n633), .ZN(G282) );
  NAND2_X1 U709 ( .A1(G123), .A2(n896), .ZN(n635) );
  XOR2_X1 U710 ( .A(KEYINPUT18), .B(n635), .Z(n636) );
  XNOR2_X1 U711 ( .A(n636), .B(KEYINPUT81), .ZN(n638) );
  NAND2_X1 U712 ( .A1(G111), .A2(n898), .ZN(n637) );
  NAND2_X1 U713 ( .A1(n638), .A2(n637), .ZN(n643) );
  NAND2_X1 U714 ( .A1(G135), .A2(n892), .ZN(n641) );
  NAND2_X1 U715 ( .A1(G99), .A2(n893), .ZN(n640) );
  NAND2_X1 U716 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U717 ( .A1(n643), .A2(n642), .ZN(n1003) );
  XNOR2_X1 U718 ( .A(n1003), .B(G2096), .ZN(n644) );
  INV_X1 U719 ( .A(G2100), .ZN(n853) );
  NAND2_X1 U720 ( .A1(n644), .A2(n853), .ZN(G156) );
  NAND2_X1 U721 ( .A1(G559), .A2(n937), .ZN(n645) );
  XOR2_X1 U722 ( .A(n923), .B(n645), .Z(n679) );
  NOR2_X1 U723 ( .A1(G860), .A2(n679), .ZN(n653) );
  NAND2_X1 U724 ( .A1(G67), .A2(n662), .ZN(n647) );
  NAND2_X1 U725 ( .A1(G55), .A2(n663), .ZN(n646) );
  NAND2_X1 U726 ( .A1(n647), .A2(n646), .ZN(n651) );
  NAND2_X1 U727 ( .A1(G93), .A2(n669), .ZN(n649) );
  NAND2_X1 U728 ( .A1(G80), .A2(n660), .ZN(n648) );
  NAND2_X1 U729 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U730 ( .A1(n651), .A2(n650), .ZN(n675) );
  XNOR2_X1 U731 ( .A(n675), .B(KEYINPUT82), .ZN(n652) );
  XNOR2_X1 U732 ( .A(n653), .B(n652), .ZN(G145) );
  NAND2_X1 U733 ( .A1(G49), .A2(n663), .ZN(n655) );
  NAND2_X1 U734 ( .A1(G74), .A2(G651), .ZN(n654) );
  NAND2_X1 U735 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U736 ( .A1(n662), .A2(n656), .ZN(n659) );
  NAND2_X1 U737 ( .A1(n657), .A2(G87), .ZN(n658) );
  NAND2_X1 U738 ( .A1(n659), .A2(n658), .ZN(G288) );
  NAND2_X1 U739 ( .A1(G75), .A2(n660), .ZN(n661) );
  XOR2_X1 U740 ( .A(KEYINPUT84), .B(n661), .Z(n668) );
  NAND2_X1 U741 ( .A1(G62), .A2(n662), .ZN(n665) );
  NAND2_X1 U742 ( .A1(G50), .A2(n663), .ZN(n664) );
  NAND2_X1 U743 ( .A1(n665), .A2(n664), .ZN(n666) );
  XOR2_X1 U744 ( .A(KEYINPUT83), .B(n666), .Z(n667) );
  NOR2_X1 U745 ( .A1(n668), .A2(n667), .ZN(n671) );
  NAND2_X1 U746 ( .A1(n669), .A2(G88), .ZN(n670) );
  NAND2_X1 U747 ( .A1(n671), .A2(n670), .ZN(G303) );
  NOR2_X1 U748 ( .A1(G868), .A2(n675), .ZN(n672) );
  XNOR2_X1 U749 ( .A(n672), .B(KEYINPUT85), .ZN(n682) );
  XNOR2_X1 U750 ( .A(KEYINPUT19), .B(G305), .ZN(n673) );
  XNOR2_X1 U751 ( .A(n673), .B(G288), .ZN(n674) );
  XNOR2_X1 U752 ( .A(n675), .B(n674), .ZN(n677) );
  XOR2_X1 U753 ( .A(G290), .B(G303), .Z(n676) );
  XNOR2_X1 U754 ( .A(n677), .B(n676), .ZN(n678) );
  XOR2_X1 U755 ( .A(G299), .B(n678), .Z(n848) );
  XNOR2_X1 U756 ( .A(n848), .B(n679), .ZN(n680) );
  NAND2_X1 U757 ( .A1(G868), .A2(n680), .ZN(n681) );
  NAND2_X1 U758 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U759 ( .A(KEYINPUT86), .B(n683), .ZN(G295) );
  NAND2_X1 U760 ( .A1(G2078), .A2(G2084), .ZN(n684) );
  XOR2_X1 U761 ( .A(KEYINPUT20), .B(n684), .Z(n685) );
  NAND2_X1 U762 ( .A1(G2090), .A2(n685), .ZN(n686) );
  XNOR2_X1 U763 ( .A(KEYINPUT21), .B(n686), .ZN(n687) );
  NAND2_X1 U764 ( .A1(n687), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U765 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U766 ( .A(KEYINPUT87), .B(KEYINPUT22), .Z(n689) );
  NAND2_X1 U767 ( .A1(G132), .A2(G82), .ZN(n688) );
  XNOR2_X1 U768 ( .A(n689), .B(n688), .ZN(n690) );
  NOR2_X1 U769 ( .A1(n690), .A2(G218), .ZN(n691) );
  NAND2_X1 U770 ( .A1(G96), .A2(n691), .ZN(n846) );
  NAND2_X1 U771 ( .A1(n846), .A2(G2106), .ZN(n695) );
  NAND2_X1 U772 ( .A1(G108), .A2(G120), .ZN(n692) );
  NOR2_X1 U773 ( .A1(G237), .A2(n692), .ZN(n693) );
  NAND2_X1 U774 ( .A1(G69), .A2(n693), .ZN(n847) );
  NAND2_X1 U775 ( .A1(n847), .A2(G567), .ZN(n694) );
  NAND2_X1 U776 ( .A1(n695), .A2(n694), .ZN(n922) );
  NAND2_X1 U777 ( .A1(G483), .A2(G661), .ZN(n696) );
  NOR2_X1 U778 ( .A1(n922), .A2(n696), .ZN(n845) );
  NAND2_X1 U779 ( .A1(n845), .A2(G36), .ZN(G176) );
  INV_X1 U780 ( .A(G303), .ZN(G166) );
  NAND2_X1 U781 ( .A1(n697), .A2(G40), .ZN(n800) );
  NAND2_X1 U782 ( .A1(G1996), .A2(n728), .ZN(n698) );
  XNOR2_X1 U783 ( .A(n698), .B(KEYINPUT26), .ZN(n699) );
  NAND2_X1 U784 ( .A1(n733), .A2(G1341), .ZN(n702) );
  NAND2_X1 U785 ( .A1(n699), .A2(n702), .ZN(n700) );
  NAND2_X1 U786 ( .A1(n700), .A2(KEYINPUT98), .ZN(n701) );
  NAND2_X1 U787 ( .A1(n701), .A2(n923), .ZN(n706) );
  INV_X1 U788 ( .A(KEYINPUT26), .ZN(n703) );
  NOR2_X1 U789 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U790 ( .A1(KEYINPUT98), .A2(n704), .ZN(n705) );
  NOR2_X1 U791 ( .A1(n708), .A2(n937), .ZN(n707) );
  XNOR2_X1 U792 ( .A(n707), .B(KEYINPUT99), .ZN(n714) );
  NAND2_X1 U793 ( .A1(n708), .A2(n937), .ZN(n712) );
  NOR2_X1 U794 ( .A1(n728), .A2(G1348), .ZN(n710) );
  NOR2_X1 U795 ( .A1(G2067), .A2(n733), .ZN(n709) );
  NOR2_X1 U796 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U797 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U798 ( .A1(n714), .A2(n713), .ZN(n720) );
  INV_X1 U799 ( .A(G299), .ZN(n722) );
  NAND2_X1 U800 ( .A1(n733), .A2(G1956), .ZN(n717) );
  NAND2_X1 U801 ( .A1(n728), .A2(G2072), .ZN(n715) );
  XOR2_X1 U802 ( .A(KEYINPUT27), .B(n715), .Z(n716) );
  NAND2_X1 U803 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U804 ( .A(n718), .B(KEYINPUT97), .ZN(n721) );
  NAND2_X1 U805 ( .A1(n722), .A2(n721), .ZN(n719) );
  NAND2_X1 U806 ( .A1(n720), .A2(n719), .ZN(n725) );
  NOR2_X1 U807 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U808 ( .A(n723), .B(KEYINPUT28), .Z(n724) );
  NAND2_X1 U809 ( .A1(n725), .A2(n724), .ZN(n727) );
  INV_X1 U810 ( .A(G1961), .ZN(n862) );
  NAND2_X1 U811 ( .A1(n733), .A2(n862), .ZN(n730) );
  XNOR2_X1 U812 ( .A(G2078), .B(KEYINPUT25), .ZN(n954) );
  NAND2_X1 U813 ( .A1(n728), .A2(n954), .ZN(n729) );
  NAND2_X1 U814 ( .A1(n730), .A2(n729), .ZN(n737) );
  NAND2_X1 U815 ( .A1(n737), .A2(G171), .ZN(n731) );
  NAND2_X1 U816 ( .A1(n732), .A2(n731), .ZN(n752) );
  NOR2_X1 U817 ( .A1(G1966), .A2(n785), .ZN(n755) );
  NOR2_X1 U818 ( .A1(G2084), .A2(n733), .ZN(n756) );
  NOR2_X1 U819 ( .A1(n755), .A2(n756), .ZN(n734) );
  NAND2_X1 U820 ( .A1(G8), .A2(n734), .ZN(n735) );
  XNOR2_X1 U821 ( .A(KEYINPUT30), .B(n735), .ZN(n736) );
  NOR2_X1 U822 ( .A1(G168), .A2(n736), .ZN(n739) );
  NOR2_X1 U823 ( .A1(G171), .A2(n737), .ZN(n738) );
  NOR2_X1 U824 ( .A1(n739), .A2(n738), .ZN(n740) );
  XOR2_X1 U825 ( .A(KEYINPUT31), .B(n740), .Z(n753) );
  NOR2_X1 U826 ( .A1(G1971), .A2(n785), .ZN(n741) );
  XNOR2_X1 U827 ( .A(n741), .B(KEYINPUT100), .ZN(n743) );
  NOR2_X1 U828 ( .A1(n733), .A2(G2090), .ZN(n742) );
  NOR2_X1 U829 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U830 ( .A1(n744), .A2(G303), .ZN(n746) );
  AND2_X1 U831 ( .A1(n753), .A2(n746), .ZN(n745) );
  NAND2_X1 U832 ( .A1(n752), .A2(n745), .ZN(n750) );
  INV_X1 U833 ( .A(n746), .ZN(n747) );
  OR2_X1 U834 ( .A1(n747), .A2(G286), .ZN(n748) );
  AND2_X1 U835 ( .A1(n748), .A2(G8), .ZN(n749) );
  NAND2_X1 U836 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U837 ( .A(n751), .B(KEYINPUT32), .ZN(n760) );
  AND2_X1 U838 ( .A1(n753), .A2(n752), .ZN(n754) );
  NOR2_X1 U839 ( .A1(n755), .A2(n754), .ZN(n758) );
  NAND2_X1 U840 ( .A1(G8), .A2(n756), .ZN(n757) );
  NAND2_X1 U841 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U842 ( .A1(n760), .A2(n759), .ZN(n775) );
  NOR2_X1 U843 ( .A1(G1976), .A2(G288), .ZN(n768) );
  NOR2_X1 U844 ( .A1(G1971), .A2(G303), .ZN(n761) );
  NOR2_X1 U845 ( .A1(n768), .A2(n761), .ZN(n926) );
  XOR2_X1 U846 ( .A(n926), .B(KEYINPUT101), .Z(n762) );
  NAND2_X1 U847 ( .A1(n775), .A2(n762), .ZN(n763) );
  XNOR2_X1 U848 ( .A(n763), .B(KEYINPUT102), .ZN(n765) );
  NAND2_X1 U849 ( .A1(G1976), .A2(G288), .ZN(n929) );
  INV_X1 U850 ( .A(n929), .ZN(n764) );
  XNOR2_X1 U851 ( .A(n766), .B(KEYINPUT64), .ZN(n767) );
  NOR2_X1 U852 ( .A1(n767), .A2(KEYINPUT33), .ZN(n771) );
  NAND2_X1 U853 ( .A1(n768), .A2(KEYINPUT33), .ZN(n769) );
  NOR2_X1 U854 ( .A1(n769), .A2(n785), .ZN(n770) );
  NOR2_X1 U855 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U856 ( .A1(n772), .A2(n932), .ZN(n779) );
  NAND2_X1 U857 ( .A1(G8), .A2(G166), .ZN(n773) );
  NOR2_X1 U858 ( .A1(G2090), .A2(n773), .ZN(n774) );
  XNOR2_X1 U859 ( .A(n774), .B(KEYINPUT103), .ZN(n776) );
  NAND2_X1 U860 ( .A1(n776), .A2(n775), .ZN(n777) );
  NAND2_X1 U861 ( .A1(n777), .A2(n785), .ZN(n778) );
  NAND2_X1 U862 ( .A1(n779), .A2(n778), .ZN(n781) );
  XNOR2_X1 U863 ( .A(n781), .B(n780), .ZN(n786) );
  NOR2_X1 U864 ( .A1(G1981), .A2(G305), .ZN(n782) );
  XOR2_X1 U865 ( .A(n782), .B(KEYINPUT96), .Z(n783) );
  XNOR2_X1 U866 ( .A(KEYINPUT24), .B(n783), .ZN(n784) );
  NAND2_X1 U867 ( .A1(n786), .A2(n520), .ZN(n823) );
  NAND2_X1 U868 ( .A1(n893), .A2(G104), .ZN(n787) );
  XOR2_X1 U869 ( .A(KEYINPUT91), .B(n787), .Z(n789) );
  NAND2_X1 U870 ( .A1(n892), .A2(G140), .ZN(n788) );
  NAND2_X1 U871 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U872 ( .A(KEYINPUT34), .B(n790), .ZN(n795) );
  NAND2_X1 U873 ( .A1(G128), .A2(n896), .ZN(n792) );
  NAND2_X1 U874 ( .A1(G116), .A2(n898), .ZN(n791) );
  NAND2_X1 U875 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U876 ( .A(n793), .B(KEYINPUT35), .Z(n794) );
  NOR2_X1 U877 ( .A1(n795), .A2(n794), .ZN(n796) );
  XOR2_X1 U878 ( .A(KEYINPUT36), .B(n796), .Z(n797) );
  XOR2_X1 U879 ( .A(KEYINPUT92), .B(n797), .Z(n906) );
  XNOR2_X1 U880 ( .A(G2067), .B(KEYINPUT37), .ZN(n824) );
  NOR2_X1 U881 ( .A1(n906), .A2(n824), .ZN(n1009) );
  INV_X1 U882 ( .A(n798), .ZN(n799) );
  NOR2_X1 U883 ( .A1(n800), .A2(n799), .ZN(n801) );
  XNOR2_X1 U884 ( .A(n801), .B(KEYINPUT90), .ZN(n836) );
  NAND2_X1 U885 ( .A1(n1009), .A2(n836), .ZN(n834) );
  NAND2_X1 U886 ( .A1(G119), .A2(n896), .ZN(n803) );
  NAND2_X1 U887 ( .A1(G107), .A2(n898), .ZN(n802) );
  NAND2_X1 U888 ( .A1(n803), .A2(n802), .ZN(n808) );
  NAND2_X1 U889 ( .A1(G131), .A2(n892), .ZN(n805) );
  NAND2_X1 U890 ( .A1(G95), .A2(n893), .ZN(n804) );
  NAND2_X1 U891 ( .A1(n805), .A2(n804), .ZN(n806) );
  XOR2_X1 U892 ( .A(KEYINPUT93), .B(n806), .Z(n807) );
  NOR2_X1 U893 ( .A1(n808), .A2(n807), .ZN(n909) );
  INV_X1 U894 ( .A(G1991), .ZN(n863) );
  NOR2_X1 U895 ( .A1(n909), .A2(n863), .ZN(n819) );
  NAND2_X1 U896 ( .A1(G105), .A2(n893), .ZN(n809) );
  XOR2_X1 U897 ( .A(KEYINPUT38), .B(n809), .Z(n815) );
  NAND2_X1 U898 ( .A1(n898), .A2(G117), .ZN(n810) );
  XNOR2_X1 U899 ( .A(n810), .B(KEYINPUT94), .ZN(n812) );
  NAND2_X1 U900 ( .A1(G129), .A2(n896), .ZN(n811) );
  NAND2_X1 U901 ( .A1(n812), .A2(n811), .ZN(n813) );
  XOR2_X1 U902 ( .A(KEYINPUT95), .B(n813), .Z(n814) );
  NOR2_X1 U903 ( .A1(n815), .A2(n814), .ZN(n817) );
  NAND2_X1 U904 ( .A1(n892), .A2(G141), .ZN(n816) );
  NAND2_X1 U905 ( .A1(n817), .A2(n816), .ZN(n905) );
  AND2_X1 U906 ( .A1(G1996), .A2(n905), .ZN(n818) );
  NOR2_X1 U907 ( .A1(n819), .A2(n818), .ZN(n1011) );
  INV_X1 U908 ( .A(n1011), .ZN(n820) );
  NAND2_X1 U909 ( .A1(n836), .A2(n820), .ZN(n825) );
  NAND2_X1 U910 ( .A1(n834), .A2(n825), .ZN(n821) );
  XNOR2_X1 U911 ( .A(G1986), .B(G290), .ZN(n928) );
  NOR2_X1 U912 ( .A1(n821), .A2(n522), .ZN(n822) );
  NAND2_X1 U913 ( .A1(n823), .A2(n822), .ZN(n839) );
  NAND2_X1 U914 ( .A1(n906), .A2(n824), .ZN(n1014) );
  XOR2_X1 U915 ( .A(KEYINPUT39), .B(KEYINPUT106), .Z(n832) );
  NOR2_X1 U916 ( .A1(G1996), .A2(n905), .ZN(n999) );
  INV_X1 U917 ( .A(n825), .ZN(n829) );
  NOR2_X1 U918 ( .A1(G1986), .A2(G290), .ZN(n826) );
  AND2_X1 U919 ( .A1(n863), .A2(n909), .ZN(n1004) );
  NOR2_X1 U920 ( .A1(n826), .A2(n1004), .ZN(n827) );
  XOR2_X1 U921 ( .A(KEYINPUT105), .B(n827), .Z(n828) );
  NOR2_X1 U922 ( .A1(n829), .A2(n828), .ZN(n830) );
  NOR2_X1 U923 ( .A1(n999), .A2(n830), .ZN(n831) );
  XOR2_X1 U924 ( .A(n832), .B(n831), .Z(n833) );
  NAND2_X1 U925 ( .A1(n834), .A2(n833), .ZN(n835) );
  NAND2_X1 U926 ( .A1(n1014), .A2(n835), .ZN(n837) );
  NAND2_X1 U927 ( .A1(n837), .A2(n836), .ZN(n838) );
  NAND2_X1 U928 ( .A1(n839), .A2(n838), .ZN(n841) );
  XOR2_X1 U929 ( .A(KEYINPUT40), .B(KEYINPUT107), .Z(n840) );
  XNOR2_X1 U930 ( .A(n841), .B(n840), .ZN(G329) );
  NAND2_X1 U931 ( .A1(G2106), .A2(n842), .ZN(G217) );
  AND2_X1 U932 ( .A1(G15), .A2(G2), .ZN(n843) );
  NAND2_X1 U933 ( .A1(G661), .A2(n843), .ZN(G259) );
  NAND2_X1 U934 ( .A1(G3), .A2(G1), .ZN(n844) );
  NAND2_X1 U935 ( .A1(n845), .A2(n844), .ZN(G188) );
  XOR2_X1 U936 ( .A(G120), .B(KEYINPUT110), .Z(G236) );
  INV_X1 U938 ( .A(G132), .ZN(G219) );
  INV_X1 U939 ( .A(G108), .ZN(G238) );
  INV_X1 U940 ( .A(G96), .ZN(G221) );
  INV_X1 U941 ( .A(G82), .ZN(G220) );
  NOR2_X1 U942 ( .A1(n847), .A2(n846), .ZN(G325) );
  INV_X1 U943 ( .A(G325), .ZN(G261) );
  INV_X1 U944 ( .A(G171), .ZN(G301) );
  XNOR2_X1 U945 ( .A(n923), .B(G286), .ZN(n849) );
  XNOR2_X1 U946 ( .A(n849), .B(n848), .ZN(n851) );
  XOR2_X1 U947 ( .A(n937), .B(G301), .Z(n850) );
  XNOR2_X1 U948 ( .A(n851), .B(n850), .ZN(n852) );
  NOR2_X1 U949 ( .A1(G37), .A2(n852), .ZN(G397) );
  XNOR2_X1 U950 ( .A(n853), .B(G2096), .ZN(n855) );
  XNOR2_X1 U951 ( .A(KEYINPUT42), .B(G2678), .ZN(n854) );
  XNOR2_X1 U952 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U953 ( .A(KEYINPUT43), .B(G2090), .Z(n857) );
  XNOR2_X1 U954 ( .A(G2067), .B(G2072), .ZN(n856) );
  XNOR2_X1 U955 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U956 ( .A(n859), .B(n858), .Z(n861) );
  XNOR2_X1 U957 ( .A(G2078), .B(G2084), .ZN(n860) );
  XNOR2_X1 U958 ( .A(n861), .B(n860), .ZN(G227) );
  XNOR2_X1 U959 ( .A(G1956), .B(n862), .ZN(n865) );
  XOR2_X1 U960 ( .A(n863), .B(G1981), .Z(n864) );
  XNOR2_X1 U961 ( .A(n865), .B(n864), .ZN(n869) );
  XOR2_X1 U962 ( .A(G1976), .B(G1971), .Z(n867) );
  XNOR2_X1 U963 ( .A(G1986), .B(G1966), .ZN(n866) );
  XNOR2_X1 U964 ( .A(n867), .B(n866), .ZN(n868) );
  XOR2_X1 U965 ( .A(n869), .B(n868), .Z(n871) );
  XNOR2_X1 U966 ( .A(G2474), .B(KEYINPUT41), .ZN(n870) );
  XNOR2_X1 U967 ( .A(n871), .B(n870), .ZN(n872) );
  XNOR2_X1 U968 ( .A(KEYINPUT111), .B(n872), .ZN(n873) );
  XOR2_X1 U969 ( .A(n873), .B(G1996), .Z(G229) );
  NAND2_X1 U970 ( .A1(n896), .A2(G124), .ZN(n874) );
  XNOR2_X1 U971 ( .A(n874), .B(KEYINPUT44), .ZN(n876) );
  NAND2_X1 U972 ( .A1(G136), .A2(n892), .ZN(n875) );
  NAND2_X1 U973 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U974 ( .A(KEYINPUT112), .B(n877), .ZN(n881) );
  NAND2_X1 U975 ( .A1(G112), .A2(n898), .ZN(n879) );
  NAND2_X1 U976 ( .A1(G100), .A2(n893), .ZN(n878) );
  NAND2_X1 U977 ( .A1(n879), .A2(n878), .ZN(n880) );
  NOR2_X1 U978 ( .A1(n881), .A2(n880), .ZN(G162) );
  XNOR2_X1 U979 ( .A(G164), .B(G162), .ZN(n891) );
  NAND2_X1 U980 ( .A1(G130), .A2(n896), .ZN(n883) );
  NAND2_X1 U981 ( .A1(G118), .A2(n898), .ZN(n882) );
  NAND2_X1 U982 ( .A1(n883), .A2(n882), .ZN(n889) );
  NAND2_X1 U983 ( .A1(G142), .A2(n892), .ZN(n885) );
  NAND2_X1 U984 ( .A1(G106), .A2(n893), .ZN(n884) );
  NAND2_X1 U985 ( .A1(n885), .A2(n884), .ZN(n886) );
  XNOR2_X1 U986 ( .A(KEYINPUT45), .B(n886), .ZN(n887) );
  XNOR2_X1 U987 ( .A(KEYINPUT113), .B(n887), .ZN(n888) );
  NOR2_X1 U988 ( .A1(n889), .A2(n888), .ZN(n890) );
  XNOR2_X1 U989 ( .A(n891), .B(n890), .ZN(n904) );
  NAND2_X1 U990 ( .A1(G139), .A2(n892), .ZN(n895) );
  NAND2_X1 U991 ( .A1(G103), .A2(n893), .ZN(n894) );
  NAND2_X1 U992 ( .A1(n895), .A2(n894), .ZN(n903) );
  NAND2_X1 U993 ( .A1(n896), .A2(G127), .ZN(n897) );
  XNOR2_X1 U994 ( .A(n897), .B(KEYINPUT114), .ZN(n900) );
  NAND2_X1 U995 ( .A1(G115), .A2(n898), .ZN(n899) );
  NAND2_X1 U996 ( .A1(n900), .A2(n899), .ZN(n901) );
  XOR2_X1 U997 ( .A(KEYINPUT47), .B(n901), .Z(n902) );
  NOR2_X1 U998 ( .A1(n903), .A2(n902), .ZN(n994) );
  XOR2_X1 U999 ( .A(n904), .B(n994), .Z(n908) );
  XOR2_X1 U1000 ( .A(n906), .B(n905), .Z(n907) );
  XNOR2_X1 U1001 ( .A(n908), .B(n907), .ZN(n914) );
  XOR2_X1 U1002 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n911) );
  XNOR2_X1 U1003 ( .A(n909), .B(n1003), .ZN(n910) );
  XNOR2_X1 U1004 ( .A(n911), .B(n910), .ZN(n912) );
  XNOR2_X1 U1005 ( .A(G160), .B(n912), .ZN(n913) );
  XNOR2_X1 U1006 ( .A(n914), .B(n913), .ZN(n915) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n915), .ZN(G395) );
  NOR2_X1 U1008 ( .A1(G401), .A2(n922), .ZN(n919) );
  NOR2_X1 U1009 ( .A1(G227), .A2(G229), .ZN(n916) );
  XNOR2_X1 U1010 ( .A(KEYINPUT49), .B(n916), .ZN(n917) );
  NOR2_X1 U1011 ( .A1(G397), .A2(n917), .ZN(n918) );
  NAND2_X1 U1012 ( .A1(n919), .A2(n918), .ZN(n920) );
  NOR2_X1 U1013 ( .A1(n920), .A2(G395), .ZN(n921) );
  XNOR2_X1 U1014 ( .A(n921), .B(KEYINPUT115), .ZN(G225) );
  XOR2_X1 U1015 ( .A(KEYINPUT116), .B(G225), .Z(G308) );
  INV_X1 U1016 ( .A(n922), .ZN(G319) );
  INV_X1 U1017 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U1018 ( .A(KEYINPUT56), .B(G16), .ZN(n947) );
  XNOR2_X1 U1019 ( .A(G1341), .B(n923), .ZN(n924) );
  XNOR2_X1 U1020 ( .A(n924), .B(KEYINPUT124), .ZN(n945) );
  NAND2_X1 U1021 ( .A1(G1971), .A2(G303), .ZN(n925) );
  NAND2_X1 U1022 ( .A1(n926), .A2(n925), .ZN(n927) );
  NOR2_X1 U1023 ( .A1(n928), .A2(n927), .ZN(n930) );
  NAND2_X1 U1024 ( .A1(n930), .A2(n929), .ZN(n943) );
  XOR2_X1 U1025 ( .A(G1966), .B(G168), .Z(n931) );
  XNOR2_X1 U1026 ( .A(KEYINPUT123), .B(n931), .ZN(n933) );
  NAND2_X1 U1027 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1028 ( .A(n934), .B(KEYINPUT57), .ZN(n941) );
  XOR2_X1 U1029 ( .A(G299), .B(G1956), .Z(n936) );
  XOR2_X1 U1030 ( .A(G301), .B(G1961), .Z(n935) );
  NAND2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n939) );
  XOR2_X1 U1032 ( .A(G1348), .B(n937), .Z(n938) );
  NOR2_X1 U1033 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1034 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1035 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1036 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1037 ( .A1(n947), .A2(n946), .ZN(n1027) );
  XOR2_X1 U1038 ( .A(G2067), .B(G26), .Z(n948) );
  NAND2_X1 U1039 ( .A1(n948), .A2(G28), .ZN(n951) );
  XOR2_X1 U1040 ( .A(KEYINPUT121), .B(G2072), .Z(n949) );
  XNOR2_X1 U1041 ( .A(G33), .B(n949), .ZN(n950) );
  NOR2_X1 U1042 ( .A1(n951), .A2(n950), .ZN(n958) );
  XOR2_X1 U1043 ( .A(G1991), .B(G25), .Z(n953) );
  XOR2_X1 U1044 ( .A(G1996), .B(G32), .Z(n952) );
  NAND2_X1 U1045 ( .A1(n953), .A2(n952), .ZN(n956) );
  XOR2_X1 U1046 ( .A(G27), .B(n954), .Z(n955) );
  NOR2_X1 U1047 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1048 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1049 ( .A(KEYINPUT53), .B(n959), .ZN(n963) );
  XOR2_X1 U1050 ( .A(G34), .B(KEYINPUT122), .Z(n961) );
  XNOR2_X1 U1051 ( .A(G2084), .B(KEYINPUT54), .ZN(n960) );
  XNOR2_X1 U1052 ( .A(n961), .B(n960), .ZN(n962) );
  NAND2_X1 U1053 ( .A1(n963), .A2(n962), .ZN(n965) );
  XNOR2_X1 U1054 ( .A(G35), .B(G2090), .ZN(n964) );
  NOR2_X1 U1055 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1056 ( .A(KEYINPUT55), .B(n966), .ZN(n968) );
  INV_X1 U1057 ( .A(G29), .ZN(n967) );
  NAND2_X1 U1058 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1059 ( .A1(n969), .A2(G11), .ZN(n1025) );
  XOR2_X1 U1060 ( .A(G5), .B(G1961), .Z(n982) );
  XNOR2_X1 U1061 ( .A(G1348), .B(KEYINPUT59), .ZN(n970) );
  XNOR2_X1 U1062 ( .A(n970), .B(G4), .ZN(n974) );
  XNOR2_X1 U1063 ( .A(G1341), .B(G19), .ZN(n972) );
  XNOR2_X1 U1064 ( .A(G1956), .B(G20), .ZN(n971) );
  NOR2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1066 ( .A1(n974), .A2(n973), .ZN(n977) );
  XOR2_X1 U1067 ( .A(KEYINPUT125), .B(G1981), .Z(n975) );
  XNOR2_X1 U1068 ( .A(G6), .B(n975), .ZN(n976) );
  NOR2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1070 ( .A(KEYINPUT60), .B(n978), .Z(n980) );
  XNOR2_X1 U1071 ( .A(G1966), .B(G21), .ZN(n979) );
  NOR2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n990) );
  XNOR2_X1 U1074 ( .A(G1971), .B(G22), .ZN(n984) );
  XNOR2_X1 U1075 ( .A(G23), .B(G1976), .ZN(n983) );
  NOR2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n987) );
  XOR2_X1 U1077 ( .A(G1986), .B(KEYINPUT126), .Z(n985) );
  XNOR2_X1 U1078 ( .A(G24), .B(n985), .ZN(n986) );
  NAND2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1080 ( .A(KEYINPUT58), .B(n988), .ZN(n989) );
  NOR2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n991) );
  XOR2_X1 U1082 ( .A(KEYINPUT61), .B(n991), .Z(n992) );
  NOR2_X1 U1083 ( .A1(G16), .A2(n992), .ZN(n993) );
  XNOR2_X1 U1084 ( .A(KEYINPUT127), .B(n993), .ZN(n1023) );
  XOR2_X1 U1085 ( .A(G2072), .B(n994), .Z(n996) );
  XOR2_X1 U1086 ( .A(G164), .B(G2078), .Z(n995) );
  NOR2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1088 ( .A(KEYINPUT50), .B(n997), .ZN(n1002) );
  XOR2_X1 U1089 ( .A(G2090), .B(G162), .Z(n998) );
  NOR2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1091 ( .A(KEYINPUT51), .B(n1000), .Z(n1001) );
  NAND2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1017) );
  NOR2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1094 ( .A(KEYINPUT117), .B(n1005), .Z(n1007) );
  XNOR2_X1 U1095 ( .A(G160), .B(G2084), .ZN(n1006) );
  NAND2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(KEYINPUT118), .B(n1010), .ZN(n1012) );
  NAND2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1100 ( .A(n1013), .B(KEYINPUT119), .ZN(n1015) );
  NAND2_X1 U1101 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1102 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1103 ( .A(KEYINPUT52), .B(n1018), .Z(n1019) );
  NOR2_X1 U1104 ( .A1(KEYINPUT55), .A2(n1019), .ZN(n1020) );
  XOR2_X1 U1105 ( .A(KEYINPUT120), .B(n1020), .Z(n1021) );
  NAND2_X1 U1106 ( .A1(n1021), .A2(G29), .ZN(n1022) );
  NAND2_X1 U1107 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1108 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1109 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1110 ( .A(KEYINPUT62), .B(n1028), .ZN(G150) );
  INV_X1 U1111 ( .A(G150), .ZN(G311) );
endmodule

