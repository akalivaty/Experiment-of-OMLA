

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586;

  AND2_X1 U324 ( .A1(n567), .A2(n436), .ZN(n437) );
  XNOR2_X1 U325 ( .A(n345), .B(n344), .ZN(n349) );
  XNOR2_X1 U326 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U327 ( .A(n347), .B(n346), .ZN(n348) );
  INV_X1 U328 ( .A(KEYINPUT11), .ZN(n346) );
  AND2_X1 U329 ( .A1(n363), .A2(n362), .ZN(n364) );
  XNOR2_X1 U330 ( .A(n345), .B(n311), .ZN(n314) );
  XNOR2_X1 U331 ( .A(n393), .B(n392), .ZN(n567) );
  XNOR2_X1 U332 ( .A(KEYINPUT119), .B(KEYINPUT54), .ZN(n392) );
  XNOR2_X1 U333 ( .A(n357), .B(n356), .ZN(n551) );
  XNOR2_X1 U334 ( .A(n349), .B(n348), .ZN(n357) );
  NOR2_X1 U335 ( .A1(n578), .A2(n366), .ZN(n367) );
  INV_X1 U336 ( .A(n542), .ZN(n362) );
  XNOR2_X1 U337 ( .A(KEYINPUT72), .B(KEYINPUT31), .ZN(n311) );
  XNOR2_X1 U338 ( .A(KEYINPUT47), .B(KEYINPUT111), .ZN(n369) );
  INV_X1 U339 ( .A(n441), .ZN(n317) );
  XNOR2_X1 U340 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U341 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U342 ( .A(n320), .B(n319), .ZN(n322) );
  XNOR2_X1 U343 ( .A(n374), .B(n373), .ZN(n525) );
  XOR2_X1 U344 ( .A(KEYINPUT36), .B(n561), .Z(n582) );
  XNOR2_X1 U345 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U346 ( .A(n452), .B(n451), .Z(n524) );
  XNOR2_X1 U347 ( .A(G169GAT), .B(KEYINPUT120), .ZN(n454) );
  XNOR2_X1 U348 ( .A(n455), .B(n454), .ZN(G1348GAT) );
  XOR2_X1 U349 ( .A(G197GAT), .B(G113GAT), .Z(n293) );
  XNOR2_X1 U350 ( .A(G50GAT), .B(G36GAT), .ZN(n292) );
  XNOR2_X1 U351 ( .A(n293), .B(n292), .ZN(n297) );
  XOR2_X1 U352 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n295) );
  XNOR2_X1 U353 ( .A(G22GAT), .B(G141GAT), .ZN(n294) );
  XNOR2_X1 U354 ( .A(n295), .B(n294), .ZN(n296) );
  XNOR2_X1 U355 ( .A(n297), .B(n296), .ZN(n308) );
  XOR2_X1 U356 ( .A(G1GAT), .B(KEYINPUT69), .Z(n299) );
  XNOR2_X1 U357 ( .A(G15GAT), .B(KEYINPUT68), .ZN(n298) );
  XNOR2_X1 U358 ( .A(n299), .B(n298), .ZN(n331) );
  XOR2_X1 U359 ( .A(G169GAT), .B(G8GAT), .Z(n378) );
  XOR2_X1 U360 ( .A(n331), .B(n378), .Z(n301) );
  NAND2_X1 U361 ( .A1(G229GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U362 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U363 ( .A(n302), .B(KEYINPUT67), .Z(n306) );
  XOR2_X1 U364 ( .A(G29GAT), .B(G43GAT), .Z(n304) );
  XNOR2_X1 U365 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n303) );
  XNOR2_X1 U366 ( .A(n304), .B(n303), .ZN(n351) );
  XNOR2_X1 U367 ( .A(n351), .B(KEYINPUT70), .ZN(n305) );
  XNOR2_X1 U368 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U369 ( .A(n308), .B(n307), .ZN(n542) );
  XOR2_X1 U370 ( .A(G85GAT), .B(G92GAT), .Z(n310) );
  XNOR2_X1 U371 ( .A(G99GAT), .B(G106GAT), .ZN(n309) );
  XNOR2_X1 U372 ( .A(n310), .B(n309), .ZN(n345) );
  XOR2_X1 U373 ( .A(G148GAT), .B(G78GAT), .Z(n397) );
  XNOR2_X1 U374 ( .A(n397), .B(KEYINPUT32), .ZN(n312) );
  XNOR2_X1 U375 ( .A(n312), .B(KEYINPUT33), .ZN(n313) );
  XOR2_X1 U376 ( .A(n314), .B(n313), .Z(n320) );
  XNOR2_X1 U377 ( .A(G57GAT), .B(KEYINPUT71), .ZN(n315) );
  XNOR2_X1 U378 ( .A(n315), .B(KEYINPUT13), .ZN(n335) );
  XNOR2_X1 U379 ( .A(G176GAT), .B(G204GAT), .ZN(n316) );
  XNOR2_X1 U380 ( .A(n316), .B(G64GAT), .ZN(n388) );
  XNOR2_X1 U381 ( .A(n335), .B(n388), .ZN(n318) );
  XOR2_X1 U382 ( .A(G120GAT), .B(G71GAT), .Z(n441) );
  NAND2_X1 U383 ( .A1(G230GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U384 ( .A(n322), .B(n321), .ZN(n574) );
  INV_X1 U385 ( .A(KEYINPUT45), .ZN(n359) );
  XOR2_X1 U386 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n324) );
  XNOR2_X1 U387 ( .A(G8GAT), .B(KEYINPUT77), .ZN(n323) );
  XNOR2_X1 U388 ( .A(n324), .B(n323), .ZN(n341) );
  XOR2_X1 U389 ( .A(KEYINPUT78), .B(G64GAT), .Z(n326) );
  XNOR2_X1 U390 ( .A(G78GAT), .B(KEYINPUT79), .ZN(n325) );
  XNOR2_X1 U391 ( .A(n326), .B(n325), .ZN(n330) );
  XOR2_X1 U392 ( .A(G211GAT), .B(G71GAT), .Z(n328) );
  XNOR2_X1 U393 ( .A(G127GAT), .B(G183GAT), .ZN(n327) );
  XNOR2_X1 U394 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U395 ( .A(n330), .B(n329), .ZN(n339) );
  XOR2_X1 U396 ( .A(G22GAT), .B(G155GAT), .Z(n400) );
  XOR2_X1 U397 ( .A(n400), .B(n331), .Z(n333) );
  NAND2_X1 U398 ( .A1(G231GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U399 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U400 ( .A(n334), .B(KEYINPUT76), .Z(n337) );
  XNOR2_X1 U401 ( .A(n335), .B(KEYINPUT15), .ZN(n336) );
  XNOR2_X1 U402 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U403 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U404 ( .A(n341), .B(n340), .ZN(n578) );
  INV_X1 U405 ( .A(n578), .ZN(n484) );
  NAND2_X1 U406 ( .A1(G232GAT), .A2(G233GAT), .ZN(n343) );
  INV_X1 U407 ( .A(KEYINPUT74), .ZN(n342) );
  XOR2_X1 U408 ( .A(G50GAT), .B(G162GAT), .Z(n403) );
  XNOR2_X1 U409 ( .A(n403), .B(KEYINPUT73), .ZN(n347) );
  XNOR2_X1 U410 ( .A(G36GAT), .B(G190GAT), .ZN(n350) );
  XNOR2_X1 U411 ( .A(n350), .B(G218GAT), .ZN(n381) );
  XNOR2_X1 U412 ( .A(n351), .B(n381), .ZN(n355) );
  XOR2_X1 U413 ( .A(KEYINPUT10), .B(KEYINPUT65), .Z(n353) );
  XNOR2_X1 U414 ( .A(G134GAT), .B(KEYINPUT9), .ZN(n352) );
  XOR2_X1 U415 ( .A(n353), .B(n352), .Z(n354) );
  XNOR2_X1 U416 ( .A(n551), .B(KEYINPUT75), .ZN(n561) );
  NOR2_X1 U417 ( .A1(n484), .A2(n582), .ZN(n358) );
  XNOR2_X1 U418 ( .A(n359), .B(n358), .ZN(n360) );
  NOR2_X1 U419 ( .A1(n574), .A2(n360), .ZN(n361) );
  XNOR2_X1 U420 ( .A(n361), .B(KEYINPUT112), .ZN(n363) );
  XNOR2_X1 U421 ( .A(KEYINPUT113), .B(n364), .ZN(n372) );
  XNOR2_X1 U422 ( .A(KEYINPUT41), .B(n574), .ZN(n544) );
  NOR2_X1 U423 ( .A1(n362), .A2(n544), .ZN(n365) );
  XNOR2_X1 U424 ( .A(n365), .B(KEYINPUT46), .ZN(n366) );
  XNOR2_X1 U425 ( .A(KEYINPUT110), .B(n367), .ZN(n368) );
  NAND2_X1 U426 ( .A1(n368), .A2(n551), .ZN(n370) );
  NAND2_X1 U427 ( .A1(n372), .A2(n371), .ZN(n374) );
  XNOR2_X1 U428 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n373) );
  XOR2_X1 U429 ( .A(KEYINPUT76), .B(G92GAT), .Z(n380) );
  XOR2_X1 U430 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n376) );
  XNOR2_X1 U431 ( .A(KEYINPUT84), .B(G183GAT), .ZN(n375) );
  XNOR2_X1 U432 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U433 ( .A(KEYINPUT19), .B(n377), .Z(n446) );
  XNOR2_X1 U434 ( .A(n378), .B(n446), .ZN(n379) );
  XNOR2_X1 U435 ( .A(n380), .B(n379), .ZN(n385) );
  XOR2_X1 U436 ( .A(n381), .B(KEYINPUT94), .Z(n383) );
  NAND2_X1 U437 ( .A1(G226GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U438 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U439 ( .A(n385), .B(n384), .Z(n390) );
  XOR2_X1 U440 ( .A(G211GAT), .B(KEYINPUT87), .Z(n387) );
  XNOR2_X1 U441 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n386) );
  XNOR2_X1 U442 ( .A(n387), .B(n386), .ZN(n402) );
  XNOR2_X1 U443 ( .A(n402), .B(n388), .ZN(n389) );
  XOR2_X1 U444 ( .A(n390), .B(n389), .Z(n512) );
  XOR2_X1 U445 ( .A(KEYINPUT118), .B(n512), .Z(n391) );
  NAND2_X1 U446 ( .A1(n525), .A2(n391), .ZN(n393) );
  XOR2_X1 U447 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n395) );
  XNOR2_X1 U448 ( .A(KEYINPUT24), .B(G204GAT), .ZN(n394) );
  XNOR2_X1 U449 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U450 ( .A(n396), .B(G106GAT), .Z(n399) );
  XNOR2_X1 U451 ( .A(n397), .B(G218GAT), .ZN(n398) );
  XNOR2_X1 U452 ( .A(n399), .B(n398), .ZN(n401) );
  XOR2_X1 U453 ( .A(n401), .B(n400), .Z(n405) );
  XNOR2_X1 U454 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U455 ( .A(n405), .B(n404), .ZN(n409) );
  XOR2_X1 U456 ( .A(KEYINPUT86), .B(KEYINPUT90), .Z(n407) );
  NAND2_X1 U457 ( .A1(G228GAT), .A2(G233GAT), .ZN(n406) );
  XNOR2_X1 U458 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U459 ( .A(n409), .B(n408), .Z(n414) );
  XOR2_X1 U460 ( .A(KEYINPUT89), .B(KEYINPUT88), .Z(n411) );
  XNOR2_X1 U461 ( .A(KEYINPUT3), .B(KEYINPUT2), .ZN(n410) );
  XNOR2_X1 U462 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U463 ( .A(G141GAT), .B(n412), .Z(n430) );
  XNOR2_X1 U464 ( .A(n430), .B(KEYINPUT85), .ZN(n413) );
  XNOR2_X1 U465 ( .A(n414), .B(n413), .ZN(n463) );
  XOR2_X1 U466 ( .A(KEYINPUT81), .B(G134GAT), .Z(n416) );
  XNOR2_X1 U467 ( .A(KEYINPUT0), .B(G127GAT), .ZN(n415) );
  XNOR2_X1 U468 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U469 ( .A(G113GAT), .B(n417), .Z(n448) );
  XOR2_X1 U470 ( .A(G57GAT), .B(G148GAT), .Z(n419) );
  XNOR2_X1 U471 ( .A(G1GAT), .B(G155GAT), .ZN(n418) );
  XNOR2_X1 U472 ( .A(n419), .B(n418), .ZN(n423) );
  XOR2_X1 U473 ( .A(G85GAT), .B(G162GAT), .Z(n421) );
  XNOR2_X1 U474 ( .A(G29GAT), .B(G120GAT), .ZN(n420) );
  XNOR2_X1 U475 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U476 ( .A(n423), .B(n422), .ZN(n434) );
  XOR2_X1 U477 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n425) );
  XNOR2_X1 U478 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n424) );
  XNOR2_X1 U479 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U480 ( .A(KEYINPUT5), .B(n426), .Z(n428) );
  NAND2_X1 U481 ( .A1(G225GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U482 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U483 ( .A(n429), .B(KEYINPUT91), .Z(n432) );
  XNOR2_X1 U484 ( .A(n430), .B(KEYINPUT4), .ZN(n431) );
  XNOR2_X1 U485 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U486 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U487 ( .A(n448), .B(n435), .ZN(n539) );
  INV_X1 U488 ( .A(n539), .ZN(n564) );
  NOR2_X1 U489 ( .A1(n463), .A2(n564), .ZN(n436) );
  XNOR2_X1 U490 ( .A(n437), .B(KEYINPUT55), .ZN(n453) );
  XOR2_X1 U491 ( .A(KEYINPUT20), .B(G190GAT), .Z(n439) );
  XNOR2_X1 U492 ( .A(G43GAT), .B(G99GAT), .ZN(n438) );
  XNOR2_X1 U493 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U494 ( .A(n440), .B(G176GAT), .Z(n443) );
  XNOR2_X1 U495 ( .A(G169GAT), .B(n441), .ZN(n442) );
  XNOR2_X1 U496 ( .A(n443), .B(n442), .ZN(n452) );
  XOR2_X1 U497 ( .A(KEYINPUT82), .B(KEYINPUT83), .Z(n445) );
  NAND2_X1 U498 ( .A1(G227GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U499 ( .A(n445), .B(n444), .ZN(n447) );
  XOR2_X1 U500 ( .A(n447), .B(n446), .Z(n450) );
  XNOR2_X1 U501 ( .A(G15GAT), .B(n448), .ZN(n449) );
  XNOR2_X1 U502 ( .A(n450), .B(n449), .ZN(n451) );
  NOR2_X2 U503 ( .A1(n453), .A2(n524), .ZN(n560) );
  NAND2_X1 U504 ( .A1(n542), .A2(n560), .ZN(n455) );
  NOR2_X1 U505 ( .A1(n574), .A2(n362), .ZN(n489) );
  INV_X1 U506 ( .A(n524), .ZN(n459) );
  XNOR2_X1 U507 ( .A(n512), .B(KEYINPUT27), .ZN(n465) );
  NOR2_X1 U508 ( .A1(n465), .A2(n539), .ZN(n457) );
  XOR2_X1 U509 ( .A(n463), .B(KEYINPUT66), .Z(n456) );
  XNOR2_X1 U510 ( .A(KEYINPUT28), .B(n456), .ZN(n520) );
  NAND2_X1 U511 ( .A1(n457), .A2(n520), .ZN(n523) );
  XOR2_X1 U512 ( .A(KEYINPUT95), .B(n523), .Z(n458) );
  NOR2_X1 U513 ( .A1(n459), .A2(n458), .ZN(n469) );
  NOR2_X1 U514 ( .A1(n524), .A2(n512), .ZN(n460) );
  NOR2_X1 U515 ( .A1(n463), .A2(n460), .ZN(n461) );
  XOR2_X1 U516 ( .A(n461), .B(KEYINPUT96), .Z(n462) );
  XNOR2_X1 U517 ( .A(KEYINPUT25), .B(n462), .ZN(n466) );
  NAND2_X1 U518 ( .A1(n463), .A2(n524), .ZN(n464) );
  XNOR2_X1 U519 ( .A(n464), .B(KEYINPUT26), .ZN(n565) );
  NOR2_X1 U520 ( .A1(n565), .A2(n465), .ZN(n538) );
  NOR2_X1 U521 ( .A1(n466), .A2(n538), .ZN(n467) );
  NOR2_X1 U522 ( .A1(n564), .A2(n467), .ZN(n468) );
  NOR2_X1 U523 ( .A1(n469), .A2(n468), .ZN(n483) );
  OR2_X1 U524 ( .A1(n484), .A2(n561), .ZN(n470) );
  XNOR2_X1 U525 ( .A(n470), .B(KEYINPUT80), .ZN(n471) );
  XNOR2_X1 U526 ( .A(n471), .B(KEYINPUT16), .ZN(n472) );
  NOR2_X1 U527 ( .A1(n483), .A2(n472), .ZN(n501) );
  NAND2_X1 U528 ( .A1(n489), .A2(n501), .ZN(n481) );
  NOR2_X1 U529 ( .A1(n539), .A2(n481), .ZN(n473) );
  XOR2_X1 U530 ( .A(KEYINPUT34), .B(n473), .Z(n474) );
  XNOR2_X1 U531 ( .A(G1GAT), .B(n474), .ZN(G1324GAT) );
  NOR2_X1 U532 ( .A1(n512), .A2(n481), .ZN(n476) );
  XNOR2_X1 U533 ( .A(KEYINPUT97), .B(KEYINPUT98), .ZN(n475) );
  XNOR2_X1 U534 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U535 ( .A(G8GAT), .B(n477), .ZN(G1325GAT) );
  NOR2_X1 U536 ( .A1(n524), .A2(n481), .ZN(n479) );
  XNOR2_X1 U537 ( .A(KEYINPUT35), .B(KEYINPUT99), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n479), .B(n478), .ZN(n480) );
  XOR2_X1 U539 ( .A(G15GAT), .B(n480), .Z(G1326GAT) );
  NOR2_X1 U540 ( .A1(n520), .A2(n481), .ZN(n482) );
  XOR2_X1 U541 ( .A(G22GAT), .B(n482), .Z(G1327GAT) );
  NOR2_X1 U542 ( .A1(n483), .A2(n582), .ZN(n485) );
  NAND2_X1 U543 ( .A1(n485), .A2(n484), .ZN(n488) );
  XOR2_X1 U544 ( .A(KEYINPUT102), .B(KEYINPUT37), .Z(n486) );
  XNOR2_X1 U545 ( .A(KEYINPUT101), .B(n486), .ZN(n487) );
  XNOR2_X1 U546 ( .A(n488), .B(n487), .ZN(n509) );
  NAND2_X1 U547 ( .A1(n509), .A2(n489), .ZN(n490) );
  XNOR2_X1 U548 ( .A(n490), .B(KEYINPUT38), .ZN(n499) );
  NOR2_X1 U549 ( .A1(n499), .A2(n539), .ZN(n492) );
  XNOR2_X1 U550 ( .A(KEYINPUT100), .B(KEYINPUT39), .ZN(n491) );
  XNOR2_X1 U551 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U552 ( .A(G29GAT), .B(n493), .ZN(G1328GAT) );
  NOR2_X1 U553 ( .A1(n499), .A2(n512), .ZN(n495) );
  XNOR2_X1 U554 ( .A(G36GAT), .B(KEYINPUT103), .ZN(n494) );
  XNOR2_X1 U555 ( .A(n495), .B(n494), .ZN(G1329GAT) );
  XNOR2_X1 U556 ( .A(KEYINPUT104), .B(KEYINPUT40), .ZN(n497) );
  NOR2_X1 U557 ( .A1(n524), .A2(n499), .ZN(n496) );
  XNOR2_X1 U558 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U559 ( .A(G43GAT), .B(n498), .Z(G1330GAT) );
  NOR2_X1 U560 ( .A1(n499), .A2(n520), .ZN(n500) );
  XOR2_X1 U561 ( .A(G50GAT), .B(n500), .Z(G1331GAT) );
  XNOR2_X1 U562 ( .A(KEYINPUT105), .B(n544), .ZN(n554) );
  AND2_X1 U563 ( .A1(n362), .A2(n554), .ZN(n510) );
  NAND2_X1 U564 ( .A1(n510), .A2(n501), .ZN(n506) );
  NOR2_X1 U565 ( .A1(n539), .A2(n506), .ZN(n502) );
  XOR2_X1 U566 ( .A(G57GAT), .B(n502), .Z(n503) );
  XNOR2_X1 U567 ( .A(KEYINPUT42), .B(n503), .ZN(G1332GAT) );
  NOR2_X1 U568 ( .A1(n512), .A2(n506), .ZN(n504) );
  XOR2_X1 U569 ( .A(G64GAT), .B(n504), .Z(G1333GAT) );
  NOR2_X1 U570 ( .A1(n524), .A2(n506), .ZN(n505) );
  XOR2_X1 U571 ( .A(G71GAT), .B(n505), .Z(G1334GAT) );
  NOR2_X1 U572 ( .A1(n520), .A2(n506), .ZN(n508) );
  XNOR2_X1 U573 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n507) );
  XNOR2_X1 U574 ( .A(n508), .B(n507), .ZN(G1335GAT) );
  NAND2_X1 U575 ( .A1(n510), .A2(n509), .ZN(n519) );
  NOR2_X1 U576 ( .A1(n539), .A2(n519), .ZN(n511) );
  XOR2_X1 U577 ( .A(G85GAT), .B(n511), .Z(G1336GAT) );
  NOR2_X1 U578 ( .A1(n512), .A2(n519), .ZN(n514) );
  XNOR2_X1 U579 ( .A(KEYINPUT106), .B(KEYINPUT107), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U581 ( .A(G92GAT), .B(n515), .ZN(G1337GAT) );
  NOR2_X1 U582 ( .A1(n524), .A2(n519), .ZN(n516) );
  XOR2_X1 U583 ( .A(G99GAT), .B(n516), .Z(G1338GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n518) );
  XNOR2_X1 U585 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n517) );
  XNOR2_X1 U586 ( .A(n518), .B(n517), .ZN(n522) );
  NOR2_X1 U587 ( .A1(n520), .A2(n519), .ZN(n521) );
  XOR2_X1 U588 ( .A(n522), .B(n521), .Z(G1339GAT) );
  NOR2_X1 U589 ( .A1(n524), .A2(n523), .ZN(n526) );
  NAND2_X1 U590 ( .A1(n526), .A2(n525), .ZN(n528) );
  NOR2_X1 U591 ( .A1(n362), .A2(n528), .ZN(n527) );
  XOR2_X1 U592 ( .A(G113GAT), .B(n527), .Z(G1340GAT) );
  XOR2_X1 U593 ( .A(G120GAT), .B(KEYINPUT115), .Z(n530) );
  INV_X1 U594 ( .A(n528), .ZN(n535) );
  NAND2_X1 U595 ( .A1(n535), .A2(n554), .ZN(n529) );
  XNOR2_X1 U596 ( .A(n530), .B(n529), .ZN(n532) );
  XOR2_X1 U597 ( .A(KEYINPUT114), .B(KEYINPUT49), .Z(n531) );
  XNOR2_X1 U598 ( .A(n532), .B(n531), .ZN(G1341GAT) );
  NAND2_X1 U599 ( .A1(n578), .A2(n535), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n533), .B(KEYINPUT50), .ZN(n534) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(n534), .ZN(G1342GAT) );
  XOR2_X1 U602 ( .A(G134GAT), .B(KEYINPUT51), .Z(n537) );
  NAND2_X1 U603 ( .A1(n535), .A2(n561), .ZN(n536) );
  XNOR2_X1 U604 ( .A(n537), .B(n536), .ZN(G1343GAT) );
  NAND2_X1 U605 ( .A1(n538), .A2(n525), .ZN(n540) );
  NOR2_X1 U606 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n541), .B(KEYINPUT116), .ZN(n548) );
  NAND2_X1 U608 ( .A1(n548), .A2(n542), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n543), .B(G141GAT), .ZN(G1344GAT) );
  INV_X1 U610 ( .A(n548), .ZN(n550) );
  NOR2_X1 U611 ( .A1(n550), .A2(n544), .ZN(n546) );
  XNOR2_X1 U612 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U614 ( .A(G148GAT), .B(n547), .ZN(G1345GAT) );
  NAND2_X1 U615 ( .A1(n548), .A2(n578), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n549), .B(G155GAT), .ZN(G1346GAT) );
  XNOR2_X1 U617 ( .A(G162GAT), .B(KEYINPUT117), .ZN(n553) );
  NOR2_X1 U618 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(G1347GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n556) );
  NAND2_X1 U621 ( .A1(n554), .A2(n560), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U623 ( .A(G176GAT), .B(n557), .ZN(G1349GAT) );
  XOR2_X1 U624 ( .A(G183GAT), .B(KEYINPUT121), .Z(n559) );
  NAND2_X1 U625 ( .A1(n560), .A2(n578), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(G1350GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(KEYINPUT58), .ZN(n563) );
  XNOR2_X1 U629 ( .A(G190GAT), .B(n563), .ZN(G1351GAT) );
  INV_X1 U630 ( .A(KEYINPUT122), .ZN(n569) );
  NOR2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  NAND2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U633 ( .A(n569), .B(n568), .Z(n583) );
  NOR2_X1 U634 ( .A1(n362), .A2(n583), .ZN(n573) );
  XOR2_X1 U635 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n571) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT123), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1352GAT) );
  INV_X1 U639 ( .A(n583), .ZN(n579) );
  NAND2_X1 U640 ( .A1(n579), .A2(n574), .ZN(n576) );
  XOR2_X1 U641 ( .A(KEYINPUT61), .B(KEYINPUT124), .Z(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(G204GAT), .B(n577), .ZN(G1353GAT) );
  XOR2_X1 U644 ( .A(G211GAT), .B(KEYINPUT125), .Z(n581) );
  NAND2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1354GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n585) );
  XNOR2_X1 U648 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(n586) );
  XOR2_X1 U650 ( .A(G218GAT), .B(n586), .Z(G1355GAT) );
endmodule

