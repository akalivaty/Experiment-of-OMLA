

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791;

  NOR2_X1 U374 ( .A1(G953), .A2(G237), .ZN(n534) );
  XNOR2_X1 U375 ( .A(n482), .B(n473), .ZN(n777) );
  XNOR2_X1 U376 ( .A(n582), .B(n581), .ZN(n587) );
  XNOR2_X1 U377 ( .A(n371), .B(KEYINPUT40), .ZN(n791) );
  NOR2_X1 U378 ( .A1(n645), .A2(n447), .ZN(n751) );
  NOR2_X2 U379 ( .A1(n355), .A2(n662), .ZN(n705) );
  XNOR2_X2 U380 ( .A(n634), .B(KEYINPUT19), .ZN(n447) );
  XNOR2_X2 U381 ( .A(n572), .B(n571), .ZN(n634) );
  NAND2_X1 U382 ( .A1(n751), .A2(n727), .ZN(n632) );
  XNOR2_X1 U383 ( .A(n380), .B(KEYINPUT82), .ZN(n379) );
  NAND2_X1 U384 ( .A1(n601), .A2(n600), .ZN(n464) );
  AND2_X1 U385 ( .A1(n466), .A2(n623), .ZN(n606) );
  OR2_X1 U386 ( .A1(n632), .A2(n430), .ZN(n429) );
  NAND2_X1 U387 ( .A1(n379), .A2(n358), .ZN(n378) );
  INV_X1 U388 ( .A(n660), .ZN(n764) );
  NAND2_X1 U389 ( .A1(n407), .A2(n406), .ZN(n394) );
  XNOR2_X1 U390 ( .A(n609), .B(KEYINPUT102), .ZN(n742) );
  AND2_X1 U391 ( .A1(n789), .A2(n633), .ZN(n437) );
  XNOR2_X1 U392 ( .A(n631), .B(n630), .ZN(n789) );
  XNOR2_X1 U393 ( .A(n372), .B(KEYINPUT39), .ZN(n652) );
  NAND2_X1 U394 ( .A1(n643), .A2(n724), .ZN(n372) );
  OR2_X1 U395 ( .A1(n591), .A2(n401), .ZN(n397) );
  NOR2_X1 U396 ( .A1(n619), .A2(n710), .ZN(n623) );
  NAND2_X1 U397 ( .A1(n426), .A2(n357), .ZN(n710) );
  XNOR2_X1 U398 ( .A(n642), .B(KEYINPUT38), .ZN(n724) );
  XNOR2_X1 U399 ( .A(n607), .B(KEYINPUT6), .ZN(n596) );
  BUF_X1 U400 ( .A(n569), .Z(n642) );
  INV_X1 U401 ( .A(n590), .ZN(n426) );
  XNOR2_X1 U402 ( .A(n451), .B(n567), .ZN(n569) );
  XNOR2_X1 U403 ( .A(n543), .B(n542), .ZN(n683) );
  XNOR2_X1 U404 ( .A(n373), .B(n477), .ZN(n700) );
  XNOR2_X1 U405 ( .A(n474), .B(n389), .ZN(n475) );
  XNOR2_X1 U406 ( .A(n480), .B(n428), .ZN(n427) );
  XNOR2_X1 U407 ( .A(n555), .B(n472), .ZN(n482) );
  XNOR2_X1 U408 ( .A(n490), .B(G125), .ZN(n553) );
  INV_X1 U409 ( .A(KEYINPUT3), .ZN(n528) );
  INV_X1 U410 ( .A(G953), .ZN(n550) );
  AND2_X2 U411 ( .A1(n384), .A2(n383), .ZN(n696) );
  NAND2_X1 U412 ( .A1(n764), .A2(n353), .ZN(n352) );
  AND2_X1 U413 ( .A1(n661), .A2(n657), .ZN(n353) );
  XNOR2_X1 U414 ( .A(n609), .B(KEYINPUT102), .ZN(n354) );
  BUF_X1 U415 ( .A(n660), .Z(n355) );
  BUF_X1 U416 ( .A(n777), .Z(n356) );
  XNOR2_X1 U417 ( .A(n543), .B(n475), .ZN(n373) );
  OR2_X1 U418 ( .A1(n759), .A2(n424), .ZN(n422) );
  XNOR2_X1 U419 ( .A(n435), .B(KEYINPUT74), .ZN(n453) );
  AND2_X1 U420 ( .A1(n722), .A2(KEYINPUT34), .ZN(n413) );
  INV_X1 U421 ( .A(KEYINPUT45), .ZN(n441) );
  NAND2_X1 U422 ( .A1(n779), .A2(KEYINPUT2), .ZN(n662) );
  NOR2_X1 U423 ( .A1(n450), .A2(KEYINPUT34), .ZN(n414) );
  NAND2_X1 U424 ( .A1(n422), .A2(n420), .ZN(n419) );
  NAND2_X1 U425 ( .A1(n421), .A2(n615), .ZN(n420) );
  INV_X1 U426 ( .A(n394), .ZN(n392) );
  XNOR2_X1 U427 ( .A(n425), .B(n367), .ZN(n462) );
  NOR2_X1 U428 ( .A1(n453), .A2(n641), .ZN(n650) );
  NAND2_X1 U429 ( .A1(n462), .A2(n458), .ZN(n457) );
  NOR2_X1 U430 ( .A1(n651), .A2(n459), .ZN(n458) );
  INV_X1 U431 ( .A(KEYINPUT83), .ZN(n459) );
  INV_X1 U432 ( .A(G237), .ZN(n546) );
  NAND2_X1 U433 ( .A1(n463), .A2(n465), .ZN(n444) );
  NAND2_X1 U434 ( .A1(n464), .A2(KEYINPUT64), .ZN(n463) );
  NOR2_X1 U435 ( .A1(n394), .A2(n391), .ZN(n465) );
  XNOR2_X1 U436 ( .A(n467), .B(n553), .ZN(n505) );
  XNOR2_X1 U437 ( .A(n390), .B(n389), .ZN(n467) );
  XNOR2_X1 U438 ( .A(KEYINPUT66), .B(KEYINPUT10), .ZN(n390) );
  XNOR2_X1 U439 ( .A(G131), .B(KEYINPUT4), .ZN(n473) );
  XNOR2_X1 U440 ( .A(n518), .B(n517), .ZN(n590) );
  XOR2_X1 U441 ( .A(G119), .B(KEYINPUT97), .Z(n507) );
  XNOR2_X1 U442 ( .A(n505), .B(n504), .ZN(n778) );
  OR2_X1 U443 ( .A1(n376), .A2(n705), .ZN(n375) );
  AND2_X1 U444 ( .A1(n440), .A2(n366), .ZN(n404) );
  NAND2_X1 U445 ( .A1(n413), .A2(n405), .ZN(n408) );
  INV_X1 U446 ( .A(KEYINPUT76), .ZN(n625) );
  XNOR2_X1 U447 ( .A(n439), .B(n438), .ZN(n614) );
  XNOR2_X1 U448 ( .A(G478), .B(KEYINPUT109), .ZN(n438) );
  OR2_X1 U449 ( .A1(n691), .A2(G902), .ZN(n439) );
  NAND2_X1 U450 ( .A1(n434), .A2(KEYINPUT47), .ZN(n432) );
  NAND2_X1 U451 ( .A1(n632), .A2(n434), .ZN(n433) );
  INV_X1 U452 ( .A(KEYINPUT75), .ZN(n434) );
  NAND2_X1 U453 ( .A1(n431), .A2(KEYINPUT75), .ZN(n430) );
  INV_X1 U454 ( .A(KEYINPUT47), .ZN(n431) );
  NAND2_X1 U455 ( .A1(n727), .A2(KEYINPUT110), .ZN(n424) );
  NOR2_X1 U456 ( .A1(n710), .A2(KEYINPUT112), .ZN(n401) );
  XNOR2_X1 U457 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U458 ( .A(G137), .B(G101), .ZN(n538) );
  XOR2_X1 U459 ( .A(KEYINPUT100), .B(KEYINPUT5), .Z(n536) );
  NOR2_X2 U460 ( .A1(n454), .A2(n460), .ZN(n661) );
  NAND2_X1 U461 ( .A1(n457), .A2(n455), .ZN(n454) );
  NOR2_X1 U462 ( .A1(n456), .A2(n788), .ZN(n455) );
  XNOR2_X1 U463 ( .A(G104), .B(G131), .ZN(n491) );
  XOR2_X1 U464 ( .A(G113), .B(G143), .Z(n492) );
  XNOR2_X1 U465 ( .A(KEYINPUT92), .B(KEYINPUT4), .ZN(n556) );
  NOR2_X1 U466 ( .A1(n402), .A2(n399), .ZN(n398) );
  AND2_X1 U467 ( .A1(n590), .A2(n469), .ZN(n618) );
  AND2_X1 U468 ( .A1(n712), .A2(n470), .ZN(n469) );
  NAND2_X1 U469 ( .A1(n700), .A2(n547), .ZN(n479) );
  XNOR2_X1 U470 ( .A(G107), .B(G116), .ZN(n483) );
  INV_X1 U471 ( .A(G134), .ZN(n472) );
  XOR2_X1 U472 ( .A(KEYINPUT107), .B(KEYINPUT7), .Z(n485) );
  NAND2_X1 U473 ( .A1(n587), .A2(n591), .ZN(n597) );
  XNOR2_X1 U474 ( .A(n778), .B(n512), .ZN(n663) );
  NAND2_X1 U475 ( .A1(n386), .A2(n385), .ZN(n384) );
  XOR2_X1 U476 ( .A(KEYINPUT90), .B(n665), .Z(n694) );
  NAND2_X1 U477 ( .A1(n374), .A2(n360), .ZN(n380) );
  OR2_X1 U478 ( .A1(n738), .A2(n645), .ZN(n646) );
  NAND2_X1 U479 ( .A1(n412), .A2(KEYINPUT35), .ZN(n406) );
  NAND2_X1 U480 ( .A1(n409), .A2(n408), .ZN(n407) );
  INV_X1 U481 ( .A(n718), .ZN(n449) );
  INV_X1 U482 ( .A(KEYINPUT113), .ZN(n630) );
  XOR2_X1 U483 ( .A(n712), .B(n577), .Z(n357) );
  AND2_X1 U484 ( .A1(n741), .A2(n740), .ZN(n358) );
  INV_X1 U485 ( .A(n651), .ZN(n461) );
  XOR2_X1 U486 ( .A(KEYINPUT96), .B(KEYINPUT24), .Z(n359) );
  XOR2_X1 U487 ( .A(n709), .B(KEYINPUT80), .Z(n360) );
  XOR2_X1 U488 ( .A(n468), .B(KEYINPUT28), .Z(n361) );
  AND2_X1 U489 ( .A1(n433), .A2(n432), .ZN(n362) );
  AND2_X1 U490 ( .A1(n613), .A2(n614), .ZN(n363) );
  INV_X1 U491 ( .A(G140), .ZN(n389) );
  AND2_X1 U492 ( .A1(n440), .A2(n628), .ZN(n364) );
  AND2_X1 U493 ( .A1(n578), .A2(n357), .ZN(n365) );
  AND2_X1 U494 ( .A1(n628), .A2(n405), .ZN(n366) );
  INV_X1 U495 ( .A(KEYINPUT112), .ZN(n403) );
  XOR2_X1 U496 ( .A(KEYINPUT48), .B(KEYINPUT84), .Z(n367) );
  XNOR2_X1 U497 ( .A(G902), .B(KEYINPUT15), .ZN(n654) );
  OR2_X1 U498 ( .A1(n602), .A2(KEYINPUT44), .ZN(n368) );
  INV_X1 U499 ( .A(KEYINPUT44), .ZN(n391) );
  OR2_X1 U500 ( .A1(n706), .A2(KEYINPUT2), .ZN(n369) );
  OR2_X1 U501 ( .A1(n707), .A2(KEYINPUT79), .ZN(n370) );
  NAND2_X1 U502 ( .A1(n375), .A2(n369), .ZN(n374) );
  NAND2_X1 U503 ( .A1(n352), .A2(n707), .ZN(n381) );
  NAND2_X1 U504 ( .A1(n652), .A2(n363), .ZN(n371) );
  XNOR2_X2 U505 ( .A(n777), .B(G146), .ZN(n543) );
  AND2_X1 U506 ( .A1(n355), .A2(n370), .ZN(n376) );
  XNOR2_X1 U507 ( .A(n378), .B(n377), .ZN(G75) );
  INV_X1 U508 ( .A(KEYINPUT53), .ZN(n377) );
  INV_X1 U509 ( .A(n705), .ZN(n383) );
  NAND2_X1 U510 ( .A1(n381), .A2(n655), .ZN(n386) );
  NOR2_X1 U511 ( .A1(n617), .A2(n616), .ZN(n382) );
  AND2_X1 U512 ( .A1(n382), .A2(n446), .ZN(n445) );
  INV_X1 U513 ( .A(n659), .ZN(n385) );
  NOR2_X1 U514 ( .A1(n423), .A2(n419), .ZN(n418) );
  XNOR2_X1 U515 ( .A(n509), .B(n387), .ZN(n511) );
  XNOR2_X1 U516 ( .A(n508), .B(n359), .ZN(n387) );
  INV_X1 U517 ( .A(n464), .ZN(n448) );
  XNOR2_X1 U518 ( .A(n388), .B(KEYINPUT30), .ZN(n622) );
  NAND2_X1 U519 ( .A1(n715), .A2(n723), .ZN(n388) );
  NAND2_X1 U520 ( .A1(n392), .A2(n391), .ZN(n603) );
  XNOR2_X1 U521 ( .A(n394), .B(n393), .ZN(G24) );
  INV_X1 U522 ( .A(G122), .ZN(n393) );
  NAND2_X1 U523 ( .A1(n395), .A2(n404), .ZN(n411) );
  NAND2_X1 U524 ( .A1(n364), .A2(n395), .ZN(n412) );
  NAND2_X1 U525 ( .A1(n415), .A2(n414), .ZN(n395) );
  NAND2_X1 U526 ( .A1(n397), .A2(n396), .ZN(n400) );
  NAND2_X1 U527 ( .A1(n591), .A2(n403), .ZN(n396) );
  NOR2_X1 U528 ( .A1(n591), .A2(n710), .ZN(n610) );
  NAND2_X1 U529 ( .A1(n400), .A2(n398), .ZN(n594) );
  AND2_X1 U530 ( .A1(n710), .A2(KEYINPUT112), .ZN(n399) );
  INV_X1 U531 ( .A(n596), .ZN(n402) );
  XNOR2_X2 U532 ( .A(n619), .B(KEYINPUT1), .ZN(n591) );
  INV_X1 U533 ( .A(KEYINPUT35), .ZN(n405) );
  NAND2_X1 U534 ( .A1(n411), .A2(n410), .ZN(n409) );
  INV_X1 U535 ( .A(n413), .ZN(n410) );
  INV_X1 U536 ( .A(n722), .ZN(n415) );
  NAND2_X1 U537 ( .A1(n416), .A2(n418), .ZN(n617) );
  NAND2_X1 U538 ( .A1(n354), .A2(n417), .ZN(n416) );
  AND2_X1 U539 ( .A1(n759), .A2(n615), .ZN(n417) );
  INV_X1 U540 ( .A(n727), .ZN(n421) );
  NOR2_X1 U541 ( .A1(n742), .A2(n424), .ZN(n423) );
  NAND2_X1 U542 ( .A1(n649), .A2(n650), .ZN(n425) );
  NAND2_X1 U543 ( .A1(n444), .A2(n368), .ZN(n443) );
  NAND2_X1 U544 ( .A1(n445), .A2(n443), .ZN(n442) );
  NAND2_X1 U545 ( .A1(n466), .A2(n365), .ZN(n582) );
  XNOR2_X2 U546 ( .A(n576), .B(KEYINPUT0), .ZN(n466) );
  NAND2_X1 U547 ( .A1(n427), .A2(G217), .ZN(n481) );
  NAND2_X1 U548 ( .A1(n427), .A2(G221), .ZN(n510) );
  INV_X1 U549 ( .A(KEYINPUT8), .ZN(n428) );
  NAND2_X1 U550 ( .A1(n362), .A2(n429), .ZN(n436) );
  NAND2_X1 U551 ( .A1(n437), .A2(n436), .ZN(n435) );
  XNOR2_X2 U552 ( .A(n479), .B(n478), .ZN(n619) );
  NAND2_X1 U553 ( .A1(n450), .A2(KEYINPUT34), .ZN(n440) );
  XNOR2_X2 U554 ( .A(n594), .B(n593), .ZN(n722) );
  XNOR2_X2 U555 ( .A(n442), .B(n441), .ZN(n660) );
  NAND2_X1 U556 ( .A1(n604), .A2(n448), .ZN(n446) );
  NOR2_X2 U557 ( .A1(n447), .A2(n575), .ZN(n576) );
  AND2_X1 U558 ( .A1(n466), .A2(n449), .ZN(n612) );
  INV_X1 U559 ( .A(n466), .ZN(n450) );
  NAND2_X1 U560 ( .A1(n668), .A2(n654), .ZN(n451) );
  XNOR2_X1 U561 ( .A(n452), .B(n770), .ZN(n668) );
  XNOR2_X2 U562 ( .A(n563), .B(n562), .ZN(n770) );
  XNOR2_X1 U563 ( .A(n559), .B(n560), .ZN(n452) );
  NOR2_X1 U564 ( .A1(n461), .A2(KEYINPUT83), .ZN(n456) );
  NOR2_X1 U565 ( .A1(n462), .A2(KEYINPUT83), .ZN(n460) );
  NAND2_X1 U566 ( .A1(n618), .A2(n715), .ZN(n468) );
  INV_X1 U567 ( .A(n621), .ZN(n470) );
  XNOR2_X2 U568 ( .A(n471), .B(n476), .ZN(n769) );
  XOR2_X2 U569 ( .A(G101), .B(G104), .Z(n471) );
  INV_X1 U570 ( .A(KEYINPUT110), .ZN(n615) );
  XNOR2_X1 U571 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U572 ( .A(n540), .B(n539), .ZN(n541) );
  BUF_X1 U573 ( .A(n668), .Z(n671) );
  XNOR2_X2 U574 ( .A(G143), .B(G128), .ZN(n555) );
  BUF_X2 U575 ( .A(n550), .Z(n780) );
  NAND2_X1 U576 ( .A1(G227), .A2(n780), .ZN(n474) );
  XNOR2_X1 U577 ( .A(G110), .B(G107), .ZN(n476) );
  XNOR2_X1 U578 ( .A(n769), .B(KEYINPUT71), .ZN(n560) );
  XOR2_X1 U579 ( .A(KEYINPUT67), .B(G137), .Z(n504) );
  XNOR2_X1 U580 ( .A(n560), .B(n504), .ZN(n477) );
  INV_X1 U581 ( .A(G902), .ZN(n547) );
  XOR2_X1 U582 ( .A(KEYINPUT68), .B(G469), .Z(n478) );
  INV_X1 U583 ( .A(n591), .ZN(n586) );
  NAND2_X1 U584 ( .A1(G234), .A2(n780), .ZN(n480) );
  XNOR2_X1 U585 ( .A(n482), .B(n481), .ZN(n489) );
  XNOR2_X1 U586 ( .A(n483), .B(KEYINPUT108), .ZN(n487) );
  XNOR2_X1 U587 ( .A(G122), .B(KEYINPUT9), .ZN(n484) );
  XNOR2_X1 U588 ( .A(n485), .B(n484), .ZN(n486) );
  XOR2_X1 U589 ( .A(n487), .B(n486), .Z(n488) );
  XNOR2_X1 U590 ( .A(n489), .B(n488), .ZN(n691) );
  INV_X1 U591 ( .A(G146), .ZN(n490) );
  XNOR2_X1 U592 ( .A(n492), .B(n491), .ZN(n496) );
  XOR2_X1 U593 ( .A(KEYINPUT104), .B(KEYINPUT12), .Z(n494) );
  XNOR2_X1 U594 ( .A(G122), .B(KEYINPUT11), .ZN(n493) );
  XNOR2_X1 U595 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U596 ( .A(n496), .B(n495), .ZN(n500) );
  XOR2_X1 U597 ( .A(KEYINPUT106), .B(KEYINPUT105), .Z(n498) );
  NAND2_X1 U598 ( .A1(n534), .A2(G214), .ZN(n497) );
  XNOR2_X1 U599 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U600 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U601 ( .A(n505), .B(n501), .ZN(n677) );
  NAND2_X1 U602 ( .A1(n677), .A2(n547), .ZN(n503) );
  XNOR2_X1 U603 ( .A(KEYINPUT13), .B(G475), .ZN(n502) );
  XNOR2_X1 U604 ( .A(n503), .B(n502), .ZN(n595) );
  INV_X1 U605 ( .A(n595), .ZN(n613) );
  INV_X1 U606 ( .A(n363), .ZN(n757) );
  XNOR2_X1 U607 ( .A(G110), .B(G128), .ZN(n506) );
  XNOR2_X1 U608 ( .A(n507), .B(n506), .ZN(n509) );
  XOR2_X1 U609 ( .A(KEYINPUT23), .B(KEYINPUT95), .Z(n508) );
  XNOR2_X1 U610 ( .A(n511), .B(n510), .ZN(n512) );
  NAND2_X1 U611 ( .A1(n663), .A2(n547), .ZN(n518) );
  NAND2_X1 U612 ( .A1(n654), .A2(G234), .ZN(n513) );
  XNOR2_X1 U613 ( .A(n513), .B(KEYINPUT20), .ZN(n519) );
  NAND2_X1 U614 ( .A1(G217), .A2(n519), .ZN(n516) );
  INV_X1 U615 ( .A(KEYINPUT77), .ZN(n514) );
  XNOR2_X1 U616 ( .A(n514), .B(KEYINPUT25), .ZN(n515) );
  XNOR2_X1 U617 ( .A(n516), .B(n515), .ZN(n517) );
  NAND2_X1 U618 ( .A1(G221), .A2(n519), .ZN(n521) );
  INV_X1 U619 ( .A(KEYINPUT21), .ZN(n520) );
  XNOR2_X1 U620 ( .A(n521), .B(n520), .ZN(n712) );
  NAND2_X1 U621 ( .A1(G237), .A2(G234), .ZN(n522) );
  XNOR2_X1 U622 ( .A(n522), .B(KEYINPUT14), .ZN(n735) );
  INV_X1 U623 ( .A(G952), .ZN(n523) );
  NAND2_X1 U624 ( .A1(n780), .A2(n523), .ZN(n525) );
  OR2_X1 U625 ( .A1(n780), .A2(G902), .ZN(n524) );
  AND2_X1 U626 ( .A1(n525), .A2(n524), .ZN(n526) );
  AND2_X1 U627 ( .A1(n735), .A2(n526), .ZN(n574) );
  NAND2_X1 U628 ( .A1(G953), .A2(G900), .ZN(n527) );
  NAND2_X1 U629 ( .A1(n574), .A2(n527), .ZN(n621) );
  XNOR2_X1 U630 ( .A(n528), .B(G119), .ZN(n530) );
  XNOR2_X1 U631 ( .A(KEYINPUT69), .B(KEYINPUT70), .ZN(n529) );
  XNOR2_X1 U632 ( .A(n530), .B(n529), .ZN(n533) );
  XNOR2_X1 U633 ( .A(G116), .B(G113), .ZN(n531) );
  XNOR2_X1 U634 ( .A(n531), .B(KEYINPUT91), .ZN(n532) );
  XNOR2_X1 U635 ( .A(n533), .B(n532), .ZN(n561) );
  NAND2_X1 U636 ( .A1(n534), .A2(G210), .ZN(n535) );
  XNOR2_X1 U637 ( .A(n536), .B(n535), .ZN(n540) );
  INV_X1 U638 ( .A(KEYINPUT101), .ZN(n537) );
  XNOR2_X1 U639 ( .A(n561), .B(n541), .ZN(n542) );
  NAND2_X1 U640 ( .A1(n683), .A2(n547), .ZN(n544) );
  XNOR2_X2 U641 ( .A(n544), .B(G472), .ZN(n715) );
  INV_X1 U642 ( .A(n715), .ZN(n607) );
  NAND2_X1 U643 ( .A1(n618), .A2(n596), .ZN(n545) );
  NOR2_X1 U644 ( .A1(n757), .A2(n545), .ZN(n635) );
  NAND2_X1 U645 ( .A1(n547), .A2(n546), .ZN(n564) );
  NAND2_X1 U646 ( .A1(n564), .A2(G214), .ZN(n723) );
  NAND2_X1 U647 ( .A1(n635), .A2(n723), .ZN(n548) );
  NOR2_X1 U648 ( .A1(n586), .A2(n548), .ZN(n549) );
  XNOR2_X1 U649 ( .A(n549), .B(KEYINPUT43), .ZN(n568) );
  XNOR2_X2 U650 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n552) );
  NAND2_X1 U651 ( .A1(n550), .A2(G224), .ZN(n551) );
  XNOR2_X1 U652 ( .A(n552), .B(n551), .ZN(n554) );
  XNOR2_X1 U653 ( .A(n554), .B(n553), .ZN(n558) );
  XNOR2_X1 U654 ( .A(n555), .B(n556), .ZN(n557) );
  XNOR2_X1 U655 ( .A(n558), .B(n557), .ZN(n559) );
  INV_X1 U656 ( .A(n561), .ZN(n563) );
  XNOR2_X1 U657 ( .A(KEYINPUT16), .B(G122), .ZN(n562) );
  NAND2_X1 U658 ( .A1(n564), .A2(G210), .ZN(n566) );
  INV_X1 U659 ( .A(KEYINPUT93), .ZN(n565) );
  INV_X1 U660 ( .A(n642), .ZN(n627) );
  NOR2_X1 U661 ( .A1(n568), .A2(n627), .ZN(n651) );
  XOR2_X1 U662 ( .A(G140), .B(n651), .Z(G42) );
  INV_X1 U663 ( .A(n569), .ZN(n570) );
  NAND2_X1 U664 ( .A1(n570), .A2(n723), .ZN(n572) );
  INV_X1 U665 ( .A(KEYINPUT86), .ZN(n571) );
  XNOR2_X1 U666 ( .A(KEYINPUT94), .B(G898), .ZN(n771) );
  NAND2_X1 U667 ( .A1(n771), .A2(G953), .ZN(n573) );
  NAND2_X1 U668 ( .A1(n574), .A2(n573), .ZN(n575) );
  NAND2_X1 U669 ( .A1(n614), .A2(n595), .ZN(n726) );
  INV_X1 U670 ( .A(n726), .ZN(n578) );
  INV_X1 U671 ( .A(KEYINPUT98), .ZN(n577) );
  XNOR2_X1 U672 ( .A(KEYINPUT73), .B(KEYINPUT22), .ZN(n580) );
  INV_X1 U673 ( .A(KEYINPUT65), .ZN(n579) );
  XNOR2_X1 U674 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U675 ( .A(n591), .B(KEYINPUT88), .ZN(n638) );
  OR2_X1 U676 ( .A1(n596), .A2(n426), .ZN(n583) );
  NOR2_X1 U677 ( .A1(n638), .A2(n583), .ZN(n584) );
  NAND2_X1 U678 ( .A1(n587), .A2(n584), .ZN(n585) );
  XNOR2_X1 U679 ( .A(n585), .B(KEYINPUT32), .ZN(n600) );
  XNOR2_X1 U680 ( .A(n600), .B(G119), .ZN(G21) );
  XNOR2_X1 U681 ( .A(n597), .B(KEYINPUT111), .ZN(n589) );
  AND2_X1 U682 ( .A1(n590), .A2(n607), .ZN(n588) );
  NAND2_X1 U683 ( .A1(n589), .A2(n588), .ZN(n601) );
  XNOR2_X1 U684 ( .A(n601), .B(G110), .ZN(G12) );
  XNOR2_X1 U685 ( .A(KEYINPUT87), .B(KEYINPUT33), .ZN(n592) );
  XNOR2_X1 U686 ( .A(n592), .B(KEYINPUT72), .ZN(n593) );
  NOR2_X1 U687 ( .A1(n614), .A2(n595), .ZN(n628) );
  NOR2_X1 U688 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U689 ( .A(n598), .B(KEYINPUT85), .ZN(n599) );
  NOR2_X1 U690 ( .A1(n599), .A2(n590), .ZN(n616) );
  XOR2_X1 U691 ( .A(G101), .B(n616), .Z(G3) );
  INV_X1 U692 ( .A(KEYINPUT64), .ZN(n602) );
  NAND2_X1 U693 ( .A1(n603), .A2(KEYINPUT64), .ZN(n604) );
  INV_X1 U694 ( .A(KEYINPUT99), .ZN(n605) );
  XNOR2_X1 U695 ( .A(n606), .B(n605), .ZN(n608) );
  NAND2_X1 U696 ( .A1(n608), .A2(n607), .ZN(n609) );
  NAND2_X1 U697 ( .A1(n715), .A2(n610), .ZN(n718) );
  XOR2_X1 U698 ( .A(KEYINPUT31), .B(KEYINPUT103), .Z(n611) );
  XNOR2_X1 U699 ( .A(n612), .B(n611), .ZN(n759) );
  NOR2_X1 U700 ( .A1(n614), .A2(n613), .ZN(n752) );
  INV_X1 U701 ( .A(n752), .ZN(n760) );
  NAND2_X1 U702 ( .A1(n760), .A2(n757), .ZN(n727) );
  INV_X1 U703 ( .A(n619), .ZN(n620) );
  NAND2_X1 U704 ( .A1(n361), .A2(n620), .ZN(n645) );
  NOR2_X1 U705 ( .A1(n622), .A2(n621), .ZN(n624) );
  NAND2_X1 U706 ( .A1(n624), .A2(n623), .ZN(n626) );
  XNOR2_X2 U707 ( .A(n626), .B(n625), .ZN(n643) );
  AND2_X1 U708 ( .A1(n628), .A2(n627), .ZN(n629) );
  NAND2_X1 U709 ( .A1(n643), .A2(n629), .ZN(n631) );
  NAND2_X1 U710 ( .A1(n632), .A2(KEYINPUT47), .ZN(n633) );
  NAND2_X1 U711 ( .A1(n634), .A2(n635), .ZN(n637) );
  XOR2_X1 U712 ( .A(KEYINPUT114), .B(KEYINPUT36), .Z(n636) );
  XNOR2_X1 U713 ( .A(n637), .B(n636), .ZN(n640) );
  INV_X1 U714 ( .A(n638), .ZN(n639) );
  NAND2_X1 U715 ( .A1(n640), .A2(n639), .ZN(n763) );
  INV_X1 U716 ( .A(n763), .ZN(n641) );
  NAND2_X1 U717 ( .A1(n724), .A2(n723), .ZN(n728) );
  NOR2_X1 U718 ( .A1(n728), .A2(n726), .ZN(n644) );
  XNOR2_X1 U719 ( .A(n644), .B(KEYINPUT41), .ZN(n738) );
  XNOR2_X1 U720 ( .A(KEYINPUT42), .B(n646), .ZN(n790) );
  NAND2_X1 U721 ( .A1(n791), .A2(n790), .ZN(n648) );
  INV_X1 U722 ( .A(KEYINPUT46), .ZN(n647) );
  XNOR2_X1 U723 ( .A(n648), .B(n647), .ZN(n649) );
  NAND2_X1 U724 ( .A1(n752), .A2(n652), .ZN(n653) );
  XNOR2_X1 U725 ( .A(n653), .B(KEYINPUT115), .ZN(n788) );
  INV_X1 U726 ( .A(KEYINPUT81), .ZN(n657) );
  INV_X1 U727 ( .A(n654), .ZN(n655) );
  NAND2_X1 U728 ( .A1(n661), .A2(n655), .ZN(n656) );
  NOR2_X1 U729 ( .A1(n660), .A2(n656), .ZN(n658) );
  NOR2_X1 U730 ( .A1(n658), .A2(n657), .ZN(n659) );
  BUF_X2 U731 ( .A(n661), .Z(n779) );
  NAND2_X1 U732 ( .A1(n696), .A2(G217), .ZN(n664) );
  XNOR2_X1 U733 ( .A(n664), .B(n663), .ZN(n666) );
  NOR2_X1 U734 ( .A1(n780), .A2(G952), .ZN(n665) );
  NAND2_X1 U735 ( .A1(n666), .A2(n694), .ZN(n667) );
  XNOR2_X1 U736 ( .A(n667), .B(KEYINPUT125), .ZN(G66) );
  NAND2_X1 U737 ( .A1(n696), .A2(G210), .ZN(n673) );
  XOR2_X1 U738 ( .A(KEYINPUT78), .B(KEYINPUT54), .Z(n669) );
  XNOR2_X1 U739 ( .A(n669), .B(KEYINPUT55), .ZN(n670) );
  XNOR2_X1 U740 ( .A(n671), .B(n670), .ZN(n672) );
  XNOR2_X1 U741 ( .A(n673), .B(n672), .ZN(n674) );
  NAND2_X1 U742 ( .A1(n674), .A2(n694), .ZN(n676) );
  INV_X1 U743 ( .A(KEYINPUT56), .ZN(n675) );
  XNOR2_X1 U744 ( .A(n676), .B(n675), .ZN(G51) );
  NAND2_X1 U745 ( .A1(n696), .A2(G475), .ZN(n679) );
  XOR2_X1 U746 ( .A(KEYINPUT59), .B(n677), .Z(n678) );
  XNOR2_X1 U747 ( .A(n679), .B(n678), .ZN(n680) );
  NAND2_X1 U748 ( .A1(n680), .A2(n694), .ZN(n682) );
  INV_X1 U749 ( .A(KEYINPUT60), .ZN(n681) );
  XNOR2_X1 U750 ( .A(n682), .B(n681), .ZN(G60) );
  NAND2_X1 U751 ( .A1(n696), .A2(G472), .ZN(n685) );
  XNOR2_X1 U752 ( .A(n683), .B(KEYINPUT62), .ZN(n684) );
  XNOR2_X1 U753 ( .A(n685), .B(n684), .ZN(n686) );
  NAND2_X1 U754 ( .A1(n686), .A2(n694), .ZN(n689) );
  XOR2_X1 U755 ( .A(KEYINPUT116), .B(KEYINPUT63), .Z(n687) );
  XNOR2_X1 U756 ( .A(n687), .B(KEYINPUT89), .ZN(n688) );
  XNOR2_X1 U757 ( .A(n689), .B(n688), .ZN(G57) );
  BUF_X1 U758 ( .A(n696), .Z(n690) );
  NAND2_X1 U759 ( .A1(n690), .A2(G478), .ZN(n693) );
  XNOR2_X1 U760 ( .A(n691), .B(KEYINPUT124), .ZN(n692) );
  XNOR2_X1 U761 ( .A(n693), .B(n692), .ZN(n695) );
  INV_X1 U762 ( .A(n694), .ZN(n703) );
  NOR2_X1 U763 ( .A1(n695), .A2(n703), .ZN(G63) );
  NAND2_X1 U764 ( .A1(n690), .A2(G469), .ZN(n702) );
  XOR2_X1 U765 ( .A(KEYINPUT123), .B(KEYINPUT122), .Z(n698) );
  XNOR2_X1 U766 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n697) );
  XNOR2_X1 U767 ( .A(n698), .B(n697), .ZN(n699) );
  XNOR2_X1 U768 ( .A(n700), .B(n699), .ZN(n701) );
  XNOR2_X1 U769 ( .A(n702), .B(n701), .ZN(n704) );
  NOR2_X1 U770 ( .A1(n704), .A2(n703), .ZN(G54) );
  INV_X1 U771 ( .A(KEYINPUT2), .ZN(n707) );
  INV_X1 U772 ( .A(KEYINPUT79), .ZN(n706) );
  XNOR2_X1 U773 ( .A(KEYINPUT79), .B(n707), .ZN(n708) );
  NOR2_X1 U774 ( .A1(n779), .A2(n708), .ZN(n709) );
  NAND2_X1 U775 ( .A1(n710), .A2(n591), .ZN(n711) );
  XNOR2_X1 U776 ( .A(n711), .B(KEYINPUT50), .ZN(n717) );
  NOR2_X1 U777 ( .A1(n426), .A2(n712), .ZN(n713) );
  XOR2_X1 U778 ( .A(KEYINPUT49), .B(n713), .Z(n714) );
  NOR2_X1 U779 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U780 ( .A1(n717), .A2(n716), .ZN(n719) );
  NAND2_X1 U781 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U782 ( .A(KEYINPUT51), .B(n720), .ZN(n721) );
  NOR2_X1 U783 ( .A1(n738), .A2(n721), .ZN(n733) );
  NOR2_X1 U784 ( .A1(n724), .A2(n723), .ZN(n725) );
  NOR2_X1 U785 ( .A1(n726), .A2(n725), .ZN(n730) );
  NOR2_X1 U786 ( .A1(n421), .A2(n728), .ZN(n729) );
  NOR2_X1 U787 ( .A1(n730), .A2(n729), .ZN(n731) );
  NOR2_X1 U788 ( .A1(n722), .A2(n731), .ZN(n732) );
  NOR2_X1 U789 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U790 ( .A(KEYINPUT52), .B(n734), .ZN(n737) );
  NAND2_X1 U791 ( .A1(G952), .A2(n735), .ZN(n736) );
  OR2_X1 U792 ( .A1(n737), .A2(n736), .ZN(n741) );
  NOR2_X1 U793 ( .A1(n722), .A2(n738), .ZN(n739) );
  NOR2_X1 U794 ( .A1(n739), .A2(G953), .ZN(n740) );
  NOR2_X1 U795 ( .A1(n354), .A2(n757), .ZN(n744) );
  XNOR2_X1 U796 ( .A(G104), .B(KEYINPUT117), .ZN(n743) );
  XNOR2_X1 U797 ( .A(n744), .B(n743), .ZN(G6) );
  XOR2_X1 U798 ( .A(KEYINPUT120), .B(KEYINPUT119), .Z(n746) );
  XNOR2_X1 U799 ( .A(KEYINPUT26), .B(KEYINPUT27), .ZN(n745) );
  XNOR2_X1 U800 ( .A(n746), .B(n745), .ZN(n750) );
  NOR2_X1 U801 ( .A1(n354), .A2(n760), .ZN(n748) );
  XNOR2_X1 U802 ( .A(G107), .B(KEYINPUT118), .ZN(n747) );
  XNOR2_X1 U803 ( .A(n748), .B(n747), .ZN(n749) );
  XNOR2_X1 U804 ( .A(n750), .B(n749), .ZN(G9) );
  XOR2_X1 U805 ( .A(KEYINPUT121), .B(KEYINPUT29), .Z(n754) );
  NAND2_X1 U806 ( .A1(n751), .A2(n752), .ZN(n753) );
  XNOR2_X1 U807 ( .A(n754), .B(n753), .ZN(n755) );
  XOR2_X1 U808 ( .A(G128), .B(n755), .Z(G30) );
  NAND2_X1 U809 ( .A1(n751), .A2(n363), .ZN(n756) );
  XNOR2_X1 U810 ( .A(n756), .B(G146), .ZN(G48) );
  NOR2_X1 U811 ( .A1(n757), .A2(n759), .ZN(n758) );
  XOR2_X1 U812 ( .A(G113), .B(n758), .Z(G15) );
  NOR2_X1 U813 ( .A1(n760), .A2(n759), .ZN(n761) );
  XOR2_X1 U814 ( .A(G116), .B(n761), .Z(G18) );
  XOR2_X1 U815 ( .A(G125), .B(KEYINPUT37), .Z(n762) );
  XNOR2_X1 U816 ( .A(n763), .B(n762), .ZN(G27) );
  NAND2_X1 U817 ( .A1(n764), .A2(n780), .ZN(n768) );
  NAND2_X1 U818 ( .A1(G953), .A2(G224), .ZN(n765) );
  XNOR2_X1 U819 ( .A(n765), .B(KEYINPUT61), .ZN(n766) );
  NAND2_X1 U820 ( .A1(n766), .A2(n771), .ZN(n767) );
  NAND2_X1 U821 ( .A1(n768), .A2(n767), .ZN(n775) );
  XOR2_X1 U822 ( .A(n770), .B(n769), .Z(n773) );
  NOR2_X1 U823 ( .A1(n771), .A2(n780), .ZN(n772) );
  NOR2_X1 U824 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U825 ( .A(n775), .B(n774), .ZN(n776) );
  XNOR2_X1 U826 ( .A(KEYINPUT126), .B(n776), .ZN(G69) );
  XNOR2_X1 U827 ( .A(n356), .B(n778), .ZN(n782) );
  XOR2_X1 U828 ( .A(n782), .B(n779), .Z(n781) );
  NAND2_X1 U829 ( .A1(n781), .A2(n780), .ZN(n787) );
  XNOR2_X1 U830 ( .A(G227), .B(n782), .ZN(n783) );
  NAND2_X1 U831 ( .A1(n783), .A2(G900), .ZN(n784) );
  XOR2_X1 U832 ( .A(KEYINPUT127), .B(n784), .Z(n785) );
  NAND2_X1 U833 ( .A1(G953), .A2(n785), .ZN(n786) );
  NAND2_X1 U834 ( .A1(n787), .A2(n786), .ZN(G72) );
  XOR2_X1 U835 ( .A(G134), .B(n788), .Z(G36) );
  XNOR2_X1 U836 ( .A(G143), .B(n789), .ZN(G45) );
  XNOR2_X1 U837 ( .A(G137), .B(n790), .ZN(G39) );
  XNOR2_X1 U838 ( .A(G131), .B(n791), .ZN(G33) );
endmodule

