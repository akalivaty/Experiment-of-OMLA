//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 1 1 0 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 1 1 0 1 0 1 1 0 0 0 0 1 0 1 0 0 1 0 0 1 1 1 1 1 0 1 1 0 1 0 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:09 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1218, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1281,
    new_n1282, new_n1283, new_n1284;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT0), .Z(new_n208));
  AOI22_X1  g0008(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n209));
  INV_X1    g0009(.A(G87), .ZN(new_n210));
  INV_X1    g0010(.A(G250), .ZN(new_n211));
  OAI21_X1  g0011(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AOI21_X1  g0012(.A(new_n212), .B1(G116), .B2(G270), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G58), .A2(G232), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G107), .A2(G264), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G50), .A2(G226), .ZN(new_n216));
  NAND4_X1  g0016(.A1(new_n213), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  AND2_X1   g0017(.A1(G68), .A2(G238), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n205), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT1), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OR2_X1    g0023(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n224), .A2(G50), .A3(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  AOI211_X1 g0027(.A(new_n208), .B(new_n220), .C1(new_n223), .C2(new_n227), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n232), .B(KEYINPUT65), .Z(new_n233));
  XOR2_X1   g0033(.A(G250), .B(G257), .Z(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G87), .B(G97), .ZN(new_n238));
  INV_X1    g0038(.A(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(KEYINPUT66), .B(G107), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G68), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  INV_X1    g0046(.A(G1), .ZN(new_n247));
  OAI211_X1 g0047(.A(new_n247), .B(G274), .C1(G41), .C2(G45), .ZN(new_n248));
  NAND2_X1  g0048(.A1(G33), .A2(G41), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n249), .A2(G1), .A3(G13), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n247), .B1(G41), .B2(G45), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G226), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n248), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  OR2_X1    g0054(.A1(new_n254), .A2(KEYINPUT67), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT3), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G222), .A2(G1698), .ZN(new_n261));
  INV_X1    g0061(.A(G1698), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(G223), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n260), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n250), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n264), .B(new_n265), .C1(G77), .C2(new_n260), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n254), .A2(KEYINPUT67), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n255), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  OR2_X1    g0068(.A1(new_n268), .A2(G179), .ZN(new_n269));
  OAI21_X1  g0069(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n270));
  INV_X1    g0070(.A(G150), .ZN(new_n271));
  NOR2_X1   g0071(.A1(G20), .A2(G33), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n257), .A2(G20), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT8), .B(G58), .ZN(new_n276));
  OAI221_X1 g0076(.A(new_n270), .B1(new_n271), .B2(new_n273), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n221), .ZN(new_n279));
  INV_X1    g0079(.A(G50), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n247), .A2(G13), .A3(G20), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  AOI22_X1  g0082(.A1(new_n277), .A2(new_n279), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n279), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n247), .A2(G20), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n284), .A2(G50), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G169), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n268), .A2(new_n288), .ZN(new_n289));
  AND3_X1   g0089(.A1(new_n269), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT9), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n292), .B(KEYINPUT70), .ZN(new_n293));
  INV_X1    g0093(.A(G190), .ZN(new_n294));
  OAI22_X1  g0094(.A1(new_n287), .A2(new_n291), .B1(new_n268), .B2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n295), .B1(G200), .B2(new_n268), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(KEYINPUT10), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT10), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n293), .A2(new_n296), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n290), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G58), .ZN(new_n302));
  INV_X1    g0102(.A(G68), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(G20), .B1(new_n304), .B2(new_n201), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n272), .A2(G159), .ZN(new_n306));
  AND3_X1   g0106(.A1(new_n305), .A2(KEYINPUT73), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(KEYINPUT73), .B1(new_n305), .B2(new_n306), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT72), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n258), .A2(new_n222), .A3(new_n259), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT7), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n258), .A2(KEYINPUT7), .A3(new_n222), .A4(new_n259), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n310), .B1(new_n315), .B2(G68), .ZN(new_n316));
  AOI211_X1 g0116(.A(KEYINPUT72), .B(new_n303), .C1(new_n313), .C2(new_n314), .ZN(new_n317));
  OAI211_X1 g0117(.A(KEYINPUT16), .B(new_n309), .C1(new_n316), .C2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT16), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n305), .A2(new_n306), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT73), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n305), .A2(KEYINPUT73), .A3(new_n306), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n303), .B1(new_n313), .B2(new_n314), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n319), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n318), .A2(new_n279), .A3(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n285), .ZN(new_n328));
  NOR3_X1   g0128(.A1(new_n276), .A2(new_n328), .A3(new_n279), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n329), .B1(new_n282), .B2(new_n276), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n250), .A2(G232), .A3(new_n251), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n248), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT74), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G223), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n262), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n253), .A2(G1698), .ZN(new_n337));
  AND2_X1   g0137(.A1(KEYINPUT3), .A2(G33), .ZN(new_n338));
  NOR2_X1   g0138(.A1(KEYINPUT3), .A2(G33), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n336), .B(new_n337), .C1(new_n338), .C2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(G33), .A2(G87), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n265), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n331), .A2(KEYINPUT74), .A3(new_n248), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n334), .A2(new_n343), .A3(new_n294), .A4(new_n344), .ZN(new_n345));
  AND3_X1   g0145(.A1(new_n331), .A2(KEYINPUT74), .A3(new_n248), .ZN(new_n346));
  AOI21_X1  g0146(.A(KEYINPUT74), .B1(new_n331), .B2(new_n248), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n250), .B1(new_n340), .B2(new_n341), .ZN(new_n348));
  NOR3_X1   g0148(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  OAI211_X1 g0149(.A(KEYINPUT75), .B(new_n345), .C1(new_n349), .C2(G200), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n334), .A2(new_n343), .A3(new_n344), .ZN(new_n352));
  INV_X1    g0152(.A(G200), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(KEYINPUT75), .B1(new_n354), .B2(new_n345), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n327), .B(new_n330), .C1(new_n351), .C2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT17), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT75), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n346), .A2(new_n347), .ZN(new_n360));
  AOI21_X1  g0160(.A(G200), .B1(new_n360), .B2(new_n343), .ZN(new_n361));
  INV_X1    g0161(.A(new_n345), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n359), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n350), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n364), .A2(KEYINPUT17), .A3(new_n327), .A4(new_n330), .ZN(new_n365));
  AND2_X1   g0165(.A1(new_n358), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT18), .ZN(new_n367));
  AND2_X1   g0167(.A1(new_n327), .A2(new_n330), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n349), .A2(G179), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n352), .A2(G169), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n367), .B1(new_n368), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n327), .A2(new_n330), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n374), .A2(KEYINPUT18), .A3(new_n371), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n260), .A2(G238), .A3(G1698), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n260), .A2(G232), .A3(new_n262), .ZN(new_n378));
  INV_X1    g0178(.A(G107), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n377), .B(new_n378), .C1(new_n379), .C2(new_n260), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(new_n265), .ZN(new_n381));
  INV_X1    g0181(.A(G244), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n381), .B(new_n248), .C1(new_n382), .C2(new_n252), .ZN(new_n383));
  AND2_X1   g0183(.A1(new_n383), .A2(G200), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n383), .A2(new_n294), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT68), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n281), .A2(new_n386), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n247), .A2(KEYINPUT68), .A3(G13), .A4(G20), .ZN(new_n388));
  AND3_X1   g0188(.A1(new_n284), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n389), .A2(G77), .A3(new_n285), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n387), .A2(new_n388), .ZN(new_n391));
  INV_X1    g0191(.A(G77), .ZN(new_n392));
  AND3_X1   g0192(.A1(new_n391), .A2(KEYINPUT69), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(KEYINPUT69), .B1(new_n391), .B2(new_n392), .ZN(new_n394));
  OAI22_X1  g0194(.A1(new_n276), .A2(new_n273), .B1(new_n222), .B2(new_n392), .ZN(new_n395));
  XOR2_X1   g0195(.A(KEYINPUT15), .B(G87), .Z(new_n396));
  AOI21_X1  g0196(.A(new_n395), .B1(new_n274), .B2(new_n396), .ZN(new_n397));
  OAI221_X1 g0197(.A(new_n390), .B1(new_n393), .B2(new_n394), .C1(new_n397), .C2(new_n284), .ZN(new_n398));
  NOR3_X1   g0198(.A1(new_n384), .A2(new_n385), .A3(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n301), .A2(new_n366), .A3(new_n376), .A4(new_n400), .ZN(new_n401));
  OAI211_X1 g0201(.A(G226), .B(new_n262), .C1(new_n338), .C2(new_n339), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(KEYINPUT71), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT71), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n260), .A2(new_n404), .A3(G226), .A4(new_n262), .ZN(new_n405));
  AND2_X1   g0205(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  OAI211_X1 g0206(.A(G232), .B(G1698), .C1(new_n338), .C2(new_n339), .ZN(new_n407));
  NAND2_X1  g0207(.A1(G33), .A2(G97), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n265), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT13), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n250), .A2(G238), .A3(new_n251), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n410), .A2(new_n411), .A3(new_n248), .A4(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n409), .B1(new_n405), .B2(new_n403), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n248), .B(new_n412), .C1(new_n414), .C2(new_n250), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT13), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(G169), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT14), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n413), .A2(new_n416), .A3(G179), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT14), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n417), .A2(new_n421), .A3(G169), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n419), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(KEYINPUT12), .B1(new_n282), .B2(new_n303), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT12), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n425), .B1(new_n387), .B2(new_n388), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n424), .B1(new_n426), .B2(new_n303), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n389), .A2(G68), .A3(new_n285), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n274), .A2(G77), .B1(G20), .B2(new_n303), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(new_n280), .B2(new_n273), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n279), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n431), .A2(KEYINPUT11), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n431), .A2(KEYINPUT11), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n427), .B(new_n428), .C1(new_n432), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n423), .A2(new_n434), .ZN(new_n435));
  OR2_X1    g0235(.A1(new_n383), .A2(G179), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n383), .A2(new_n288), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n436), .A2(new_n398), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n434), .B1(new_n417), .B2(G200), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n413), .A2(new_n416), .A3(G190), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  NOR3_X1   g0243(.A1(new_n401), .A2(new_n439), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n239), .B1(new_n247), .B2(G33), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n389), .A2(new_n445), .B1(new_n239), .B2(new_n391), .ZN(new_n446));
  AOI21_X1  g0246(.A(G20), .B1(G33), .B2(G283), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n257), .A2(G97), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(KEYINPUT79), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT79), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n447), .A2(new_n448), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  AOI22_X1  g0253(.A1(new_n278), .A2(new_n221), .B1(G20), .B2(new_n239), .ZN(new_n454));
  AOI21_X1  g0254(.A(KEYINPUT20), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AND3_X1   g0255(.A1(new_n447), .A2(new_n448), .A3(new_n451), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n451), .B1(new_n447), .B2(new_n448), .ZN(new_n457));
  OAI211_X1 g0257(.A(KEYINPUT20), .B(new_n454), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n446), .B1(new_n455), .B2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n260), .A2(G264), .A3(G1698), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n260), .A2(G257), .A3(new_n262), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n338), .A2(new_n339), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(G303), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n461), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(new_n265), .ZN(new_n466));
  INV_X1    g0266(.A(G45), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n467), .A2(G1), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(G274), .ZN(new_n469));
  INV_X1    g0269(.A(G41), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(KEYINPUT5), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT5), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(G41), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n474), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n265), .B1(new_n477), .B2(new_n468), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(G270), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n466), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n460), .A2(new_n480), .A3(G169), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT80), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(KEYINPUT21), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT21), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n481), .A2(KEYINPUT80), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n466), .A2(new_n479), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n487), .A2(new_n460), .A3(G179), .A4(new_n476), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n480), .A2(G200), .ZN(new_n489));
  INV_X1    g0289(.A(new_n460), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n489), .B(new_n490), .C1(new_n294), .C2(new_n480), .ZN(new_n491));
  AND4_X1   g0291(.A1(new_n483), .A2(new_n485), .A3(new_n488), .A4(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n468), .ZN(new_n493));
  OAI211_X1 g0293(.A(G264), .B(new_n250), .C1(new_n474), .C2(new_n493), .ZN(new_n494));
  XNOR2_X1  g0294(.A(new_n494), .B(KEYINPUT81), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n260), .A2(G257), .A3(G1698), .ZN(new_n496));
  NAND2_X1  g0296(.A1(G33), .A2(G294), .ZN(new_n497));
  OAI211_X1 g0297(.A(G250), .B(new_n262), .C1(new_n338), .C2(new_n339), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n475), .B1(new_n499), .B2(new_n265), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n495), .A2(G179), .A3(new_n500), .ZN(new_n501));
  AND2_X1   g0301(.A1(new_n500), .A2(new_n494), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n501), .B1(new_n502), .B2(new_n288), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n222), .B(G87), .C1(new_n338), .C2(new_n339), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(KEYINPUT22), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT22), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n260), .A2(new_n506), .A3(new_n222), .A4(G87), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT24), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT23), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n510), .B1(new_n222), .B2(G107), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n379), .A2(KEYINPUT23), .A3(G20), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n511), .A2(new_n512), .B1(new_n274), .B2(G116), .ZN(new_n513));
  AND3_X1   g0313(.A1(new_n508), .A2(new_n509), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n509), .B1(new_n508), .B2(new_n513), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n279), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n247), .A2(G33), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n284), .A2(new_n281), .A3(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT25), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n520), .B1(new_n281), .B2(G107), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n282), .A2(KEYINPUT25), .A3(new_n379), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n519), .A2(G107), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n516), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n503), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(KEYINPUT82), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT82), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n503), .A2(new_n524), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(G200), .B1(new_n495), .B2(new_n500), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n499), .A2(new_n265), .ZN(new_n531));
  AND4_X1   g0331(.A1(new_n294), .A2(new_n531), .A3(new_n476), .A4(new_n494), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n516), .B(new_n523), .C1(new_n530), .C2(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(KEYINPUT7), .B1(new_n463), .B2(new_n222), .ZN(new_n534));
  INV_X1    g0334(.A(new_n314), .ZN(new_n535));
  OAI21_X1  g0335(.A(G107), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT6), .ZN(new_n537));
  AND2_X1   g0337(.A1(G97), .A2(G107), .ZN(new_n538));
  NOR2_X1   g0338(.A1(G97), .A2(G107), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n379), .A2(KEYINPUT6), .A3(G97), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n542), .A2(G20), .B1(G77), .B2(new_n272), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n284), .B1(new_n536), .B2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(G97), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n518), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n281), .A2(G97), .ZN(new_n547));
  NOR3_X1   g0347(.A1(new_n544), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  OAI211_X1 g0348(.A(G244), .B(new_n262), .C1(new_n338), .C2(new_n339), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT4), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n260), .A2(KEYINPUT4), .A3(G244), .A4(new_n262), .ZN(new_n552));
  NAND2_X1  g0352(.A1(G33), .A2(G283), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n260), .A2(G250), .A3(G1698), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n551), .A2(new_n552), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n265), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n475), .B1(new_n478), .B2(G257), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(G200), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n556), .A2(G190), .A3(new_n557), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n548), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n558), .A2(new_n288), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n542), .A2(G20), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n272), .A2(G77), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n379), .B1(new_n313), .B2(new_n314), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n279), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n546), .ZN(new_n568));
  INV_X1    g0368(.A(new_n547), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(G179), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n556), .A2(new_n571), .A3(new_n557), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n562), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n533), .A2(new_n561), .A3(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(G244), .B(G1698), .C1(new_n338), .C2(new_n339), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT76), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n260), .A2(KEYINPUT76), .A3(G244), .A4(G1698), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n260), .A2(G238), .A3(new_n262), .ZN(new_n579));
  NAND2_X1  g0379(.A1(G33), .A2(G116), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n577), .A2(new_n578), .A3(new_n579), .A4(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n265), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n493), .A2(new_n250), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n469), .B1(new_n583), .B2(new_n211), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(G200), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n584), .B1(new_n581), .B2(new_n265), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(G190), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT19), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n222), .B1(new_n408), .B2(new_n590), .ZN(new_n591));
  NOR4_X1   g0391(.A1(KEYINPUT77), .A2(G87), .A3(G97), .A4(G107), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT77), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n593), .B1(new_n539), .B2(new_n210), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n591), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n260), .A2(new_n222), .A3(G68), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n590), .B1(new_n275), .B2(new_n545), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n279), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n519), .A2(G87), .ZN(new_n600));
  INV_X1    g0400(.A(new_n396), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n391), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n599), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n587), .A2(new_n589), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n519), .A2(new_n396), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n599), .A2(new_n602), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(KEYINPUT78), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT78), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n599), .A2(new_n608), .A3(new_n602), .A4(new_n605), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n288), .B1(new_n582), .B2(new_n585), .ZN(new_n611));
  AOI211_X1 g0411(.A(new_n571), .B(new_n584), .C1(new_n581), .C2(new_n265), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n604), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n574), .A2(new_n614), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n444), .A2(new_n492), .A3(new_n529), .A4(new_n615), .ZN(new_n616));
  XNOR2_X1  g0416(.A(new_n616), .B(KEYINPUT83), .ZN(G372));
  OAI21_X1  g0417(.A(new_n606), .B1(new_n611), .B2(new_n612), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n604), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n574), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n483), .A2(new_n485), .A3(new_n488), .ZN(new_n621));
  INV_X1    g0421(.A(new_n525), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n619), .A2(new_n573), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT26), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g0426(.A(new_n618), .B(KEYINPUT84), .Z(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n562), .A2(new_n570), .A3(new_n572), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n629), .B(new_n604), .C1(new_n613), .C2(new_n610), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(KEYINPUT26), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n623), .A2(new_n626), .A3(new_n628), .A4(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n444), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n439), .A2(new_n366), .A3(new_n442), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n376), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n298), .A2(new_n300), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n290), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n633), .A2(new_n637), .ZN(G369));
  XNOR2_X1  g0438(.A(KEYINPUT85), .B(KEYINPUT27), .ZN(new_n639));
  INV_X1    g0439(.A(G13), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n640), .A2(G20), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  OR3_X1    g0442(.A1(new_n639), .A2(new_n642), .A3(G1), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n639), .B1(new_n642), .B2(G1), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(G213), .A3(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(G343), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n492), .B1(new_n490), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n621), .A2(new_n460), .A3(new_n647), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g0451(.A(KEYINPUT86), .B(G330), .Z(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n503), .A2(new_n524), .A3(new_n527), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n527), .B1(new_n503), .B2(new_n524), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n533), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n524), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n659), .B1(new_n660), .B2(new_n648), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n661), .B1(new_n525), .B2(new_n648), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n654), .A2(new_n662), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n621), .A2(new_n648), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n659), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n622), .A2(new_n648), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n663), .A2(new_n668), .ZN(G399));
  INV_X1    g0469(.A(new_n206), .ZN(new_n670));
  OR3_X1    g0470(.A1(new_n670), .A2(KEYINPUT87), .A3(G41), .ZN(new_n671));
  OAI21_X1  g0471(.A(KEYINPUT87), .B1(new_n670), .B2(G41), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n592), .A2(new_n594), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n239), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n673), .A2(new_n676), .A3(G1), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n226), .B2(new_n673), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n678), .B(KEYINPUT28), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n632), .A2(new_n648), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(KEYINPUT29), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n630), .A2(new_n625), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT90), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n624), .A2(KEYINPUT26), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n630), .A2(KEYINPUT90), .A3(new_n625), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n620), .B1(new_n657), .B2(new_n621), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT91), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OAI211_X1 g0490(.A(new_n620), .B(KEYINPUT91), .C1(new_n657), .C2(new_n621), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n687), .A2(new_n690), .A3(new_n628), .A4(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(new_n648), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n681), .B1(new_n693), .B2(KEYINPUT29), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT31), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n558), .A2(new_n486), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n495), .A2(new_n500), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n696), .A2(KEYINPUT30), .A3(new_n697), .A4(new_n612), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(KEYINPUT88), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n495), .A2(new_n500), .ZN(new_n700));
  NOR3_X1   g0500(.A1(new_n700), .A2(new_n558), .A3(new_n486), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT88), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n701), .A2(new_n702), .A3(KEYINPUT30), .A4(new_n612), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n558), .A2(new_n586), .A3(new_n571), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n705), .A2(new_n480), .A3(new_n700), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT30), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n696), .A2(new_n697), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n588), .A2(G179), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  AOI211_X1 g0511(.A(new_n695), .B(new_n648), .C1(new_n707), .C2(new_n711), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n492), .A2(new_n615), .A3(new_n529), .A4(new_n648), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n711), .A2(KEYINPUT89), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT89), .ZN(new_n715));
  OAI211_X1 g0515(.A(new_n715), .B(new_n708), .C1(new_n709), .C2(new_n710), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n714), .A2(new_n704), .A3(new_n706), .A4(new_n716), .ZN(new_n717));
  AOI22_X1  g0517(.A1(new_n713), .A2(KEYINPUT31), .B1(new_n717), .B2(new_n647), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n652), .B1(new_n712), .B2(new_n718), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n694), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n679), .B1(new_n720), .B2(G1), .ZN(G364));
  INV_X1    g0521(.A(new_n673), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n247), .B1(new_n641), .B2(G45), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n654), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n726), .B1(new_n652), .B2(new_n651), .ZN(new_n727));
  INV_X1    g0527(.A(new_n725), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n670), .A2(new_n260), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n730), .B1(new_n245), .B2(G45), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n731), .B1(G45), .B2(new_n226), .ZN(new_n732));
  INV_X1    g0532(.A(G355), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n260), .A2(new_n206), .ZN(new_n734));
  OAI221_X1 g0534(.A(new_n732), .B1(G116), .B2(new_n206), .C1(new_n733), .C2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(G13), .A2(G33), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(G20), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n221), .B1(G20), .B2(new_n288), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n728), .B1(new_n735), .B2(new_n740), .ZN(new_n741));
  XOR2_X1   g0541(.A(new_n741), .B(KEYINPUT92), .Z(new_n742));
  INV_X1    g0542(.A(new_n738), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n222), .A2(new_n294), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n571), .A2(new_n353), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(G326), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n222), .A2(G190), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n571), .A2(G200), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(G311), .ZN(new_n751));
  OAI22_X1  g0551(.A1(new_n746), .A2(new_n747), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(G179), .A2(G200), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n222), .B1(new_n753), .B2(G190), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n752), .B1(G294), .B2(new_n755), .ZN(new_n756));
  XOR2_X1   g0556(.A(new_n756), .B(KEYINPUT93), .Z(new_n757));
  NAND2_X1  g0557(.A1(new_n748), .A2(new_n753), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI211_X1 g0559(.A(new_n260), .B(new_n757), .C1(G329), .C2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n353), .A2(G179), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n748), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G283), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n744), .A2(new_n761), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n744), .A2(new_n749), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI22_X1  g0568(.A1(G303), .A2(new_n766), .B1(new_n768), .B2(G322), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n745), .A2(new_n748), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(KEYINPUT33), .A2(G317), .ZN(new_n772));
  AND2_X1   g0572(.A1(KEYINPUT33), .A2(G317), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n771), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND4_X1  g0574(.A1(new_n760), .A2(new_n764), .A3(new_n769), .A4(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n754), .A2(new_n545), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n303), .A2(new_n770), .B1(new_n765), .B2(new_n210), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n776), .B(new_n777), .C1(G58), .C2(new_n768), .ZN(new_n778));
  INV_X1    g0578(.A(new_n750), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G77), .ZN(new_n780));
  INV_X1    g0580(.A(G159), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n758), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n782), .B(KEYINPUT32), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n762), .A2(new_n379), .ZN(new_n784));
  INV_X1    g0584(.A(new_n746), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n463), .B(new_n784), .C1(G50), .C2(new_n785), .ZN(new_n786));
  NAND4_X1  g0586(.A1(new_n778), .A2(new_n780), .A3(new_n783), .A4(new_n786), .ZN(new_n787));
  AND2_X1   g0587(.A1(new_n775), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n739), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n742), .B1(new_n651), .B2(new_n743), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  AND2_X1   g0590(.A1(new_n727), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(G396));
  INV_X1    g0592(.A(new_n438), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(KEYINPUT94), .ZN(new_n794));
  INV_X1    g0594(.A(KEYINPUT94), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n438), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n399), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n398), .A2(new_n647), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n797), .A2(new_n798), .B1(new_n793), .B2(new_n647), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n680), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n632), .A2(new_n648), .A3(new_n797), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XOR2_X1   g0602(.A(new_n802), .B(new_n719), .Z(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(new_n728), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n799), .A2(new_n736), .ZN(new_n805));
  INV_X1    g0605(.A(G303), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n746), .A2(new_n806), .B1(new_n762), .B2(new_n210), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n260), .B(new_n807), .C1(G283), .C2(new_n771), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n768), .A2(G294), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n759), .A2(G311), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n750), .A2(new_n239), .ZN(new_n811));
  AOI211_X1 g0611(.A(new_n776), .B(new_n811), .C1(G107), .C2(new_n766), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n808), .A2(new_n809), .A3(new_n810), .A4(new_n812), .ZN(new_n813));
  AOI22_X1  g0613(.A1(G143), .A2(new_n768), .B1(new_n779), .B2(G159), .ZN(new_n814));
  INV_X1    g0614(.A(G137), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n814), .B1(new_n815), .B2(new_n746), .C1(new_n271), .C2(new_n770), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT34), .Z(new_n817));
  AOI21_X1  g0617(.A(new_n817), .B1(G132), .B2(new_n759), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n766), .A2(G50), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n755), .A2(G58), .ZN(new_n820));
  NAND4_X1  g0620(.A1(new_n818), .A2(new_n260), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n762), .A2(new_n303), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n813), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(new_n739), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n739), .A2(new_n736), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n392), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n805), .A2(new_n725), .A3(new_n824), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n804), .A2(new_n827), .ZN(G384));
  INV_X1    g0628(.A(KEYINPUT38), .ZN(new_n829));
  INV_X1    g0629(.A(new_n645), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n374), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n831), .B1(new_n366), .B2(new_n376), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n374), .B1(new_n371), .B2(new_n830), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT37), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n833), .A2(new_n834), .A3(new_n356), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n834), .B1(new_n833), .B2(new_n356), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n829), .B1(new_n832), .B2(new_n838), .ZN(new_n839));
  OR2_X1    g0639(.A1(new_n316), .A2(new_n317), .ZN(new_n840));
  AOI21_X1  g0640(.A(KEYINPUT16), .B1(new_n840), .B2(new_n309), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n318), .A2(new_n279), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n330), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AOI221_X4 g0643(.A(new_n367), .B1(new_n370), .B2(new_n369), .C1(new_n327), .C2(new_n330), .ZN(new_n844));
  AOI21_X1  g0644(.A(KEYINPUT18), .B1(new_n374), .B2(new_n371), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n358), .A2(new_n365), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n830), .B(new_n843), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n372), .A2(new_n645), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n843), .A2(new_n849), .B1(new_n368), .B2(new_n364), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n835), .B1(new_n850), .B2(new_n834), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n848), .A2(KEYINPUT38), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n839), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT96), .ZN(new_n854));
  OR3_X1    g0654(.A1(new_n853), .A2(new_n854), .A3(KEYINPUT39), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n839), .A2(new_n854), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n848), .A2(new_n851), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n829), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n852), .ZN(new_n859));
  OAI21_X1  g0659(.A(KEYINPUT39), .B1(new_n856), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n855), .A2(new_n860), .ZN(new_n861));
  AND3_X1   g0661(.A1(new_n423), .A2(new_n434), .A3(new_n648), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n794), .A2(new_n648), .A3(new_n796), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n801), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n434), .A2(new_n647), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n423), .A2(new_n434), .B1(new_n442), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n862), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  AND3_X1   g0669(.A1(new_n848), .A2(KEYINPUT38), .A3(new_n851), .ZN(new_n870));
  AOI21_X1  g0670(.A(KEYINPUT38), .B1(new_n848), .B2(new_n851), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n873), .B1(new_n846), .B2(new_n645), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n863), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n444), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n637), .B1(new_n694), .B2(new_n876), .ZN(new_n877));
  XNOR2_X1  g0677(.A(new_n875), .B(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT40), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n794), .A2(new_n796), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n880), .A2(new_n400), .A3(new_n798), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n793), .A2(new_n647), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AND3_X1   g0683(.A1(new_n717), .A2(KEYINPUT31), .A3(new_n647), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n868), .B(new_n883), .C1(new_n718), .C2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n879), .B1(new_n872), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n713), .A2(KEYINPUT31), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n717), .A2(new_n647), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n717), .A2(KEYINPUT31), .A3(new_n647), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n799), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n891), .A2(new_n853), .A3(KEYINPUT40), .A4(new_n868), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n886), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n889), .A2(new_n890), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n444), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n893), .B(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n652), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n878), .B(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n898), .B1(new_n247), .B2(new_n641), .ZN(new_n899));
  NOR3_X1   g0699(.A1(new_n226), .A2(new_n392), .A3(new_n304), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n303), .A2(G50), .ZN(new_n901));
  OAI211_X1 g0701(.A(G1), .B(new_n640), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n239), .B1(new_n542), .B2(KEYINPUT35), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n903), .B(new_n223), .C1(KEYINPUT35), .C2(new_n542), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n904), .B(KEYINPUT95), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n905), .B(KEYINPUT36), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n899), .A2(new_n902), .A3(new_n906), .ZN(G367));
  INV_X1    g0707(.A(new_n663), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n561), .B(new_n573), .C1(new_n548), .C2(new_n648), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n629), .A2(new_n647), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n603), .A2(new_n648), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n627), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT43), .ZN(new_n915));
  OR2_X1    g0715(.A1(new_n619), .A2(new_n913), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT97), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n917), .B(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(KEYINPUT42), .B1(new_n665), .B2(new_n909), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT42), .ZN(new_n921));
  INV_X1    g0721(.A(new_n909), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n659), .A2(new_n664), .A3(new_n921), .A4(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n629), .B1(new_n657), .B2(new_n922), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n920), .B(new_n923), .C1(new_n647), .C2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n914), .A2(new_n916), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(KEYINPUT43), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n919), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n928), .B(KEYINPUT98), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n925), .A2(new_n919), .A3(new_n927), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT100), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n925), .A2(new_n919), .A3(KEYINPUT100), .A4(new_n927), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n929), .A2(KEYINPUT99), .A3(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT99), .B1(new_n929), .B2(new_n934), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n912), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n937), .ZN(new_n939));
  INV_X1    g0739(.A(new_n912), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n939), .A2(new_n940), .A3(new_n935), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n673), .B(KEYINPUT41), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT44), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n668), .B2(new_n911), .ZN(new_n944));
  INV_X1    g0744(.A(new_n911), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n667), .A2(KEYINPUT44), .A3(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n944), .A2(KEYINPUT103), .A3(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT103), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n948), .B(new_n943), .C1(new_n668), .C2(new_n911), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT45), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n668), .A2(new_n951), .A3(new_n911), .ZN(new_n952));
  OAI21_X1  g0752(.A(KEYINPUT45), .B1(new_n667), .B2(new_n945), .ZN(new_n953));
  XNOR2_X1  g0753(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n952), .A2(new_n953), .ZN(new_n956));
  INV_X1    g0756(.A(new_n954), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n950), .A2(new_n663), .A3(new_n955), .A4(new_n958), .ZN(new_n959));
  NAND4_X1  g0759(.A1(new_n958), .A2(new_n947), .A3(new_n955), .A4(new_n949), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n908), .ZN(new_n961));
  AND2_X1   g0761(.A1(new_n663), .A2(KEYINPUT104), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n665), .B1(new_n662), .B2(new_n664), .ZN(new_n963));
  AND2_X1   g0763(.A1(new_n963), .A2(new_n653), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n663), .A2(KEYINPUT104), .ZN(new_n965));
  NOR3_X1   g0765(.A1(new_n962), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n959), .A2(new_n961), .A3(new_n720), .A4(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n942), .B1(new_n967), .B2(new_n720), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n938), .B(new_n941), .C1(new_n968), .C2(new_n724), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n740), .B1(new_n236), .B2(new_n730), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(new_n670), .B2(new_n396), .ZN(new_n971));
  AOI22_X1  g0771(.A1(G143), .A2(new_n785), .B1(new_n768), .B2(G150), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n972), .B1(new_n302), .B2(new_n765), .C1(new_n781), .C2(new_n770), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n463), .B1(new_n763), .B2(G77), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n974), .A2(KEYINPUT105), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n754), .A2(new_n303), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n976), .B1(G137), .B2(new_n759), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n974), .A2(KEYINPUT105), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n975), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  AOI211_X1 g0779(.A(new_n973), .B(new_n979), .C1(G50), .C2(new_n779), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n260), .B1(new_n755), .B2(G107), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n763), .A2(G97), .ZN(new_n982));
  INV_X1    g0782(.A(G294), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n981), .B(new_n982), .C1(new_n983), .C2(new_n770), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n766), .A2(G116), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT46), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n985), .A2(new_n986), .B1(G311), .B2(new_n785), .ZN(new_n987));
  AOI22_X1  g0787(.A1(G303), .A2(new_n768), .B1(new_n779), .B2(G283), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n987), .B(new_n988), .C1(new_n986), .C2(new_n985), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n984), .B(new_n989), .C1(G317), .C2(new_n759), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n980), .A2(new_n990), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n991), .B(KEYINPUT47), .Z(new_n992));
  AOI21_X1  g0792(.A(new_n971), .B1(new_n992), .B2(new_n739), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n993), .B(new_n725), .C1(new_n743), .C2(new_n926), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n969), .A2(new_n994), .ZN(G387));
  NOR2_X1   g0795(.A1(new_n662), .A2(new_n743), .ZN(new_n996));
  AOI211_X1 g0796(.A(G45), .B(new_n675), .C1(G68), .C2(G77), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT106), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n276), .A2(G50), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT50), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n730), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n1001), .B(KEYINPUT107), .Z(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n467), .B2(new_n232), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n1003), .B1(G107), .B2(new_n206), .C1(new_n676), .C2(new_n734), .ZN(new_n1004));
  AND2_X1   g0804(.A1(new_n1004), .A2(new_n740), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(G68), .A2(new_n779), .B1(new_n759), .B2(G150), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n601), .B2(new_n754), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n767), .A2(new_n280), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n770), .A2(new_n276), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n765), .A2(new_n392), .ZN(new_n1010));
  NOR4_X1   g0810(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n785), .A2(G159), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1011), .A2(new_n260), .A3(new_n982), .A4(new_n1012), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(G322), .A2(new_n785), .B1(new_n771), .B2(G311), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(KEYINPUT108), .Z(new_n1015));
  INV_X1    g0815(.A(G317), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1015), .B1(new_n806), .B2(new_n750), .C1(new_n1016), .C2(new_n767), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT48), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n755), .A2(G283), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1018), .B(new_n1019), .C1(new_n983), .C2(new_n765), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT49), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n260), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n1022), .B1(new_n1021), .B2(new_n1020), .C1(new_n239), .C2(new_n762), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n758), .A2(new_n747), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1013), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n996), .B(new_n1005), .C1(new_n739), .C2(new_n1025), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n1026), .A2(new_n725), .B1(new_n724), .B2(new_n966), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n966), .A2(new_n720), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n966), .A2(new_n720), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1028), .A2(new_n722), .A3(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1027), .A2(new_n1030), .ZN(G393));
  NAND3_X1  g0831(.A1(new_n959), .A2(new_n961), .A3(KEYINPUT109), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT109), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n960), .A2(new_n1033), .A3(new_n908), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1032), .A2(new_n1029), .A3(new_n1034), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1035), .A2(new_n722), .A3(new_n967), .ZN(new_n1036));
  INV_X1    g0836(.A(G143), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n750), .A2(new_n276), .B1(new_n758), .B2(new_n1037), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n746), .A2(new_n271), .B1(new_n767), .B2(new_n781), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT51), .Z(new_n1040));
  AOI211_X1 g0840(.A(new_n1038), .B(new_n1040), .C1(G77), .C2(new_n755), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1041), .B1(new_n280), .B2(new_n770), .C1(new_n303), .C2(new_n765), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n463), .B(new_n1042), .C1(G87), .C2(new_n763), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n746), .A2(new_n1016), .B1(new_n767), .B2(new_n751), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT52), .Z(new_n1045));
  AOI22_X1  g0845(.A1(G303), .A2(new_n771), .B1(new_n779), .B2(G294), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n766), .A2(G283), .B1(new_n755), .B2(G116), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n784), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n260), .B1(new_n759), .B2(G322), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .A4(new_n1049), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1045), .A2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n739), .B1(new_n1043), .B2(new_n1051), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n740), .B1(new_n545), .B2(new_n206), .C1(new_n242), .C2(new_n730), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1052), .A2(new_n725), .A3(new_n1053), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n1054), .A2(KEYINPUT111), .B1(new_n738), .B2(new_n945), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(KEYINPUT111), .B2(new_n1054), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1036), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT110), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1032), .A2(KEYINPUT110), .A3(new_n1034), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1061), .A2(new_n724), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1058), .A2(new_n1063), .ZN(G390));
  INV_X1    g0864(.A(new_n862), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n869), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n855), .A2(new_n860), .A3(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n862), .B1(new_n839), .B2(new_n852), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n692), .A2(new_n648), .A3(new_n797), .ZN(new_n1069));
  AND2_X1   g0869(.A1(new_n1069), .A2(new_n864), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n868), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1068), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n652), .B(new_n883), .C1(new_n712), .C2(new_n718), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n868), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT112), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n891), .A2(new_n1077), .A3(G330), .ZN(new_n1078));
  AND4_X1   g0878(.A1(new_n1067), .A2(new_n1072), .A3(new_n1076), .A4(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(G330), .ZN(new_n1080));
  NOR3_X1   g0880(.A1(new_n885), .A2(new_n1077), .A3(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(new_n1067), .B2(new_n1072), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1079), .A2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n444), .A2(G330), .A3(new_n894), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1084), .B(new_n637), .C1(new_n694), .C2(new_n876), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1074), .A2(new_n868), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n885), .A2(new_n1080), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n865), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n891), .A2(G330), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n1071), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1090), .A2(new_n1075), .A3(new_n1070), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1085), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n673), .B1(new_n1083), .B2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1092), .B1(new_n1079), .B2(new_n1082), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1067), .A2(new_n1072), .A3(new_n1076), .A4(new_n1078), .ZN(new_n1097));
  AND2_X1   g0897(.A1(new_n1067), .A2(new_n1072), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1097), .B1(new_n1098), .B2(new_n1081), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n724), .ZN(new_n1100));
  INV_X1    g0900(.A(G128), .ZN(new_n1101));
  INV_X1    g0901(.A(G132), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n746), .A2(new_n1101), .B1(new_n767), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT53), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n766), .B2(G150), .ZN(new_n1105));
  XOR2_X1   g0905(.A(KEYINPUT54), .B(G143), .Z(new_n1106));
  AOI211_X1 g0906(.A(new_n1103), .B(new_n1105), .C1(new_n779), .C2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n770), .A2(new_n815), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n260), .B1(new_n762), .B2(new_n280), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n1108), .B(new_n1109), .C1(G125), .C2(new_n759), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n755), .A2(G159), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n766), .A2(new_n1104), .A3(G150), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1107), .A2(new_n1110), .A3(new_n1111), .A4(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n463), .B1(new_n765), .B2(new_n210), .ZN(new_n1114));
  XOR2_X1   g0914(.A(new_n1114), .B(KEYINPUT113), .Z(new_n1115));
  OAI22_X1  g0915(.A1(new_n767), .A2(new_n239), .B1(new_n758), .B2(new_n983), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n822), .B(new_n1116), .C1(G107), .C2(new_n771), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n779), .A2(G97), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n785), .A2(G283), .B1(new_n755), .B2(G77), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1115), .A2(new_n1117), .A3(new_n1118), .A4(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n789), .B1(new_n1113), .B2(new_n1120), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n728), .B(new_n1121), .C1(new_n276), .C2(new_n825), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1122), .B1(new_n861), .B2(new_n737), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1096), .A2(new_n1100), .A3(new_n1123), .ZN(G378));
  INV_X1    g0924(.A(KEYINPUT57), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n886), .A2(G330), .A3(new_n892), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT117), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n886), .A2(new_n892), .A3(KEYINPUT117), .A4(G330), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT115), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n301), .B(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n287), .A2(new_n830), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1133), .B(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1130), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n863), .A2(new_n874), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1135), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1136), .A2(new_n1137), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1135), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n875), .B1(new_n1142), .B2(new_n1138), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1088), .A2(new_n1091), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1085), .B1(new_n1099), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1125), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1085), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1095), .A2(new_n1148), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1149), .A2(KEYINPUT57), .A3(new_n1143), .A4(new_n1140), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1147), .A2(new_n722), .A3(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1140), .A2(new_n724), .A3(new_n1143), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1135), .A2(new_n736), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n754), .A2(new_n271), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n770), .A2(new_n1102), .B1(new_n750), .B2(new_n815), .ZN(new_n1155));
  XOR2_X1   g0955(.A(new_n1155), .B(KEYINPUT114), .Z(new_n1156));
  AOI211_X1 g0956(.A(new_n1154), .B(new_n1156), .C1(G125), .C2(new_n785), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n1101), .B2(new_n767), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(new_n766), .B2(new_n1106), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n1159), .B(KEYINPUT59), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n257), .B1(new_n762), .B2(new_n781), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(G124), .B2(new_n759), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1160), .A2(new_n470), .A3(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n280), .B1(new_n338), .B2(G41), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n601), .A2(new_n750), .B1(new_n302), .B2(new_n762), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n463), .B1(new_n746), .B2(new_n239), .ZN(new_n1166));
  NOR4_X1   g0966(.A1(new_n1165), .A2(new_n1166), .A3(G41), .A4(new_n976), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1010), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(G97), .A2(new_n771), .B1(new_n759), .B2(G283), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n768), .A2(G107), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1167), .A2(new_n1168), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT58), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1163), .A2(new_n1164), .A3(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n739), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n825), .A2(new_n280), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1153), .A2(new_n725), .A3(new_n1174), .A4(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT116), .ZN(new_n1177));
  AND2_X1   g0977(.A1(new_n1152), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1151), .A2(new_n1178), .ZN(G375));
  INV_X1    g0979(.A(new_n942), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1088), .A2(new_n1091), .A3(new_n1085), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1093), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n260), .B1(new_n762), .B2(new_n302), .ZN(new_n1183));
  XOR2_X1   g0983(.A(new_n1183), .B(KEYINPUT119), .Z(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(new_n771), .B2(new_n1106), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n765), .A2(new_n781), .B1(new_n758), .B2(new_n1101), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1186), .B(KEYINPUT120), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n750), .A2(new_n271), .B1(new_n754), .B2(new_n280), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n785), .A2(G132), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n768), .A2(G137), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1185), .A2(new_n1189), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n770), .A2(new_n239), .B1(new_n762), .B2(new_n392), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n260), .B(new_n1193), .C1(G303), .C2(new_n759), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n766), .A2(G97), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n768), .A2(G283), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n601), .A2(new_n754), .B1(new_n983), .B2(new_n746), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(G107), .B2(new_n779), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .A4(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n789), .B1(new_n1192), .B2(new_n1199), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n728), .B(new_n1200), .C1(new_n303), .C2(new_n825), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1071), .A2(new_n736), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n1202), .B(KEYINPUT118), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n1145), .A2(new_n724), .B1(new_n1201), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1182), .A2(new_n1204), .ZN(G381));
  NOR2_X1   g1005(.A1(G390), .A2(G381), .ZN(new_n1206));
  INV_X1    g1006(.A(G387), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1027), .A2(new_n1030), .A3(new_n791), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1208), .A2(G384), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(KEYINPUT121), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1206), .A2(new_n1207), .A3(new_n1210), .ZN(new_n1211));
  XOR2_X1   g1011(.A(new_n1211), .B(KEYINPUT122), .Z(new_n1212));
  NAND2_X1  g1012(.A1(new_n1100), .A2(new_n1123), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(new_n1095), .B2(new_n1094), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(G375), .A2(KEYINPUT123), .ZN(new_n1215));
  OR2_X1    g1015(.A1(G375), .A2(KEYINPUT123), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1212), .A2(new_n1214), .A3(new_n1215), .A4(new_n1216), .ZN(G407));
  NAND4_X1  g1017(.A1(new_n1216), .A2(new_n646), .A3(new_n1214), .A4(new_n1215), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(G407), .A2(G213), .A3(new_n1218), .ZN(G409));
  NAND3_X1  g1019(.A1(new_n1151), .A2(G378), .A3(new_n1178), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1149), .A2(new_n1180), .A3(new_n1143), .A4(new_n1140), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1221), .A2(new_n1152), .A3(new_n1176), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(new_n1214), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1220), .A2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT60), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1093), .B(new_n722), .C1(new_n1225), .C2(new_n1181), .ZN(new_n1226));
  AND2_X1   g1026(.A1(new_n1181), .A2(new_n1225), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1204), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1228), .A2(new_n804), .A3(new_n827), .ZN(new_n1229));
  OAI211_X1 g1029(.A(G384), .B(new_n1204), .C1(new_n1226), .C2(new_n1227), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(G213), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1233), .A2(G343), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1224), .A2(new_n1232), .A3(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT124), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT62), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1234), .B1(new_n1220), .B2(new_n1223), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1240), .A2(KEYINPUT124), .A3(new_n1232), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1238), .A2(new_n1239), .A3(new_n1241), .ZN(new_n1242));
  AND2_X1   g1042(.A1(new_n1234), .A2(G2897), .ZN(new_n1243));
  AND3_X1   g1043(.A1(new_n1229), .A2(new_n1230), .A3(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1243), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1239), .B1(new_n1240), .B2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(KEYINPUT61), .B1(new_n1247), .B2(new_n1236), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1242), .A2(new_n1248), .ZN(new_n1249));
  AND3_X1   g1049(.A1(new_n1061), .A2(new_n724), .A3(new_n1062), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n969), .B(new_n994), .C1(new_n1250), .C2(new_n1057), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT126), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(G393), .A2(G396), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(new_n1208), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(G387), .A2(new_n1058), .A3(new_n1063), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n1253), .A2(new_n1255), .B1(new_n1251), .B2(new_n1256), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1256), .A2(new_n1251), .A3(KEYINPUT126), .A4(new_n1255), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT127), .ZN(new_n1260));
  NOR3_X1   g1060(.A1(new_n1257), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1256), .A2(new_n1251), .ZN(new_n1262));
  AOI21_X1  g1062(.A(KEYINPUT126), .B1(new_n1207), .B2(G390), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1255), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1262), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(KEYINPUT127), .B1(new_n1265), .B2(new_n1258), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1261), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1249), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT63), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1241), .ZN(new_n1270));
  AOI21_X1  g1070(.A(KEYINPUT124), .B1(new_n1240), .B2(new_n1232), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1269), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT125), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1240), .B1(new_n1273), .B2(new_n1246), .ZN(new_n1274));
  OAI21_X1  g1074(.A(KEYINPUT125), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n1274), .A2(new_n1275), .B1(new_n1258), .B2(new_n1265), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1236), .A2(new_n1269), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1277), .A2(KEYINPUT61), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1272), .A2(new_n1276), .A3(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1268), .A2(new_n1279), .ZN(G405));
  INV_X1    g1080(.A(new_n1220), .ZN(new_n1281));
  AOI21_X1  g1081(.A(G378), .B1(new_n1151), .B2(new_n1178), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  XNOR2_X1  g1083(.A(new_n1283), .B(new_n1231), .ZN(new_n1284));
  XNOR2_X1  g1084(.A(new_n1267), .B(new_n1284), .ZN(G402));
endmodule


