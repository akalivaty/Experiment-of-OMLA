//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 1 0 1 1 0 1 0 0 1 1 1 0 1 1 0 1 1 1 0 0 0 0 1 1 1 0 0 1 1 0 0 0 1 1 0 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:59 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000;
  INV_X1    g000(.A(KEYINPUT71), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT67), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  OAI211_X1 g007(.A(KEYINPUT64), .B(KEYINPUT1), .C1(new_n191), .C2(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G128), .ZN(new_n195));
  AOI21_X1  g009(.A(KEYINPUT64), .B1(new_n190), .B2(KEYINPUT1), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n193), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  XNOR2_X1  g011(.A(G143), .B(G146), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT1), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n198), .A2(new_n199), .A3(G128), .ZN(new_n200));
  AND3_X1   g014(.A1(new_n197), .A2(KEYINPUT66), .A3(new_n200), .ZN(new_n201));
  AOI21_X1  g015(.A(KEYINPUT66), .B1(new_n197), .B2(new_n200), .ZN(new_n202));
  INV_X1    g016(.A(G134), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G137), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n203), .A2(G137), .ZN(new_n206));
  OAI21_X1  g020(.A(G131), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT11), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n208), .B1(new_n203), .B2(G137), .ZN(new_n209));
  INV_X1    g023(.A(G137), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(KEYINPUT11), .A3(G134), .ZN(new_n211));
  INV_X1    g025(.A(G131), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n209), .A2(new_n211), .A3(new_n212), .A4(new_n204), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n207), .A2(new_n213), .ZN(new_n214));
  NOR3_X1   g028(.A1(new_n201), .A2(new_n202), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(KEYINPUT0), .A2(G128), .ZN(new_n216));
  OR2_X1    g030(.A1(KEYINPUT0), .A2(G128), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n193), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n198), .A2(KEYINPUT0), .A3(G128), .ZN(new_n219));
  AND2_X1   g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n209), .A2(new_n204), .A3(new_n211), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G131), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(new_n213), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n188), .B1(new_n215), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G119), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G116), .ZN(new_n228));
  INV_X1    g042(.A(G116), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G119), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT65), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT2), .B(G113), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT65), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n228), .A2(new_n230), .A3(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n232), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  OR2_X1    g050(.A1(new_n231), .A2(new_n233), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n197), .A2(new_n200), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT66), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n214), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n197), .A2(KEYINPUT66), .A3(new_n200), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n242), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n245), .A2(KEYINPUT67), .A3(new_n224), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n226), .A2(new_n239), .A3(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT28), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NOR2_X1   g063(.A1(G237), .A2(G953), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G210), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n251), .B(KEYINPUT27), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT26), .B(G101), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n252), .B(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n245), .A2(new_n239), .A3(new_n224), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n214), .B1(new_n197), .B2(new_n200), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n238), .B1(new_n225), .B2(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n248), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n249), .A2(new_n254), .A3(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n245), .A2(KEYINPUT30), .A3(new_n224), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT30), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n262), .B1(new_n225), .B2(new_n256), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n261), .A2(new_n263), .A3(new_n238), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(new_n255), .ZN(new_n265));
  INV_X1    g079(.A(new_n254), .ZN(new_n266));
  AOI21_X1  g080(.A(KEYINPUT29), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n260), .A2(new_n267), .ZN(new_n268));
  XOR2_X1   g082(.A(KEYINPUT69), .B(G902), .Z(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n254), .A2(KEYINPUT29), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n271), .B1(new_n247), .B2(new_n248), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n238), .B1(new_n215), .B2(new_n225), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n273), .A2(KEYINPUT68), .A3(new_n255), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n245), .A2(new_n224), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT68), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n275), .A2(new_n276), .A3(new_n238), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n274), .A2(KEYINPUT28), .A3(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n270), .B1(new_n272), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n268), .B1(new_n279), .B2(KEYINPUT70), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT70), .ZN(new_n281));
  AOI211_X1 g095(.A(new_n281), .B(new_n270), .C1(new_n272), .C2(new_n278), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n187), .B(G472), .C1(new_n280), .C2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n249), .A2(new_n259), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n264), .A2(new_n255), .A3(new_n254), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT31), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n264), .A2(KEYINPUT31), .A3(new_n255), .A4(new_n254), .ZN(new_n288));
  AOI22_X1  g102(.A1(new_n266), .A2(new_n284), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NOR2_X1   g103(.A1(G472), .A2(G902), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(KEYINPUT32), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n287), .A2(new_n288), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n238), .B1(new_n275), .B2(new_n188), .ZN(new_n294));
  AOI21_X1  g108(.A(KEYINPUT28), .B1(new_n294), .B2(new_n246), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n266), .B1(new_n295), .B2(new_n258), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT32), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n297), .A2(new_n298), .A3(new_n290), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n292), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n283), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n272), .A2(new_n278), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n269), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n281), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n279), .A2(KEYINPUT70), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n304), .A2(new_n305), .A3(new_n268), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n187), .B1(new_n306), .B2(G472), .ZN(new_n307));
  OAI21_X1  g121(.A(KEYINPUT72), .B1(new_n301), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G475), .ZN(new_n309));
  INV_X1    g123(.A(G140), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G125), .ZN(new_n311));
  INV_X1    g125(.A(G125), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G140), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n311), .A2(new_n313), .A3(KEYINPUT16), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n312), .A2(G140), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT16), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AND3_X1   g131(.A1(new_n314), .A2(G146), .A3(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(G146), .B1(new_n314), .B2(new_n317), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G237), .ZN(new_n321));
  INV_X1    g135(.A(G953), .ZN(new_n322));
  AND4_X1   g136(.A1(G143), .A2(new_n321), .A3(new_n322), .A4(G214), .ZN(new_n323));
  AOI21_X1  g137(.A(G143), .B1(new_n250), .B2(G214), .ZN(new_n324));
  OAI21_X1  g138(.A(G131), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT88), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n321), .A2(new_n322), .A3(G214), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n191), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n250), .A2(G143), .A3(G214), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(KEYINPUT88), .A3(G131), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT17), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n329), .A2(new_n212), .A3(new_n330), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n327), .A2(new_n332), .A3(new_n333), .A4(new_n334), .ZN(new_n335));
  AND2_X1   g149(.A1(new_n327), .A2(new_n332), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n320), .B(new_n335), .C1(new_n336), .C2(new_n333), .ZN(new_n337));
  XNOR2_X1  g151(.A(G125), .B(G140), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n189), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n310), .A2(G125), .ZN(new_n340));
  OAI21_X1  g154(.A(G146), .B1(new_n315), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(KEYINPUT87), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT87), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n339), .A2(new_n341), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT18), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n331), .B1(new_n347), .B2(new_n212), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n329), .A2(KEYINPUT18), .A3(G131), .A4(new_n330), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n337), .A2(new_n351), .ZN(new_n352));
  XOR2_X1   g166(.A(G113), .B(G122), .Z(new_n353));
  XOR2_X1   g167(.A(KEYINPUT90), .B(G104), .Z(new_n354));
  XOR2_X1   g168(.A(new_n353), .B(new_n354), .Z(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n352), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n337), .A2(new_n355), .A3(new_n351), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(G902), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n309), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NOR2_X1   g175(.A1(G475), .A2(G902), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n327), .A2(new_n332), .A3(new_n334), .ZN(new_n363));
  AND3_X1   g177(.A1(new_n311), .A2(new_n313), .A3(KEYINPUT19), .ZN(new_n364));
  AOI21_X1  g178(.A(KEYINPUT19), .B1(new_n311), .B2(new_n313), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n189), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n318), .B1(new_n366), .B2(KEYINPUT89), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT19), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n368), .B1(new_n315), .B2(new_n340), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n311), .A2(new_n313), .A3(KEYINPUT19), .ZN(new_n370));
  AOI21_X1  g184(.A(G146), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT89), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n363), .A2(new_n367), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n351), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT91), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(new_n376), .A3(new_n356), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n358), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n376), .B1(new_n375), .B2(new_n356), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n362), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT20), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT20), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n382), .B(new_n362), .C1(new_n378), .C2(new_n379), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n361), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT15), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G478), .ZN(new_n386));
  XNOR2_X1  g200(.A(KEYINPUT9), .B(G234), .ZN(new_n387));
  INV_X1    g201(.A(G217), .ZN(new_n388));
  NOR3_X1   g202(.A1(new_n387), .A2(new_n388), .A3(G953), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT94), .ZN(new_n391));
  INV_X1    g205(.A(G128), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G143), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n191), .A2(G128), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n393), .A2(new_n394), .A3(KEYINPUT93), .A4(new_n203), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n229), .A2(G122), .ZN(new_n396));
  INV_X1    g210(.A(G122), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G116), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G107), .ZN(new_n400));
  XNOR2_X1  g214(.A(G116), .B(G122), .ZN(new_n401));
  INV_X1    g215(.A(G107), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT93), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n393), .A2(new_n394), .A3(new_n203), .ZN(new_n405));
  AOI22_X1  g219(.A1(new_n400), .A2(new_n403), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(KEYINPUT13), .B1(new_n191), .B2(G128), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT92), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n407), .A2(new_n408), .A3(new_n394), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n408), .B1(new_n407), .B2(new_n394), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n392), .A2(G143), .ZN(new_n412));
  AND2_X1   g226(.A1(new_n412), .A2(KEYINPUT13), .ZN(new_n413));
  NOR3_X1   g227(.A1(new_n410), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n395), .B(new_n406), .C1(new_n414), .C2(new_n203), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n393), .A2(new_n394), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(G134), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n405), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n229), .A2(KEYINPUT14), .A3(G122), .ZN(new_n419));
  OAI211_X1 g233(.A(G107), .B(new_n419), .C1(new_n399), .C2(KEYINPUT14), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n418), .A2(new_n420), .A3(new_n403), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n391), .B1(new_n415), .B2(new_n421), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n411), .A2(new_n413), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n203), .B1(new_n423), .B2(new_n409), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n400), .A2(new_n403), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n405), .A2(new_n404), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(new_n395), .A3(new_n426), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n391), .B(new_n421), .C1(new_n424), .C2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n390), .B1(new_n422), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n421), .B1(new_n424), .B2(new_n427), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT94), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n432), .A2(new_n389), .A3(new_n428), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n270), .B1(new_n430), .B2(new_n433), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n434), .A2(KEYINPUT95), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT95), .ZN(new_n436));
  AOI211_X1 g250(.A(new_n436), .B(new_n270), .C1(new_n430), .C2(new_n433), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n386), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  OR2_X1    g252(.A1(new_n437), .A2(new_n386), .ZN(new_n439));
  AND2_X1   g253(.A1(new_n322), .A2(G952), .ZN(new_n440));
  NAND2_X1  g254(.A1(G234), .A2(G237), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  XOR2_X1   g256(.A(new_n442), .B(KEYINPUT96), .Z(new_n443));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(G898), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n270), .A2(G953), .A3(new_n441), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n443), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n384), .A2(new_n438), .A3(new_n439), .A4(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(G210), .B1(G237), .B2(G902), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(G104), .ZN(new_n451));
  OAI21_X1  g265(.A(KEYINPUT3), .B1(new_n451), .B2(G107), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT3), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n453), .A2(new_n402), .A3(G104), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n451), .A2(G107), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n452), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT4), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n456), .A2(new_n457), .A3(G101), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(G101), .ZN(new_n459));
  INV_X1    g273(.A(G101), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n452), .A2(new_n454), .A3(new_n460), .A4(new_n455), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n459), .A2(KEYINPUT4), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n238), .A2(new_n458), .A3(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n402), .A2(G104), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n451), .A2(G107), .ZN(new_n465));
  OAI21_X1  g279(.A(G101), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n461), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT5), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n468), .B1(new_n232), .B2(new_n235), .ZN(new_n469));
  OAI21_X1  g283(.A(G113), .B1(new_n228), .B2(KEYINPUT5), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n237), .B(new_n467), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n463), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(G110), .B(G122), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n463), .A2(new_n471), .A3(new_n473), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n475), .A2(KEYINPUT6), .A3(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT6), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n472), .A2(new_n478), .A3(new_n474), .ZN(new_n479));
  OAI21_X1  g293(.A(KEYINPUT84), .B1(new_n220), .B2(new_n312), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n197), .A2(new_n312), .A3(new_n200), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n218), .A2(new_n219), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT84), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(new_n483), .A3(G125), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n480), .A2(new_n481), .A3(new_n484), .ZN(new_n485));
  XOR2_X1   g299(.A(KEYINPUT85), .B(G224), .Z(new_n486));
  NOR2_X1   g300(.A1(new_n486), .A2(G953), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n487), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n480), .A2(new_n489), .A3(new_n481), .A4(new_n484), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n477), .A2(new_n479), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT7), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n485), .B1(new_n493), .B2(new_n487), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n487), .A2(new_n493), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n480), .A2(new_n481), .A3(new_n495), .A4(new_n484), .ZN(new_n496));
  XOR2_X1   g310(.A(new_n473), .B(KEYINPUT8), .Z(new_n497));
  NOR2_X1   g311(.A1(new_n231), .A2(new_n468), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n237), .B1(new_n498), .B2(new_n470), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n497), .B1(new_n499), .B2(new_n467), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n237), .B1(new_n469), .B2(new_n470), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n500), .B1(new_n501), .B2(new_n467), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n494), .A2(new_n476), .A3(new_n496), .A4(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n360), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n450), .B1(new_n492), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n477), .A2(new_n491), .A3(new_n479), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n506), .A2(new_n360), .A3(new_n449), .A4(new_n503), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(G214), .B1(G237), .B2(G902), .ZN(new_n509));
  AOI21_X1  g323(.A(KEYINPUT86), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT86), .ZN(new_n511));
  INV_X1    g325(.A(new_n509), .ZN(new_n512));
  AOI211_X1 g326(.A(new_n511), .B(new_n512), .C1(new_n505), .C2(new_n507), .ZN(new_n513));
  NOR3_X1   g327(.A1(new_n448), .A2(new_n510), .A3(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(G221), .B1(new_n387), .B2(G902), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n461), .A2(new_n466), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT10), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n242), .A2(new_n244), .A3(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n223), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n392), .B1(new_n190), .B2(KEYINPUT1), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n200), .B1(new_n198), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n467), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n518), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n462), .A2(new_n220), .A3(new_n458), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n520), .A2(new_n521), .A3(new_n525), .A4(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT80), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AND2_X1   g343(.A1(new_n525), .A2(new_n526), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n530), .A2(KEYINPUT80), .A3(new_n521), .A4(new_n520), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n530), .A2(new_n520), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n223), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g349(.A(G110), .B(G140), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n322), .A2(G227), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n536), .B(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n535), .A2(KEYINPUT83), .A3(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT83), .ZN(new_n540));
  AOI22_X1  g354(.A1(new_n529), .A2(new_n531), .B1(new_n223), .B2(new_n533), .ZN(new_n541));
  INV_X1    g355(.A(new_n538), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n197), .A2(new_n517), .A3(new_n200), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n521), .B1(new_n524), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT81), .ZN(new_n546));
  AOI21_X1  g360(.A(KEYINPUT12), .B1(new_n223), .B2(new_n546), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n545), .B(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n538), .B1(new_n529), .B2(new_n531), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT82), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AOI211_X1 g366(.A(KEYINPUT82), .B(new_n538), .C1(new_n529), .C2(new_n531), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n539), .B(new_n543), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(G469), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n554), .A2(new_n555), .A3(new_n269), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n555), .A2(new_n360), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n532), .A2(new_n549), .ZN(new_n558));
  AOI22_X1  g372(.A1(new_n558), .A2(new_n538), .B1(new_n550), .B2(new_n534), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n557), .B1(new_n559), .B2(G469), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n516), .B1(new_n556), .B2(new_n560), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n514), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT78), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT25), .ZN(new_n564));
  AOI21_X1  g378(.A(KEYINPUT79), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n565), .B1(KEYINPUT79), .B2(new_n564), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n392), .A2(G119), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n227), .A2(G128), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n569), .B(KEYINPUT74), .ZN(new_n570));
  XOR2_X1   g384(.A(KEYINPUT24), .B(G110), .Z(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(G110), .ZN(new_n573));
  OAI21_X1  g387(.A(KEYINPUT75), .B1(new_n227), .B2(G128), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(KEYINPUT23), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT23), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n567), .A2(KEYINPUT75), .A3(new_n576), .ZN(new_n577));
  AND3_X1   g391(.A1(new_n575), .A2(new_n577), .A3(new_n568), .ZN(new_n578));
  OAI221_X1 g392(.A(new_n572), .B1(new_n573), .B2(new_n578), .C1(new_n319), .C2(new_n318), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n314), .A2(new_n317), .A3(G146), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n570), .A2(new_n571), .ZN(new_n581));
  XNOR2_X1  g395(.A(KEYINPUT76), .B(G110), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n580), .B(new_n339), .C1(new_n581), .C2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n322), .A2(G221), .A3(G234), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(KEYINPUT77), .ZN(new_n586));
  XNOR2_X1  g400(.A(KEYINPUT22), .B(G137), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n586), .B(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n579), .A2(new_n584), .A3(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n588), .B1(new_n579), .B2(new_n584), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n269), .B(new_n566), .C1(new_n590), .C2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n388), .B1(new_n269), .B2(G234), .ZN(new_n593));
  XOR2_X1   g407(.A(new_n593), .B(KEYINPUT73), .Z(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n591), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n270), .B1(new_n596), .B2(new_n589), .ZN(new_n597));
  INV_X1    g411(.A(new_n565), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n592), .B(new_n595), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n360), .B(new_n594), .C1(new_n590), .C2(new_n591), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(G472), .B1(new_n280), .B2(new_n282), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(KEYINPUT71), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT72), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n604), .A2(new_n605), .A3(new_n300), .A4(new_n283), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n308), .A2(new_n562), .A3(new_n602), .A4(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(KEYINPUT97), .B(G101), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(G3));
  OAI21_X1  g423(.A(G472), .B1(new_n289), .B2(new_n270), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n297), .A2(new_n290), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n612), .A2(new_n601), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT98), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT33), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n432), .A2(new_n389), .A3(new_n428), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n389), .B1(new_n432), .B2(new_n428), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n430), .A2(KEYINPUT33), .A3(new_n433), .ZN(new_n619));
  INV_X1    g433(.A(G478), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n270), .A2(new_n620), .ZN(new_n621));
  AND4_X1   g435(.A1(new_n614), .A2(new_n618), .A3(new_n619), .A4(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n618), .A2(new_n619), .A3(new_n621), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n430), .A2(new_n433), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n269), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n614), .B1(new_n625), .B2(new_n620), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n622), .B1(new_n623), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n359), .A2(new_n360), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(G475), .ZN(new_n629));
  INV_X1    g443(.A(new_n383), .ZN(new_n630));
  AOI22_X1  g444(.A1(new_n343), .A2(new_n345), .B1(new_n348), .B2(new_n349), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n580), .B1(new_n371), .B2(new_n372), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n366), .A2(KEYINPUT89), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n631), .B1(new_n634), .B2(new_n363), .ZN(new_n635));
  OAI21_X1  g449(.A(KEYINPUT91), .B1(new_n635), .B2(new_n355), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n636), .A2(new_n358), .A3(new_n377), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n382), .B1(new_n637), .B2(new_n362), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n629), .B1(new_n630), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n627), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n447), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n508), .A2(new_n509), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n613), .A2(new_n561), .A3(new_n642), .A4(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT34), .B(G104), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G6));
  NAND2_X1  g461(.A1(new_n438), .A2(new_n439), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n447), .B(KEYINPUT99), .Z(new_n649));
  NAND3_X1  g463(.A1(new_n648), .A2(new_n384), .A3(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT100), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n652), .A2(new_n561), .A3(new_n644), .A4(new_n613), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT102), .B(G107), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(KEYINPUT101), .B(KEYINPUT35), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G9));
  INV_X1    g471(.A(KEYINPUT104), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n579), .A2(new_n584), .ZN(new_n659));
  OR2_X1    g473(.A1(new_n588), .A2(KEYINPUT36), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n594), .A2(new_n360), .ZN(new_n662));
  OR3_X1    g476(.A1(new_n661), .A2(KEYINPUT103), .A3(new_n662), .ZN(new_n663));
  OAI21_X1  g477(.A(KEYINPUT103), .B1(new_n661), .B2(new_n662), .ZN(new_n664));
  AND3_X1   g478(.A1(new_n663), .A2(new_n599), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n658), .B1(new_n612), .B2(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n663), .A2(new_n599), .A3(new_n664), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n610), .A2(new_n611), .A3(KEYINPUT104), .A4(new_n667), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n666), .A2(new_n561), .A3(new_n514), .A4(new_n668), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT37), .B(G110), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G12));
  NAND2_X1  g485(.A1(new_n556), .A2(new_n560), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n443), .B1(G900), .B2(new_n446), .ZN(new_n673));
  AND3_X1   g487(.A1(new_n648), .A2(new_n384), .A3(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n665), .A2(new_n643), .ZN(new_n675));
  AND4_X1   g489(.A1(new_n515), .A2(new_n672), .A3(new_n674), .A4(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n308), .A2(new_n676), .A3(new_n606), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G128), .ZN(G30));
  XNOR2_X1  g492(.A(new_n673), .B(KEYINPUT39), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n561), .A2(new_n679), .ZN(new_n680));
  OR2_X1    g494(.A1(new_n680), .A2(KEYINPUT40), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n274), .A2(new_n277), .A3(new_n266), .ZN(new_n682));
  AND2_X1   g496(.A1(new_n682), .A2(KEYINPUT105), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n285), .B1(new_n682), .B2(KEYINPUT105), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n360), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(G472), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n300), .A2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n508), .B(KEYINPUT38), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n384), .B1(new_n438), .B2(new_n439), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n691), .A2(new_n509), .A3(new_n665), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n688), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n680), .A2(KEYINPUT40), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n681), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT106), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(new_n191), .ZN(G45));
  NAND2_X1  g511(.A1(new_n626), .A2(new_n623), .ZN(new_n698));
  AND2_X1   g512(.A1(new_n618), .A2(new_n619), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n699), .A2(new_n614), .A3(new_n621), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n639), .A2(new_n698), .A3(new_n700), .A4(new_n673), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n561), .A2(new_n702), .A3(new_n675), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n308), .A2(new_n703), .A3(new_n606), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G146), .ZN(G48));
  NAND3_X1  g519(.A1(new_n308), .A2(new_n602), .A3(new_n606), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n554), .A2(new_n269), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(G469), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n708), .A2(KEYINPUT107), .A3(new_n556), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT107), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n707), .A2(new_n710), .A3(G469), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n712), .A2(new_n515), .A3(new_n644), .A4(new_n642), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n706), .A2(new_n713), .ZN(new_n714));
  XOR2_X1   g528(.A(KEYINPUT41), .B(G113), .Z(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G15));
  NAND4_X1  g530(.A1(new_n712), .A2(new_n652), .A3(new_n515), .A4(new_n644), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n706), .A2(new_n717), .ZN(new_n718));
  XOR2_X1   g532(.A(KEYINPUT108), .B(G116), .Z(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(G18));
  AOI21_X1  g534(.A(new_n516), .B1(new_n709), .B2(new_n711), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n448), .A2(new_n643), .A3(new_n665), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n721), .A2(new_n308), .A3(new_n606), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(KEYINPUT109), .B(G119), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(G21));
  NAND2_X1  g539(.A1(new_n278), .A2(new_n249), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n254), .B1(new_n726), .B2(KEYINPUT110), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT110), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n278), .A2(new_n728), .A3(new_n249), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n293), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n290), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT111), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n732), .A2(new_n733), .A3(new_n602), .A4(new_n610), .ZN(new_n734));
  AOI22_X1  g548(.A1(new_n727), .A2(new_n729), .B1(new_n287), .B2(new_n288), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n602), .B(new_n610), .C1(new_n735), .C2(new_n291), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(KEYINPUT111), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  AND2_X1   g552(.A1(new_n691), .A2(new_n649), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n738), .A2(new_n721), .A3(new_n644), .A4(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G122), .ZN(G24));
  NAND2_X1  g555(.A1(new_n701), .A2(KEYINPUT112), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT112), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n627), .A2(new_n743), .A3(new_n639), .A4(new_n673), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n610), .B(new_n667), .C1(new_n735), .C2(new_n291), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n747), .A2(new_n712), .A3(new_n515), .A4(new_n644), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G125), .ZN(G27));
  INV_X1    g563(.A(KEYINPUT42), .ZN(new_n750));
  INV_X1    g564(.A(new_n508), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n516), .A2(new_n512), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n558), .A2(KEYINPUT113), .A3(new_n538), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT113), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n548), .B1(new_n529), .B2(new_n531), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n755), .B1(new_n756), .B2(new_n542), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n550), .A2(new_n534), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n754), .A2(new_n757), .A3(G469), .A4(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(new_n557), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n753), .B1(new_n761), .B2(new_n556), .ZN(new_n762));
  AND4_X1   g576(.A1(new_n750), .A2(new_n762), .A3(new_n742), .A4(new_n744), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n763), .A2(new_n602), .A3(new_n308), .A4(new_n606), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n602), .B1(new_n301), .B2(new_n307), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n762), .A2(new_n742), .A3(new_n744), .ZN(new_n766));
  OAI21_X1  g580(.A(KEYINPUT42), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n764), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(new_n212), .ZN(G33));
  AND2_X1   g583(.A1(new_n762), .A2(new_n674), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n308), .A2(new_n770), .A3(new_n602), .A4(new_n606), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G134), .ZN(G36));
  NAND2_X1  g586(.A1(new_n751), .A2(new_n509), .ZN(new_n773));
  INV_X1    g587(.A(new_n627), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n774), .A2(new_n639), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(KEYINPUT43), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n776), .A2(new_n612), .A3(new_n667), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT44), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n773), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n779), .B1(new_n778), .B2(new_n777), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n754), .A2(new_n757), .A3(KEYINPUT45), .A4(new_n758), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n781), .B(G469), .C1(new_n559), .C2(KEYINPUT45), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(new_n760), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT46), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n556), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n783), .A2(new_n784), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n515), .B(new_n679), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n780), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(new_n210), .ZN(G39));
  OAI21_X1  g604(.A(new_n515), .B1(new_n786), .B2(new_n787), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT114), .ZN(new_n792));
  AOI22_X1  g606(.A1(new_n791), .A2(new_n792), .B1(KEYINPUT115), .B2(KEYINPUT47), .ZN(new_n793));
  OAI211_X1 g607(.A(KEYINPUT114), .B(new_n515), .C1(new_n786), .C2(new_n787), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(KEYINPUT115), .A2(KEYINPUT47), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n795), .A2(new_n796), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n702), .A2(new_n601), .A3(new_n509), .A4(new_n751), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n800), .B1(new_n308), .B2(new_n606), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G140), .ZN(G42));
  OAI21_X1  g617(.A(new_n607), .B1(new_n706), .B2(new_n713), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n804), .A2(new_n718), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n764), .A2(new_n767), .A3(new_n771), .ZN(new_n806));
  INV_X1    g620(.A(new_n649), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n648), .A2(new_n384), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n807), .B1(new_n640), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n510), .A2(new_n513), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n613), .A2(new_n809), .A3(new_n561), .A4(new_n810), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n669), .A2(new_n811), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n812), .A2(new_n740), .A3(new_n723), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n667), .A2(new_n384), .A3(new_n673), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n814), .A2(new_n773), .A3(new_n648), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n308), .A2(new_n606), .A3(new_n561), .A4(new_n815), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n766), .A2(new_n746), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n805), .A2(new_n806), .A3(new_n813), .A4(new_n819), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n748), .A2(new_n677), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT52), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n691), .A2(new_n644), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n761), .A2(new_n556), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n665), .A2(new_n515), .A3(new_n673), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n823), .A2(new_n687), .A3(new_n824), .A4(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n821), .A2(new_n822), .A3(new_n704), .A4(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n704), .A2(new_n748), .A3(new_n677), .A4(new_n826), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(KEYINPUT52), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n748), .A2(new_n677), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n831), .B1(new_n832), .B2(KEYINPUT52), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n820), .A2(new_n830), .A3(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n831), .B1(new_n820), .B2(new_n830), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT116), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI211_X1 g652(.A(KEYINPUT116), .B(new_n831), .C1(new_n820), .C2(new_n830), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n835), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT54), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n812), .A2(new_n740), .A3(new_n723), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n843), .A2(new_n804), .A3(new_n718), .ZN(new_n844));
  INV_X1    g658(.A(new_n771), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n768), .A2(new_n845), .A3(new_n818), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n844), .A2(new_n846), .A3(new_n829), .A4(new_n827), .ZN(new_n847));
  AOI21_X1  g661(.A(KEYINPUT53), .B1(new_n832), .B2(KEYINPUT52), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n836), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(KEYINPUT54), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n842), .A2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n443), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n776), .A2(new_n852), .A3(new_n738), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n721), .A2(new_n512), .A3(new_n690), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n855), .A2(KEYINPUT50), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n855), .A2(KEYINPUT50), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n712), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n797), .B(new_n798), .C1(new_n515), .C2(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n853), .A2(new_n773), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n858), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n776), .A2(new_n852), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n863), .A2(new_n859), .A3(new_n753), .ZN(new_n864));
  INV_X1    g678(.A(new_n746), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n688), .A2(new_n602), .A3(new_n852), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n859), .A2(new_n867), .A3(new_n753), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n868), .A2(new_n384), .A3(new_n774), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(KEYINPUT51), .B1(new_n870), .B2(KEYINPUT117), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n871), .B1(KEYINPUT117), .B2(new_n870), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n862), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(new_n870), .ZN(new_n874));
  AOI21_X1  g688(.A(KEYINPUT51), .B1(new_n862), .B2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n765), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n864), .A2(new_n876), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n877), .B(KEYINPUT48), .Z(new_n878));
  NAND3_X1  g692(.A1(new_n868), .A2(new_n639), .A3(new_n627), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n721), .A2(new_n644), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n879), .B(new_n440), .C1(new_n881), .C2(new_n853), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n878), .A2(new_n882), .ZN(new_n883));
  NOR4_X1   g697(.A1(new_n851), .A2(new_n873), .A3(new_n875), .A4(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(G952), .A2(G953), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n859), .A2(KEYINPUT49), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n775), .A2(new_n602), .A3(new_n752), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n887), .A2(new_n687), .A3(new_n689), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT49), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n888), .B1(new_n889), .B2(new_n712), .ZN(new_n890));
  OAI22_X1  g704(.A1(new_n884), .A2(new_n885), .B1(new_n886), .B2(new_n890), .ZN(G75));
  NAND2_X1  g705(.A1(new_n477), .A2(new_n479), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(new_n491), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT55), .Z(new_n894));
  NOR3_X1   g708(.A1(new_n840), .A2(new_n269), .A3(new_n449), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n894), .B1(new_n895), .B2(KEYINPUT56), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT56), .ZN(new_n897));
  INV_X1    g711(.A(new_n894), .ZN(new_n898));
  INV_X1    g712(.A(new_n835), .ZN(new_n899));
  INV_X1    g713(.A(new_n839), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT116), .B1(new_n847), .B2(new_n831), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n270), .ZN(new_n903));
  OAI211_X1 g717(.A(new_n897), .B(new_n898), .C1(new_n903), .C2(new_n449), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n322), .A2(G952), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n896), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT118), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n896), .A2(KEYINPUT118), .A3(new_n904), .A4(new_n906), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(G51));
  NOR2_X1   g725(.A1(new_n903), .A2(new_n782), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n557), .B(KEYINPUT57), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n838), .A2(new_n839), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n841), .B1(new_n914), .B2(new_n899), .ZN(new_n915));
  AOI211_X1 g729(.A(KEYINPUT54), .B(new_n835), .C1(new_n838), .C2(new_n839), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n913), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n912), .B1(new_n917), .B2(new_n554), .ZN(new_n918));
  OAI21_X1  g732(.A(KEYINPUT119), .B1(new_n918), .B2(new_n905), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT119), .ZN(new_n920));
  INV_X1    g734(.A(new_n554), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n902), .A2(KEYINPUT54), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(new_n842), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n921), .B1(new_n923), .B2(new_n913), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n920), .B(new_n906), .C1(new_n924), .C2(new_n912), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n919), .A2(new_n925), .ZN(G54));
  AND2_X1   g740(.A1(KEYINPUT58), .A2(G475), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n902), .A2(new_n270), .A3(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(new_n637), .ZN(new_n929));
  OAI21_X1  g743(.A(KEYINPUT120), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n905), .B1(new_n928), .B2(new_n929), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n840), .A2(new_n269), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT120), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n932), .A2(new_n933), .A3(new_n637), .A4(new_n927), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n930), .A2(new_n931), .A3(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT121), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n930), .A2(new_n931), .A3(new_n934), .A4(KEYINPUT121), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(G60));
  NAND2_X1  g753(.A1(G478), .A2(G902), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT59), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n923), .A2(new_n699), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n699), .B1(new_n851), .B2(new_n941), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n942), .A2(new_n943), .A3(new_n905), .ZN(G63));
  NAND2_X1  g758(.A1(G217), .A2(G902), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT60), .Z(new_n946));
  NAND2_X1  g760(.A1(new_n902), .A2(new_n946), .ZN(new_n947));
  OR2_X1    g761(.A1(new_n947), .A2(new_n661), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n947), .A2(new_n589), .A3(new_n596), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n948), .A2(new_n906), .A3(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n948), .A2(KEYINPUT61), .A3(new_n906), .A4(new_n949), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(G66));
  XNOR2_X1  g768(.A(new_n844), .B(KEYINPUT122), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n322), .ZN(new_n956));
  OAI21_X1  g770(.A(G953), .B1(new_n486), .B2(new_n444), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n892), .B1(G898), .B2(new_n322), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n958), .B(new_n959), .ZN(G69));
  AOI21_X1  g774(.A(new_n322), .B1(G227), .B2(G900), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n261), .A2(new_n263), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n369), .A2(new_n370), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n962), .B(new_n963), .Z(new_n964));
  AOI21_X1  g778(.A(new_n789), .B1(new_n799), .B2(new_n801), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n821), .A2(new_n704), .ZN(new_n966));
  OR3_X1    g780(.A1(new_n696), .A2(KEYINPUT62), .A3(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(KEYINPUT62), .B1(new_n696), .B2(new_n966), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n640), .A2(new_n808), .ZN(new_n969));
  OR4_X1    g783(.A1(new_n706), .A2(new_n680), .A3(new_n773), .A4(new_n969), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n965), .A2(new_n967), .A3(new_n968), .A4(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n964), .B1(new_n971), .B2(new_n322), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(KEYINPUT123), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n806), .B(KEYINPUT125), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n876), .A2(new_n823), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n976), .A2(new_n788), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n966), .A2(new_n977), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n965), .A2(new_n322), .A3(new_n975), .A4(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n964), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n980), .B1(G900), .B2(G953), .ZN(new_n981));
  AOI21_X1  g795(.A(KEYINPUT124), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n982), .B1(new_n972), .B2(KEYINPUT123), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n961), .B1(new_n974), .B2(new_n983), .ZN(new_n984));
  OR2_X1    g798(.A1(new_n972), .A2(KEYINPUT123), .ZN(new_n985));
  INV_X1    g799(.A(new_n961), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n985), .A2(new_n986), .A3(new_n973), .A4(new_n982), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n984), .A2(new_n987), .ZN(G72));
  XOR2_X1   g802(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n989));
  NAND2_X1  g803(.A1(G472), .A2(G902), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n989), .B(new_n990), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT127), .Z(new_n992));
  OAI21_X1  g806(.A(new_n992), .B1(new_n971), .B2(new_n955), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n993), .A2(new_n254), .A3(new_n265), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n965), .A2(new_n975), .A3(new_n978), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n992), .B1(new_n995), .B2(new_n955), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n996), .A2(new_n255), .A3(new_n266), .A4(new_n264), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n265), .A2(new_n266), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n991), .B1(new_n998), .B2(new_n285), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n905), .B1(new_n849), .B2(new_n999), .ZN(new_n1000));
  AND3_X1   g814(.A1(new_n994), .A2(new_n997), .A3(new_n1000), .ZN(G57));
endmodule


