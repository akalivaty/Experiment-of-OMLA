

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585;

  XNOR2_X1 U319 ( .A(n411), .B(KEYINPUT54), .ZN(n412) );
  XNOR2_X1 U320 ( .A(KEYINPUT26), .B(KEYINPUT95), .ZN(n446) );
  XNOR2_X1 U321 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U322 ( .A(n335), .B(n334), .ZN(n339) );
  NOR2_X1 U323 ( .A1(n393), .A2(n392), .ZN(n394) );
  XNOR2_X1 U324 ( .A(n385), .B(n384), .ZN(n393) );
  XNOR2_X1 U325 ( .A(n448), .B(KEYINPUT123), .ZN(n581) );
  XNOR2_X1 U326 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U327 ( .A(n426), .B(n425), .ZN(n535) );
  XOR2_X1 U328 ( .A(KEYINPUT93), .B(n473), .Z(n522) );
  XOR2_X1 U329 ( .A(n419), .B(n330), .Z(n287) );
  NOR2_X1 U330 ( .A1(n389), .A2(n388), .ZN(n390) );
  INV_X1 U331 ( .A(KEYINPUT79), .ZN(n314) );
  XNOR2_X1 U332 ( .A(KEYINPUT109), .B(KEYINPUT47), .ZN(n384) );
  XNOR2_X1 U333 ( .A(n315), .B(n314), .ZN(n317) );
  XNOR2_X1 U334 ( .A(n347), .B(n346), .ZN(n348) );
  INV_X1 U335 ( .A(KEYINPUT29), .ZN(n332) );
  XNOR2_X1 U336 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U337 ( .A(n317), .B(n316), .ZN(n416) );
  XNOR2_X1 U338 ( .A(n427), .B(n348), .ZN(n349) );
  XNOR2_X1 U339 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U340 ( .A(n476), .B(KEYINPUT96), .ZN(n491) );
  XNOR2_X1 U341 ( .A(n447), .B(n446), .ZN(n553) );
  INV_X1 U342 ( .A(n491), .ZN(n494) );
  AND2_X1 U343 ( .A1(n455), .A2(n468), .ZN(n448) );
  XNOR2_X1 U344 ( .A(n382), .B(n381), .ZN(n386) );
  INV_X1 U345 ( .A(G218GAT), .ZN(n452) );
  INV_X1 U346 ( .A(G29GAT), .ZN(n481) );
  XNOR2_X1 U347 ( .A(n452), .B(KEYINPUT62), .ZN(n453) );
  XNOR2_X1 U348 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U349 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U350 ( .A(n454), .B(n453), .ZN(G1355GAT) );
  XNOR2_X1 U351 ( .A(n488), .B(n487), .ZN(G1351GAT) );
  XNOR2_X1 U352 ( .A(n484), .B(n483), .ZN(G1328GAT) );
  XOR2_X1 U353 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n289) );
  XNOR2_X1 U354 ( .A(G64GAT), .B(KEYINPUT15), .ZN(n288) );
  XNOR2_X1 U355 ( .A(n289), .B(n288), .ZN(n293) );
  XOR2_X1 U356 ( .A(KEYINPUT13), .B(KEYINPUT77), .Z(n291) );
  XNOR2_X1 U357 ( .A(KEYINPUT76), .B(KEYINPUT78), .ZN(n290) );
  XNOR2_X1 U358 ( .A(n291), .B(n290), .ZN(n292) );
  XNOR2_X1 U359 ( .A(n293), .B(n292), .ZN(n307) );
  XOR2_X1 U360 ( .A(G211GAT), .B(G78GAT), .Z(n295) );
  XNOR2_X1 U361 ( .A(G127GAT), .B(G71GAT), .ZN(n294) );
  XNOR2_X1 U362 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U363 ( .A(G57GAT), .B(G155GAT), .Z(n297) );
  XNOR2_X1 U364 ( .A(G1GAT), .B(G8GAT), .ZN(n296) );
  XNOR2_X1 U365 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U366 ( .A(n299), .B(n298), .Z(n305) );
  XNOR2_X1 U367 ( .A(G22GAT), .B(KEYINPUT70), .ZN(n300) );
  XNOR2_X1 U368 ( .A(n300), .B(KEYINPUT69), .ZN(n330) );
  XOR2_X1 U369 ( .A(G183GAT), .B(n330), .Z(n302) );
  NAND2_X1 U370 ( .A1(G231GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U371 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U372 ( .A(G15GAT), .B(n303), .ZN(n304) );
  XNOR2_X1 U373 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U374 ( .A(n307), .B(n306), .Z(n572) );
  INV_X1 U375 ( .A(n572), .ZN(n563) );
  XOR2_X1 U376 ( .A(KEYINPUT4), .B(KEYINPUT92), .Z(n309) );
  XNOR2_X1 U377 ( .A(KEYINPUT1), .B(KEYINPUT5), .ZN(n308) );
  XNOR2_X1 U378 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U379 ( .A(KEYINPUT91), .B(n310), .Z(n312) );
  NAND2_X1 U380 ( .A1(G225GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U381 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U382 ( .A(n313), .B(KEYINPUT6), .Z(n319) );
  XNOR2_X1 U383 ( .A(G127GAT), .B(G120GAT), .ZN(n315) );
  XOR2_X1 U384 ( .A(KEYINPUT0), .B(G134GAT), .Z(n316) );
  XNOR2_X1 U385 ( .A(n416), .B(KEYINPUT75), .ZN(n318) );
  XNOR2_X1 U386 ( .A(n319), .B(n318), .ZN(n321) );
  XNOR2_X1 U387 ( .A(G148GAT), .B(G85GAT), .ZN(n320) );
  XNOR2_X1 U388 ( .A(n320), .B(G57GAT), .ZN(n350) );
  XOR2_X1 U389 ( .A(n321), .B(n350), .Z(n329) );
  XOR2_X1 U390 ( .A(G1GAT), .B(G141GAT), .Z(n323) );
  XNOR2_X1 U391 ( .A(G29GAT), .B(G113GAT), .ZN(n322) );
  XNOR2_X1 U392 ( .A(n323), .B(n322), .ZN(n342) );
  XNOR2_X1 U393 ( .A(KEYINPUT87), .B(KEYINPUT2), .ZN(n324) );
  XNOR2_X1 U394 ( .A(n324), .B(KEYINPUT3), .ZN(n325) );
  XOR2_X1 U395 ( .A(n325), .B(KEYINPUT86), .Z(n327) );
  XNOR2_X1 U396 ( .A(G155GAT), .B(G162GAT), .ZN(n326) );
  XNOR2_X1 U397 ( .A(n327), .B(n326), .ZN(n431) );
  XNOR2_X1 U398 ( .A(n342), .B(n431), .ZN(n328) );
  XNOR2_X1 U399 ( .A(n329), .B(n328), .ZN(n473) );
  INV_X1 U400 ( .A(KEYINPUT48), .ZN(n395) );
  XOR2_X1 U401 ( .A(G43GAT), .B(G15GAT), .Z(n419) );
  NAND2_X1 U402 ( .A1(G229GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U403 ( .A(n287), .B(n331), .ZN(n335) );
  XOR2_X1 U404 ( .A(G197GAT), .B(G8GAT), .Z(n408) );
  XNOR2_X1 U405 ( .A(G169GAT), .B(n408), .ZN(n333) );
  XOR2_X1 U406 ( .A(KEYINPUT30), .B(KEYINPUT66), .Z(n337) );
  XNOR2_X1 U407 ( .A(KEYINPUT67), .B(KEYINPUT68), .ZN(n336) );
  XNOR2_X1 U408 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U409 ( .A(n339), .B(n338), .Z(n344) );
  XOR2_X1 U410 ( .A(G36GAT), .B(G50GAT), .Z(n341) );
  XNOR2_X1 U411 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n340) );
  XNOR2_X1 U412 ( .A(n341), .B(n340), .ZN(n376) );
  XNOR2_X1 U413 ( .A(n376), .B(n342), .ZN(n343) );
  XNOR2_X1 U414 ( .A(n344), .B(n343), .ZN(n576) );
  XNOR2_X1 U415 ( .A(G106GAT), .B(G78GAT), .ZN(n345) );
  XNOR2_X1 U416 ( .A(n345), .B(KEYINPUT73), .ZN(n427) );
  NAND2_X1 U417 ( .A1(G230GAT), .A2(G233GAT), .ZN(n347) );
  INV_X1 U418 ( .A(KEYINPUT74), .ZN(n346) );
  XOR2_X1 U419 ( .A(G92GAT), .B(G64GAT), .Z(n401) );
  XNOR2_X1 U420 ( .A(n349), .B(n401), .ZN(n352) );
  XOR2_X1 U421 ( .A(G99GAT), .B(G71GAT), .Z(n415) );
  XOR2_X1 U422 ( .A(n415), .B(n350), .Z(n351) );
  XNOR2_X1 U423 ( .A(n352), .B(n351), .ZN(n360) );
  XOR2_X1 U424 ( .A(KEYINPUT13), .B(G204GAT), .Z(n354) );
  XNOR2_X1 U425 ( .A(G176GAT), .B(G120GAT), .ZN(n353) );
  XNOR2_X1 U426 ( .A(n354), .B(n353), .ZN(n358) );
  XOR2_X1 U427 ( .A(KEYINPUT72), .B(KEYINPUT31), .Z(n356) );
  XNOR2_X1 U428 ( .A(KEYINPUT33), .B(KEYINPUT32), .ZN(n355) );
  XNOR2_X1 U429 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U430 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U431 ( .A(n360), .B(n359), .ZN(n580) );
  XOR2_X1 U432 ( .A(KEYINPUT41), .B(n580), .Z(n560) );
  NOR2_X1 U433 ( .A1(n576), .A2(n560), .ZN(n361) );
  XNOR2_X1 U434 ( .A(n361), .B(KEYINPUT46), .ZN(n362) );
  NOR2_X1 U435 ( .A1(n572), .A2(n362), .ZN(n364) );
  INV_X1 U436 ( .A(KEYINPUT108), .ZN(n363) );
  XNOR2_X1 U437 ( .A(n364), .B(n363), .ZN(n383) );
  XOR2_X1 U438 ( .A(G85GAT), .B(G99GAT), .Z(n366) );
  XNOR2_X1 U439 ( .A(G29GAT), .B(G43GAT), .ZN(n365) );
  XNOR2_X1 U440 ( .A(n366), .B(n365), .ZN(n368) );
  XOR2_X1 U441 ( .A(G106GAT), .B(G218GAT), .Z(n367) );
  XNOR2_X1 U442 ( .A(n368), .B(n367), .ZN(n374) );
  XOR2_X1 U443 ( .A(KEYINPUT10), .B(KEYINPUT65), .Z(n370) );
  XNOR2_X1 U444 ( .A(KEYINPUT75), .B(G92GAT), .ZN(n369) );
  XNOR2_X1 U445 ( .A(n370), .B(n369), .ZN(n372) );
  NAND2_X1 U446 ( .A1(G232GAT), .A2(G233GAT), .ZN(n371) );
  XOR2_X1 U447 ( .A(n375), .B(G162GAT), .Z(n382) );
  XNOR2_X1 U448 ( .A(n376), .B(G134GAT), .ZN(n380) );
  XOR2_X1 U449 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n378) );
  XNOR2_X1 U450 ( .A(G190GAT), .B(KEYINPUT64), .ZN(n377) );
  XNOR2_X1 U451 ( .A(n378), .B(n377), .ZN(n379) );
  NOR2_X1 U452 ( .A1(n383), .A2(n386), .ZN(n385) );
  XNOR2_X1 U453 ( .A(n576), .B(KEYINPUT71), .ZN(n569) );
  INV_X1 U454 ( .A(n580), .ZN(n389) );
  XOR2_X1 U455 ( .A(n386), .B(KEYINPUT36), .Z(n477) );
  NOR2_X1 U456 ( .A1(n563), .A2(n477), .ZN(n387) );
  XOR2_X1 U457 ( .A(KEYINPUT45), .B(n387), .Z(n388) );
  XOR2_X1 U458 ( .A(KEYINPUT110), .B(n390), .Z(n391) );
  NOR2_X1 U459 ( .A1(n569), .A2(n391), .ZN(n392) );
  XNOR2_X1 U460 ( .A(n395), .B(n394), .ZN(n551) );
  XOR2_X1 U461 ( .A(KEYINPUT21), .B(G218GAT), .Z(n397) );
  XNOR2_X1 U462 ( .A(G211GAT), .B(G204GAT), .ZN(n396) );
  XNOR2_X1 U463 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U464 ( .A(KEYINPUT85), .B(n398), .Z(n434) );
  XOR2_X1 U465 ( .A(n434), .B(G36GAT), .Z(n400) );
  NAND2_X1 U466 ( .A1(G226GAT), .A2(G233GAT), .ZN(n399) );
  XNOR2_X1 U467 ( .A(n400), .B(n399), .ZN(n402) );
  XOR2_X1 U468 ( .A(n402), .B(n401), .Z(n410) );
  XOR2_X1 U469 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n404) );
  XNOR2_X1 U470 ( .A(G190GAT), .B(KEYINPUT17), .ZN(n403) );
  XNOR2_X1 U471 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U472 ( .A(n405), .B(G183GAT), .Z(n407) );
  XNOR2_X1 U473 ( .A(G169GAT), .B(G176GAT), .ZN(n406) );
  XNOR2_X1 U474 ( .A(n407), .B(n406), .ZN(n426) );
  XNOR2_X1 U475 ( .A(n408), .B(n426), .ZN(n409) );
  XOR2_X1 U476 ( .A(n410), .B(n409), .Z(n524) );
  AND2_X1 U477 ( .A1(n551), .A2(n524), .ZN(n413) );
  INV_X1 U478 ( .A(KEYINPUT118), .ZN(n411) );
  XNOR2_X1 U479 ( .A(n413), .B(n412), .ZN(n414) );
  NOR2_X1 U480 ( .A1(n522), .A2(n414), .ZN(n455) );
  XOR2_X1 U481 ( .A(n415), .B(KEYINPUT20), .Z(n418) );
  XNOR2_X1 U482 ( .A(n416), .B(KEYINPUT81), .ZN(n417) );
  XNOR2_X1 U483 ( .A(n418), .B(n417), .ZN(n424) );
  XOR2_X1 U484 ( .A(KEYINPUT80), .B(n419), .Z(n421) );
  NAND2_X1 U485 ( .A1(G227GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U486 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U487 ( .A(G113GAT), .B(n422), .Z(n423) );
  XNOR2_X1 U488 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U489 ( .A(n427), .B(G141GAT), .Z(n429) );
  NAND2_X1 U490 ( .A1(G228GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U491 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U492 ( .A(n431), .B(n430), .ZN(n445) );
  XOR2_X1 U493 ( .A(KEYINPUT84), .B(KEYINPUT89), .Z(n433) );
  XNOR2_X1 U494 ( .A(KEYINPUT22), .B(G148GAT), .ZN(n432) );
  XNOR2_X1 U495 ( .A(n433), .B(n432), .ZN(n435) );
  XOR2_X1 U496 ( .A(n435), .B(n434), .Z(n443) );
  XOR2_X1 U497 ( .A(KEYINPUT88), .B(KEYINPUT83), .Z(n437) );
  XNOR2_X1 U498 ( .A(G197GAT), .B(KEYINPUT24), .ZN(n436) );
  XNOR2_X1 U499 ( .A(n437), .B(n436), .ZN(n441) );
  XOR2_X1 U500 ( .A(KEYINPUT90), .B(KEYINPUT23), .Z(n439) );
  XNOR2_X1 U501 ( .A(G50GAT), .B(G22GAT), .ZN(n438) );
  XNOR2_X1 U502 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U503 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U504 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U505 ( .A(n445), .B(n444), .ZN(n466) );
  NOR2_X1 U506 ( .A1(n535), .A2(n466), .ZN(n447) );
  INV_X1 U507 ( .A(n553), .ZN(n468) );
  NOR2_X1 U508 ( .A1(n563), .A2(n581), .ZN(n451) );
  INV_X1 U509 ( .A(G211GAT), .ZN(n449) );
  XNOR2_X1 U510 ( .A(n449), .B(KEYINPUT126), .ZN(n450) );
  XNOR2_X1 U511 ( .A(n451), .B(n450), .ZN(G1354GAT) );
  NOR2_X1 U512 ( .A1(n477), .A2(n581), .ZN(n454) );
  NAND2_X1 U513 ( .A1(n466), .A2(n455), .ZN(n456) );
  XNOR2_X1 U514 ( .A(n456), .B(KEYINPUT55), .ZN(n457) );
  NAND2_X1 U515 ( .A1(n457), .A2(n535), .ZN(n458) );
  XNOR2_X1 U516 ( .A(n458), .B(KEYINPUT119), .ZN(n573) );
  INV_X1 U517 ( .A(n560), .ZN(n541) );
  NAND2_X1 U518 ( .A1(n573), .A2(n541), .ZN(n461) );
  XOR2_X1 U519 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n459) );
  XNOR2_X1 U520 ( .A(n459), .B(G176GAT), .ZN(n460) );
  XNOR2_X1 U521 ( .A(n461), .B(n460), .ZN(G1349GAT) );
  XNOR2_X1 U522 ( .A(n524), .B(KEYINPUT27), .ZN(n469) );
  NAND2_X1 U523 ( .A1(n469), .A2(n522), .ZN(n462) );
  XOR2_X1 U524 ( .A(KEYINPUT94), .B(n462), .Z(n554) );
  XOR2_X1 U525 ( .A(n466), .B(KEYINPUT28), .Z(n530) );
  INV_X1 U526 ( .A(n530), .ZN(n463) );
  NAND2_X1 U527 ( .A1(n554), .A2(n463), .ZN(n537) );
  XNOR2_X1 U528 ( .A(KEYINPUT82), .B(n535), .ZN(n464) );
  NOR2_X1 U529 ( .A1(n537), .A2(n464), .ZN(n475) );
  NAND2_X1 U530 ( .A1(n535), .A2(n524), .ZN(n465) );
  NAND2_X1 U531 ( .A1(n466), .A2(n465), .ZN(n467) );
  XNOR2_X1 U532 ( .A(n467), .B(KEYINPUT25), .ZN(n471) );
  AND2_X1 U533 ( .A1(n469), .A2(n468), .ZN(n470) );
  NOR2_X1 U534 ( .A1(n471), .A2(n470), .ZN(n472) );
  NOR2_X1 U535 ( .A1(n473), .A2(n472), .ZN(n474) );
  NOR2_X1 U536 ( .A1(n475), .A2(n474), .ZN(n476) );
  NOR2_X1 U537 ( .A1(n491), .A2(n477), .ZN(n478) );
  NAND2_X1 U538 ( .A1(n478), .A2(n563), .ZN(n479) );
  XOR2_X1 U539 ( .A(KEYINPUT37), .B(n479), .Z(n521) );
  NAND2_X1 U540 ( .A1(n580), .A2(n569), .ZN(n495) );
  NOR2_X1 U541 ( .A1(n521), .A2(n495), .ZN(n480) );
  XNOR2_X1 U542 ( .A(KEYINPUT38), .B(n480), .ZN(n507) );
  NAND2_X1 U543 ( .A1(n522), .A2(n507), .ZN(n484) );
  XOR2_X1 U544 ( .A(KEYINPUT99), .B(KEYINPUT39), .Z(n482) );
  NAND2_X1 U545 ( .A1(n573), .A2(n386), .ZN(n488) );
  XOR2_X1 U546 ( .A(KEYINPUT122), .B(KEYINPUT58), .Z(n486) );
  INV_X1 U547 ( .A(G190GAT), .ZN(n485) );
  XNOR2_X1 U548 ( .A(G1GAT), .B(KEYINPUT98), .ZN(n489) );
  XNOR2_X1 U549 ( .A(n489), .B(KEYINPUT97), .ZN(n490) );
  XOR2_X1 U550 ( .A(KEYINPUT34), .B(n490), .Z(n497) );
  NOR2_X1 U551 ( .A1(n386), .A2(n563), .ZN(n492) );
  XNOR2_X1 U552 ( .A(n492), .B(KEYINPUT16), .ZN(n493) );
  NAND2_X1 U553 ( .A1(n494), .A2(n493), .ZN(n510) );
  NOR2_X1 U554 ( .A1(n495), .A2(n510), .ZN(n501) );
  NAND2_X1 U555 ( .A1(n501), .A2(n522), .ZN(n496) );
  XNOR2_X1 U556 ( .A(n497), .B(n496), .ZN(G1324GAT) );
  NAND2_X1 U557 ( .A1(n524), .A2(n501), .ZN(n498) );
  XNOR2_X1 U558 ( .A(n498), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U559 ( .A(G15GAT), .B(KEYINPUT35), .Z(n500) );
  NAND2_X1 U560 ( .A1(n501), .A2(n535), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n500), .B(n499), .ZN(G1326GAT) );
  NAND2_X1 U562 ( .A1(n501), .A2(n530), .ZN(n502) );
  XNOR2_X1 U563 ( .A(n502), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U564 ( .A1(n507), .A2(n524), .ZN(n503) );
  XNOR2_X1 U565 ( .A(n503), .B(KEYINPUT100), .ZN(n504) );
  XNOR2_X1 U566 ( .A(G36GAT), .B(n504), .ZN(G1329GAT) );
  NAND2_X1 U567 ( .A1(n507), .A2(n535), .ZN(n505) );
  XNOR2_X1 U568 ( .A(n505), .B(KEYINPUT40), .ZN(n506) );
  XNOR2_X1 U569 ( .A(G43GAT), .B(n506), .ZN(G1330GAT) );
  XOR2_X1 U570 ( .A(G50GAT), .B(KEYINPUT101), .Z(n509) );
  NAND2_X1 U571 ( .A1(n530), .A2(n507), .ZN(n508) );
  XNOR2_X1 U572 ( .A(n509), .B(n508), .ZN(G1331GAT) );
  XOR2_X1 U573 ( .A(KEYINPUT42), .B(KEYINPUT102), .Z(n512) );
  NAND2_X1 U574 ( .A1(n576), .A2(n541), .ZN(n520) );
  NOR2_X1 U575 ( .A1(n520), .A2(n510), .ZN(n516) );
  NAND2_X1 U576 ( .A1(n516), .A2(n522), .ZN(n511) );
  XNOR2_X1 U577 ( .A(n512), .B(n511), .ZN(n513) );
  XOR2_X1 U578 ( .A(G57GAT), .B(n513), .Z(G1332GAT) );
  NAND2_X1 U579 ( .A1(n524), .A2(n516), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n514), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U581 ( .A1(n516), .A2(n535), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n515), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U583 ( .A(KEYINPUT103), .B(KEYINPUT43), .Z(n518) );
  NAND2_X1 U584 ( .A1(n516), .A2(n530), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n518), .B(n517), .ZN(n519) );
  XOR2_X1 U586 ( .A(G78GAT), .B(n519), .Z(G1335GAT) );
  NOR2_X1 U587 ( .A1(n521), .A2(n520), .ZN(n531) );
  NAND2_X1 U588 ( .A1(n522), .A2(n531), .ZN(n523) );
  XNOR2_X1 U589 ( .A(G85GAT), .B(n523), .ZN(G1336GAT) );
  NAND2_X1 U590 ( .A1(n524), .A2(n531), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n525), .B(KEYINPUT104), .ZN(n526) );
  XNOR2_X1 U592 ( .A(G92GAT), .B(n526), .ZN(G1337GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n528) );
  NAND2_X1 U594 ( .A1(n531), .A2(n535), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U596 ( .A(G99GAT), .B(n529), .ZN(G1338GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT44), .B(KEYINPUT107), .Z(n533) );
  NAND2_X1 U598 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U600 ( .A(G106GAT), .B(n534), .ZN(G1339GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n539) );
  NAND2_X1 U602 ( .A1(n535), .A2(n551), .ZN(n536) );
  NOR2_X1 U603 ( .A1(n537), .A2(n536), .ZN(n548) );
  NAND2_X1 U604 ( .A1(n548), .A2(n569), .ZN(n538) );
  XNOR2_X1 U605 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U606 ( .A(G113GAT), .B(n540), .ZN(G1340GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT113), .B(KEYINPUT49), .Z(n543) );
  NAND2_X1 U608 ( .A1(n548), .A2(n541), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U610 ( .A(G120GAT), .B(n544), .Z(G1341GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n546) );
  NAND2_X1 U612 ( .A1(n548), .A2(n572), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U614 ( .A(G127GAT), .B(n547), .Z(G1342GAT) );
  XOR2_X1 U615 ( .A(G134GAT), .B(KEYINPUT51), .Z(n550) );
  NAND2_X1 U616 ( .A1(n548), .A2(n386), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  INV_X1 U618 ( .A(n551), .ZN(n552) );
  NOR2_X1 U619 ( .A1(n553), .A2(n552), .ZN(n555) );
  NAND2_X1 U620 ( .A1(n555), .A2(n554), .ZN(n566) );
  NOR2_X1 U621 ( .A1(n576), .A2(n566), .ZN(n557) );
  XNOR2_X1 U622 ( .A(G141GAT), .B(KEYINPUT115), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(G1344GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n559) );
  XNOR2_X1 U625 ( .A(G148GAT), .B(KEYINPUT116), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(n562) );
  NOR2_X1 U627 ( .A1(n560), .A2(n566), .ZN(n561) );
  XOR2_X1 U628 ( .A(n562), .B(n561), .Z(G1345GAT) );
  NOR2_X1 U629 ( .A1(n563), .A2(n566), .ZN(n565) );
  XNOR2_X1 U630 ( .A(G155GAT), .B(KEYINPUT117), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(G1346GAT) );
  INV_X1 U632 ( .A(n386), .ZN(n567) );
  NOR2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U634 ( .A(G162GAT), .B(n568), .Z(G1347GAT) );
  XNOR2_X1 U635 ( .A(G169GAT), .B(KEYINPUT120), .ZN(n571) );
  NAND2_X1 U636 ( .A1(n573), .A2(n569), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(G1348GAT) );
  XOR2_X1 U638 ( .A(G183GAT), .B(KEYINPUT121), .Z(n575) );
  NAND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1350GAT) );
  NOR2_X1 U641 ( .A1(n576), .A2(n581), .ZN(n578) );
  XNOR2_X1 U642 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(n579), .ZN(G1352GAT) );
  NOR2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n585) );
  XOR2_X1 U646 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n583) );
  XNOR2_X1 U647 ( .A(G204GAT), .B(KEYINPUT125), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(G1353GAT) );
endmodule

