

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591;

  XOR2_X2 U324 ( .A(KEYINPUT13), .B(KEYINPUT69), .Z(n346) );
  NOR2_X1 U325 ( .A1(n540), .A2(n555), .ZN(n433) );
  NOR2_X1 U326 ( .A1(n387), .A2(n568), .ZN(n388) );
  AND2_X1 U327 ( .A1(n558), .A2(n575), .ZN(n364) );
  XNOR2_X1 U328 ( .A(n313), .B(n312), .ZN(n314) );
  INV_X1 U329 ( .A(n353), .ZN(n318) );
  XNOR2_X1 U330 ( .A(n319), .B(n318), .ZN(n320) );
  INV_X1 U331 ( .A(n406), .ZN(n357) );
  XNOR2_X1 U332 ( .A(n321), .B(n320), .ZN(n323) );
  XNOR2_X1 U333 ( .A(n358), .B(n357), .ZN(n359) );
  NOR2_X1 U334 ( .A1(n583), .A2(n470), .ZN(n472) );
  AND2_X1 U335 ( .A1(n573), .A2(n485), .ZN(n486) );
  XNOR2_X1 U336 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U337 ( .A(n315), .B(n314), .ZN(n407) );
  XOR2_X1 U338 ( .A(n307), .B(n343), .Z(n575) );
  INV_X1 U339 ( .A(KEYINPUT108), .ZN(n478) );
  XNOR2_X1 U340 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U341 ( .A(G113GAT), .B(KEYINPUT118), .ZN(n453) );
  XNOR2_X1 U342 ( .A(n478), .B(G36GAT), .ZN(n479) );
  XNOR2_X1 U343 ( .A(n491), .B(n490), .ZN(G1349GAT) );
  XNOR2_X1 U344 ( .A(n480), .B(n479), .ZN(G1329GAT) );
  XNOR2_X1 U345 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n292) );
  XNOR2_X1 U346 ( .A(n292), .B(KEYINPUT8), .ZN(n370) );
  XOR2_X1 U347 ( .A(G50GAT), .B(n370), .Z(n294) );
  NAND2_X1 U348 ( .A1(G229GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U349 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U350 ( .A(n295), .B(G29GAT), .Z(n303) );
  XOR2_X1 U351 ( .A(G169GAT), .B(G141GAT), .Z(n297) );
  XNOR2_X1 U352 ( .A(G43GAT), .B(G197GAT), .ZN(n296) );
  XNOR2_X1 U353 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U354 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n299) );
  XNOR2_X1 U355 ( .A(G113GAT), .B(KEYINPUT67), .ZN(n298) );
  XNOR2_X1 U356 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U357 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U358 ( .A(n303), .B(n302), .ZN(n307) );
  XOR2_X1 U359 ( .A(G15GAT), .B(G22GAT), .Z(n305) );
  XNOR2_X1 U360 ( .A(KEYINPUT68), .B(G8GAT), .ZN(n304) );
  XNOR2_X1 U361 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U362 ( .A(G1GAT), .B(n306), .ZN(n343) );
  XOR2_X1 U363 ( .A(G43GAT), .B(G134GAT), .Z(n376) );
  XOR2_X1 U364 ( .A(KEYINPUT85), .B(KEYINPUT84), .Z(n309) );
  XNOR2_X1 U365 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n308) );
  XNOR2_X1 U366 ( .A(n309), .B(n308), .ZN(n311) );
  INV_X1 U367 ( .A(KEYINPUT19), .ZN(n310) );
  XNOR2_X1 U368 ( .A(n311), .B(n310), .ZN(n315) );
  XNOR2_X1 U369 ( .A(G169GAT), .B(G176GAT), .ZN(n313) );
  XNOR2_X1 U370 ( .A(G190GAT), .B(G183GAT), .ZN(n312) );
  XNOR2_X1 U371 ( .A(G15GAT), .B(n407), .ZN(n321) );
  XOR2_X1 U372 ( .A(G120GAT), .B(G127GAT), .Z(n317) );
  XNOR2_X1 U373 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n316) );
  XNOR2_X1 U374 ( .A(n317), .B(n316), .ZN(n416) );
  XOR2_X1 U375 ( .A(n416), .B(KEYINPUT20), .Z(n319) );
  XOR2_X1 U376 ( .A(G99GAT), .B(G71GAT), .Z(n353) );
  XNOR2_X1 U377 ( .A(KEYINPUT82), .B(KEYINPUT83), .ZN(n322) );
  XNOR2_X1 U378 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U379 ( .A(n376), .B(n324), .Z(n326) );
  NAND2_X1 U380 ( .A1(G227GAT), .A2(G233GAT), .ZN(n325) );
  XOR2_X1 U381 ( .A(n326), .B(n325), .Z(n507) );
  INV_X1 U382 ( .A(n507), .ZN(n540) );
  XOR2_X1 U383 ( .A(KEYINPUT79), .B(KEYINPUT14), .Z(n328) );
  XNOR2_X1 U384 ( .A(KEYINPUT81), .B(KEYINPUT12), .ZN(n327) );
  XNOR2_X1 U385 ( .A(n328), .B(n327), .ZN(n341) );
  XOR2_X1 U386 ( .A(G183GAT), .B(G78GAT), .Z(n330) );
  XNOR2_X1 U387 ( .A(G155GAT), .B(G211GAT), .ZN(n329) );
  XNOR2_X1 U388 ( .A(n330), .B(n329), .ZN(n334) );
  XOR2_X1 U389 ( .A(G57GAT), .B(G64GAT), .Z(n332) );
  XNOR2_X1 U390 ( .A(G71GAT), .B(G127GAT), .ZN(n331) );
  XNOR2_X1 U391 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U392 ( .A(n334), .B(n333), .Z(n339) );
  XOR2_X1 U393 ( .A(KEYINPUT15), .B(KEYINPUT80), .Z(n336) );
  NAND2_X1 U394 ( .A1(G231GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U395 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U396 ( .A(n346), .B(n337), .ZN(n338) );
  XNOR2_X1 U397 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U398 ( .A(n341), .B(n340), .Z(n342) );
  XOR2_X1 U399 ( .A(n343), .B(n342), .Z(n492) );
  INV_X1 U400 ( .A(n492), .ZN(n583) );
  XOR2_X1 U401 ( .A(KEYINPUT31), .B(KEYINPUT70), .Z(n345) );
  XNOR2_X1 U402 ( .A(G120GAT), .B(KEYINPUT32), .ZN(n344) );
  XNOR2_X1 U403 ( .A(n345), .B(n344), .ZN(n362) );
  XOR2_X1 U404 ( .A(G85GAT), .B(n346), .Z(n348) );
  XOR2_X1 U405 ( .A(G148GAT), .B(G57GAT), .Z(n413) );
  XNOR2_X1 U406 ( .A(G176GAT), .B(n413), .ZN(n347) );
  XNOR2_X1 U407 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U408 ( .A(KEYINPUT73), .B(KEYINPUT33), .Z(n350) );
  NAND2_X1 U409 ( .A1(G230GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U410 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U411 ( .A(n352), .B(n351), .ZN(n355) );
  XOR2_X1 U412 ( .A(n353), .B(KEYINPUT74), .Z(n354) );
  XNOR2_X1 U413 ( .A(n355), .B(n354), .ZN(n360) );
  XOR2_X1 U414 ( .A(G106GAT), .B(G78GAT), .Z(n436) );
  XOR2_X1 U415 ( .A(KEYINPUT71), .B(G92GAT), .Z(n381) );
  XNOR2_X1 U416 ( .A(n436), .B(n381), .ZN(n358) );
  XNOR2_X1 U417 ( .A(G204GAT), .B(G64GAT), .ZN(n356) );
  XNOR2_X1 U418 ( .A(n356), .B(KEYINPUT72), .ZN(n406) );
  XOR2_X1 U419 ( .A(n362), .B(n361), .Z(n389) );
  XOR2_X2 U420 ( .A(n389), .B(KEYINPUT41), .Z(n558) );
  XNOR2_X1 U421 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n363) );
  XNOR2_X1 U422 ( .A(n364), .B(n363), .ZN(n365) );
  NOR2_X1 U423 ( .A1(n583), .A2(n365), .ZN(n366) );
  XNOR2_X1 U424 ( .A(n366), .B(KEYINPUT113), .ZN(n387) );
  XOR2_X1 U425 ( .A(KEYINPUT78), .B(KEYINPUT76), .Z(n372) );
  XOR2_X1 U426 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n368) );
  XNOR2_X1 U427 ( .A(G162GAT), .B(KEYINPUT11), .ZN(n367) );
  XNOR2_X1 U428 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U429 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U430 ( .A(n372), .B(n371), .ZN(n380) );
  XOR2_X1 U431 ( .A(KEYINPUT65), .B(G99GAT), .Z(n374) );
  XNOR2_X1 U432 ( .A(G106GAT), .B(G190GAT), .ZN(n373) );
  XNOR2_X1 U433 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U434 ( .A(n375), .B(KEYINPUT77), .Z(n378) );
  XNOR2_X1 U435 ( .A(G218GAT), .B(n376), .ZN(n377) );
  XNOR2_X1 U436 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U437 ( .A(n380), .B(n379), .Z(n386) );
  XOR2_X1 U438 ( .A(G50GAT), .B(KEYINPUT75), .Z(n437) );
  XOR2_X1 U439 ( .A(G29GAT), .B(G85GAT), .Z(n417) );
  XOR2_X1 U440 ( .A(n417), .B(n381), .Z(n383) );
  NAND2_X1 U441 ( .A1(G232GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U442 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U443 ( .A(n437), .B(n384), .ZN(n385) );
  XNOR2_X1 U444 ( .A(n386), .B(n385), .ZN(n568) );
  XNOR2_X1 U445 ( .A(n388), .B(KEYINPUT47), .ZN(n395) );
  BUF_X1 U446 ( .A(n389), .Z(n579) );
  XNOR2_X1 U447 ( .A(KEYINPUT36), .B(n568), .ZN(n587) );
  NAND2_X1 U448 ( .A1(n587), .A2(n583), .ZN(n390) );
  XNOR2_X1 U449 ( .A(n390), .B(KEYINPUT45), .ZN(n391) );
  XNOR2_X1 U450 ( .A(n391), .B(KEYINPUT64), .ZN(n392) );
  NOR2_X1 U451 ( .A1(n579), .A2(n392), .ZN(n393) );
  INV_X1 U452 ( .A(n575), .ZN(n455) );
  NAND2_X1 U453 ( .A1(n393), .A2(n455), .ZN(n394) );
  NAND2_X1 U454 ( .A1(n395), .A2(n394), .ZN(n397) );
  XNOR2_X1 U455 ( .A(KEYINPUT114), .B(KEYINPUT48), .ZN(n396) );
  XNOR2_X1 U456 ( .A(n397), .B(n396), .ZN(n481) );
  XOR2_X1 U457 ( .A(G211GAT), .B(KEYINPUT21), .Z(n399) );
  XNOR2_X1 U458 ( .A(G197GAT), .B(G218GAT), .ZN(n398) );
  XNOR2_X1 U459 ( .A(n399), .B(n398), .ZN(n445) );
  XOR2_X1 U460 ( .A(n445), .B(KEYINPUT96), .Z(n401) );
  NAND2_X1 U461 ( .A1(G226GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U462 ( .A(n401), .B(n400), .ZN(n405) );
  XOR2_X1 U463 ( .A(KEYINPUT95), .B(G92GAT), .Z(n403) );
  XNOR2_X1 U464 ( .A(G8GAT), .B(G36GAT), .ZN(n402) );
  XNOR2_X1 U465 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U466 ( .A(n405), .B(n404), .Z(n409) );
  XNOR2_X1 U467 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U468 ( .A(n409), .B(n408), .Z(n538) );
  XNOR2_X1 U469 ( .A(n538), .B(KEYINPUT27), .ZN(n462) );
  XOR2_X1 U470 ( .A(KEYINPUT4), .B(KEYINPUT91), .Z(n411) );
  XNOR2_X1 U471 ( .A(G134GAT), .B(KEYINPUT93), .ZN(n410) );
  XNOR2_X1 U472 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U473 ( .A(n412), .B(KEYINPUT1), .Z(n415) );
  XNOR2_X1 U474 ( .A(G1GAT), .B(n413), .ZN(n414) );
  XNOR2_X1 U475 ( .A(n415), .B(n414), .ZN(n421) );
  XOR2_X1 U476 ( .A(n417), .B(n416), .Z(n419) );
  NAND2_X1 U477 ( .A1(G225GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U478 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U479 ( .A(n421), .B(n420), .Z(n430) );
  XNOR2_X1 U480 ( .A(G155GAT), .B(KEYINPUT88), .ZN(n422) );
  XNOR2_X1 U481 ( .A(n422), .B(KEYINPUT3), .ZN(n423) );
  XOR2_X1 U482 ( .A(n423), .B(KEYINPUT2), .Z(n425) );
  XNOR2_X1 U483 ( .A(G141GAT), .B(G162GAT), .ZN(n424) );
  XNOR2_X1 U484 ( .A(n425), .B(n424), .ZN(n449) );
  XOR2_X1 U485 ( .A(KEYINPUT90), .B(KEYINPUT5), .Z(n427) );
  XNOR2_X1 U486 ( .A(KEYINPUT6), .B(KEYINPUT92), .ZN(n426) );
  XNOR2_X1 U487 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U488 ( .A(n449), .B(n428), .ZN(n429) );
  XNOR2_X1 U489 ( .A(n430), .B(n429), .ZN(n466) );
  XOR2_X1 U490 ( .A(KEYINPUT94), .B(n466), .Z(n498) );
  INV_X1 U491 ( .A(n498), .ZN(n536) );
  NOR2_X1 U492 ( .A1(n462), .A2(n536), .ZN(n457) );
  NAND2_X1 U493 ( .A1(n481), .A2(n457), .ZN(n432) );
  INV_X1 U494 ( .A(KEYINPUT115), .ZN(n431) );
  XNOR2_X1 U495 ( .A(n432), .B(n431), .ZN(n555) );
  XNOR2_X1 U496 ( .A(n433), .B(KEYINPUT116), .ZN(n451) );
  XNOR2_X1 U497 ( .A(KEYINPUT66), .B(KEYINPUT28), .ZN(n450) );
  XOR2_X1 U498 ( .A(KEYINPUT89), .B(KEYINPUT23), .Z(n435) );
  XNOR2_X1 U499 ( .A(G22GAT), .B(G148GAT), .ZN(n434) );
  XNOR2_X1 U500 ( .A(n435), .B(n434), .ZN(n441) );
  XOR2_X1 U501 ( .A(G204GAT), .B(KEYINPUT24), .Z(n439) );
  XNOR2_X1 U502 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U503 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U504 ( .A(n441), .B(n440), .Z(n443) );
  NAND2_X1 U505 ( .A1(G228GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U506 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U507 ( .A(n444), .B(KEYINPUT87), .Z(n447) );
  XNOR2_X1 U508 ( .A(n445), .B(KEYINPUT22), .ZN(n446) );
  XNOR2_X1 U509 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U510 ( .A(n449), .B(n448), .ZN(n485) );
  XOR2_X1 U511 ( .A(n450), .B(n485), .Z(n512) );
  INV_X1 U512 ( .A(n512), .ZN(n543) );
  NAND2_X1 U513 ( .A1(n451), .A2(n543), .ZN(n452) );
  XNOR2_X2 U514 ( .A(n452), .B(KEYINPUT117), .ZN(n551) );
  NAND2_X1 U515 ( .A1(n575), .A2(n551), .ZN(n454) );
  XNOR2_X1 U516 ( .A(n454), .B(n453), .ZN(G1340GAT) );
  NOR2_X1 U517 ( .A1(n455), .A2(n579), .ZN(n496) );
  INV_X1 U518 ( .A(KEYINPUT37), .ZN(n471) );
  XOR2_X1 U519 ( .A(KEYINPUT86), .B(n540), .Z(n456) );
  NOR2_X1 U520 ( .A1(n512), .A2(n456), .ZN(n458) );
  NAND2_X1 U521 ( .A1(n458), .A2(n457), .ZN(n469) );
  INV_X1 U522 ( .A(n538), .ZN(n503) );
  NAND2_X1 U523 ( .A1(n503), .A2(n507), .ZN(n459) );
  NAND2_X1 U524 ( .A1(n485), .A2(n459), .ZN(n460) );
  XNOR2_X1 U525 ( .A(n460), .B(KEYINPUT25), .ZN(n464) );
  NOR2_X1 U526 ( .A1(n485), .A2(n507), .ZN(n461) );
  XOR2_X1 U527 ( .A(KEYINPUT26), .B(n461), .Z(n554) );
  NOR2_X1 U528 ( .A1(n462), .A2(n554), .ZN(n463) );
  NOR2_X1 U529 ( .A1(n464), .A2(n463), .ZN(n465) );
  XNOR2_X1 U530 ( .A(n465), .B(KEYINPUT97), .ZN(n467) );
  NAND2_X1 U531 ( .A1(n467), .A2(n466), .ZN(n468) );
  NAND2_X1 U532 ( .A1(n469), .A2(n468), .ZN(n494) );
  NAND2_X1 U533 ( .A1(n587), .A2(n494), .ZN(n470) );
  NAND2_X1 U534 ( .A1(n471), .A2(n472), .ZN(n475) );
  INV_X1 U535 ( .A(n472), .ZN(n473) );
  NAND2_X1 U536 ( .A1(KEYINPUT37), .A2(n473), .ZN(n474) );
  NAND2_X1 U537 ( .A1(n475), .A2(n474), .ZN(n535) );
  NAND2_X1 U538 ( .A1(n496), .A2(n535), .ZN(n477) );
  XOR2_X1 U539 ( .A(KEYINPUT38), .B(KEYINPUT107), .Z(n476) );
  XNOR2_X1 U540 ( .A(n477), .B(n476), .ZN(n522) );
  NOR2_X1 U541 ( .A1(n522), .A2(n538), .ZN(n480) );
  XOR2_X1 U542 ( .A(KEYINPUT121), .B(KEYINPUT54), .Z(n483) );
  NAND2_X1 U543 ( .A1(n481), .A2(n503), .ZN(n482) );
  XNOR2_X1 U544 ( .A(n483), .B(n482), .ZN(n484) );
  NOR2_X1 U545 ( .A1(n484), .A2(n498), .ZN(n573) );
  XNOR2_X1 U546 ( .A(n486), .B(KEYINPUT55), .ZN(n487) );
  NOR2_X2 U547 ( .A1(n540), .A2(n487), .ZN(n569) );
  NAND2_X1 U548 ( .A1(n569), .A2(n558), .ZN(n491) );
  XOR2_X1 U549 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n489) );
  XNOR2_X1 U550 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n488) );
  NOR2_X1 U551 ( .A1(n568), .A2(n492), .ZN(n493) );
  XNOR2_X1 U552 ( .A(KEYINPUT16), .B(n493), .ZN(n495) );
  AND2_X1 U553 ( .A1(n495), .A2(n494), .ZN(n525) );
  NAND2_X1 U554 ( .A1(n496), .A2(n525), .ZN(n497) );
  XOR2_X1 U555 ( .A(KEYINPUT98), .B(n497), .Z(n511) );
  NAND2_X1 U556 ( .A1(n511), .A2(n498), .ZN(n502) );
  XOR2_X1 U557 ( .A(KEYINPUT34), .B(KEYINPUT100), .Z(n500) );
  XNOR2_X1 U558 ( .A(G1GAT), .B(KEYINPUT99), .ZN(n499) );
  XNOR2_X1 U559 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U560 ( .A(n502), .B(n501), .ZN(G1324GAT) );
  XOR2_X1 U561 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n505) );
  NAND2_X1 U562 ( .A1(n503), .A2(n511), .ZN(n504) );
  XNOR2_X1 U563 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U564 ( .A(G8GAT), .B(n506), .ZN(G1325GAT) );
  XOR2_X1 U565 ( .A(KEYINPUT103), .B(KEYINPUT35), .Z(n509) );
  NAND2_X1 U566 ( .A1(n511), .A2(n507), .ZN(n508) );
  XNOR2_X1 U567 ( .A(n509), .B(n508), .ZN(n510) );
  XOR2_X1 U568 ( .A(G15GAT), .B(n510), .Z(G1326GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n514) );
  NAND2_X1 U570 ( .A1(n512), .A2(n511), .ZN(n513) );
  XNOR2_X1 U571 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U572 ( .A(G22GAT), .B(n515), .ZN(G1327GAT) );
  NOR2_X1 U573 ( .A1(n522), .A2(n536), .ZN(n517) );
  XNOR2_X1 U574 ( .A(KEYINPUT106), .B(KEYINPUT39), .ZN(n516) );
  XNOR2_X1 U575 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U576 ( .A(G29GAT), .B(n518), .ZN(G1328GAT) );
  XNOR2_X1 U577 ( .A(KEYINPUT40), .B(KEYINPUT109), .ZN(n520) );
  NOR2_X1 U578 ( .A1(n540), .A2(n522), .ZN(n519) );
  XNOR2_X1 U579 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U580 ( .A(G43GAT), .B(n521), .ZN(G1330GAT) );
  NOR2_X1 U581 ( .A1(n522), .A2(n543), .ZN(n523) );
  XOR2_X1 U582 ( .A(G50GAT), .B(n523), .Z(G1331GAT) );
  INV_X1 U583 ( .A(n558), .ZN(n524) );
  NOR2_X1 U584 ( .A1(n575), .A2(n524), .ZN(n534) );
  NAND2_X1 U585 ( .A1(n525), .A2(n534), .ZN(n530) );
  NOR2_X1 U586 ( .A1(n536), .A2(n530), .ZN(n526) );
  XOR2_X1 U587 ( .A(G57GAT), .B(n526), .Z(n527) );
  XNOR2_X1 U588 ( .A(KEYINPUT42), .B(n527), .ZN(G1332GAT) );
  NOR2_X1 U589 ( .A1(n538), .A2(n530), .ZN(n528) );
  XOR2_X1 U590 ( .A(G64GAT), .B(n528), .Z(G1333GAT) );
  NOR2_X1 U591 ( .A1(n540), .A2(n530), .ZN(n529) );
  XOR2_X1 U592 ( .A(G71GAT), .B(n529), .Z(G1334GAT) );
  NOR2_X1 U593 ( .A1(n543), .A2(n530), .ZN(n532) );
  XNOR2_X1 U594 ( .A(KEYINPUT110), .B(KEYINPUT43), .ZN(n531) );
  XNOR2_X1 U595 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U596 ( .A(G78GAT), .B(n533), .ZN(G1335GAT) );
  NAND2_X1 U597 ( .A1(n535), .A2(n534), .ZN(n542) );
  NOR2_X1 U598 ( .A1(n536), .A2(n542), .ZN(n537) );
  XOR2_X1 U599 ( .A(G85GAT), .B(n537), .Z(G1336GAT) );
  NOR2_X1 U600 ( .A1(n538), .A2(n542), .ZN(n539) );
  XOR2_X1 U601 ( .A(G92GAT), .B(n539), .Z(G1337GAT) );
  NOR2_X1 U602 ( .A1(n540), .A2(n542), .ZN(n541) );
  XOR2_X1 U603 ( .A(G99GAT), .B(n541), .Z(G1338GAT) );
  NOR2_X1 U604 ( .A1(n543), .A2(n542), .ZN(n545) );
  XNOR2_X1 U605 ( .A(KEYINPUT111), .B(KEYINPUT44), .ZN(n544) );
  XNOR2_X1 U606 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U607 ( .A(G106GAT), .B(n546), .ZN(G1339GAT) );
  XOR2_X1 U608 ( .A(G120GAT), .B(KEYINPUT49), .Z(n548) );
  NAND2_X1 U609 ( .A1(n551), .A2(n558), .ZN(n547) );
  XNOR2_X1 U610 ( .A(n548), .B(n547), .ZN(G1341GAT) );
  NAND2_X1 U611 ( .A1(n551), .A2(n583), .ZN(n549) );
  XNOR2_X1 U612 ( .A(n549), .B(KEYINPUT50), .ZN(n550) );
  XNOR2_X1 U613 ( .A(G127GAT), .B(n550), .ZN(G1342GAT) );
  XOR2_X1 U614 ( .A(G134GAT), .B(KEYINPUT51), .Z(n553) );
  NAND2_X1 U615 ( .A1(n551), .A2(n568), .ZN(n552) );
  XNOR2_X1 U616 ( .A(n553), .B(n552), .ZN(G1343GAT) );
  NOR2_X1 U617 ( .A1(n554), .A2(n555), .ZN(n556) );
  XOR2_X1 U618 ( .A(KEYINPUT119), .B(n556), .Z(n564) );
  NAND2_X1 U619 ( .A1(n575), .A2(n564), .ZN(n557) );
  XNOR2_X1 U620 ( .A(n557), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n560) );
  NAND2_X1 U622 ( .A1(n564), .A2(n558), .ZN(n559) );
  XNOR2_X1 U623 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U624 ( .A(G148GAT), .B(n561), .ZN(G1345GAT) );
  NAND2_X1 U625 ( .A1(n564), .A2(n583), .ZN(n562) );
  XNOR2_X1 U626 ( .A(n562), .B(KEYINPUT120), .ZN(n563) );
  XNOR2_X1 U627 ( .A(G155GAT), .B(n563), .ZN(G1346GAT) );
  NAND2_X1 U628 ( .A1(n564), .A2(n568), .ZN(n565) );
  XNOR2_X1 U629 ( .A(n565), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U630 ( .A1(n575), .A2(n569), .ZN(n566) );
  XNOR2_X1 U631 ( .A(n566), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U632 ( .A1(n569), .A2(n583), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n567), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n571) );
  XOR2_X1 U635 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U637 ( .A(G190GAT), .B(n572), .ZN(G1351GAT) );
  INV_X1 U638 ( .A(n573), .ZN(n574) );
  NOR2_X1 U639 ( .A1(n574), .A2(n554), .ZN(n588) );
  AND2_X1 U640 ( .A1(n575), .A2(n588), .ZN(n577) );
  XNOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(n578), .ZN(G1352GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n581) );
  NAND2_X1 U645 ( .A1(n588), .A2(n579), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(G204GAT), .B(n582), .ZN(G1353GAT) );
  XOR2_X1 U648 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n585) );
  NAND2_X1 U649 ( .A1(n588), .A2(n583), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(G211GAT), .B(n586), .ZN(G1354GAT) );
  XOR2_X1 U652 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n590) );
  NAND2_X1 U653 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

