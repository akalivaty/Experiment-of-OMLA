//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 1 0 0 0 1 1 1 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 1 1 0 0 0 0 0 1 0 1 0 0 1 1 0 1 1 0 0 0 0 0 0 0 0 1 0 0 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n762, new_n764, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n865, new_n866, new_n867, new_n868, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n991, new_n992, new_n993, new_n994,
    new_n996, new_n997, new_n998;
  XNOR2_X1  g000(.A(KEYINPUT92), .B(KEYINPUT15), .ZN(new_n202));
  INV_X1    g001(.A(G43gat), .ZN(new_n203));
  AOI21_X1  g002(.A(KEYINPUT93), .B1(new_n203), .B2(G50gat), .ZN(new_n204));
  INV_X1    g003(.A(G50gat), .ZN(new_n205));
  AOI21_X1  g004(.A(new_n204), .B1(G43gat), .B2(new_n205), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n203), .A2(KEYINPUT93), .A3(G50gat), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n202), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  OR3_X1    g007(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n205), .A2(G43gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n203), .A2(G50gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n212), .A2(new_n213), .A3(KEYINPUT15), .ZN(new_n214));
  INV_X1    g013(.A(G29gat), .ZN(new_n215));
  INV_X1    g014(.A(G36gat), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n211), .B(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n208), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n210), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT91), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n219), .B1(new_n209), .B2(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(new_n220), .B2(new_n209), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n222), .B1(new_n215), .B2(new_n216), .ZN(new_n223));
  INV_X1    g022(.A(new_n214), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n218), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  OR2_X1    g024(.A1(new_n225), .A2(KEYINPUT17), .ZN(new_n226));
  XNOR2_X1  g025(.A(G15gat), .B(G22gat), .ZN(new_n227));
  OR2_X1    g026(.A1(new_n227), .A2(G1gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT16), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n227), .B1(new_n229), .B2(G1gat), .ZN(new_n230));
  INV_X1    g029(.A(G8gat), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n228), .B(new_n230), .C1(KEYINPUT94), .C2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n228), .A2(KEYINPUT94), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n228), .A2(new_n230), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(new_n234), .A3(G8gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n225), .A2(KEYINPUT17), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n226), .A2(new_n232), .A3(new_n235), .A4(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(G229gat), .A2(G233gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n235), .A2(new_n232), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT95), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n239), .B(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n225), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n237), .A2(new_n238), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT18), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n237), .A2(new_n243), .A3(KEYINPUT18), .A4(new_n238), .ZN(new_n247));
  XOR2_X1   g046(.A(new_n238), .B(KEYINPUT13), .Z(new_n248));
  INV_X1    g047(.A(new_n243), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n241), .A2(new_n242), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n246), .A2(new_n247), .A3(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(G113gat), .B(G141gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(G197gat), .ZN(new_n254));
  XOR2_X1   g053(.A(KEYINPUT11), .B(G169gat), .Z(new_n255));
  XNOR2_X1  g054(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XOR2_X1   g055(.A(new_n256), .B(KEYINPUT12), .Z(new_n257));
  NAND2_X1  g056(.A1(new_n252), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n257), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n246), .A2(new_n251), .A3(new_n259), .A4(new_n247), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT22), .ZN(new_n263));
  AOI22_X1  g062(.A1(new_n263), .A2(KEYINPUT72), .B1(G211gat), .B2(G218gat), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n264), .B1(KEYINPUT72), .B2(new_n263), .ZN(new_n265));
  XNOR2_X1  g064(.A(G197gat), .B(G204gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  XOR2_X1   g066(.A(G211gat), .B(G218gat), .Z(new_n268));
  OR3_X1    g067(.A1(new_n267), .A2(KEYINPUT74), .A3(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(KEYINPUT74), .B1(new_n267), .B2(new_n268), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n268), .ZN(new_n272));
  INV_X1    g071(.A(new_n267), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT73), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n267), .A2(KEYINPUT73), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AND2_X1   g076(.A1(new_n271), .A2(new_n277), .ZN(new_n278));
  NOR2_X1   g077(.A1(G155gat), .A2(G162gat), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n279), .A2(KEYINPUT76), .ZN(new_n280));
  XNOR2_X1  g079(.A(G155gat), .B(G162gat), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n280), .B1(new_n281), .B2(KEYINPUT76), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT2), .ZN(new_n283));
  XNOR2_X1  g082(.A(G141gat), .B(G148gat), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n283), .B1(new_n284), .B2(KEYINPUT77), .ZN(new_n285));
  INV_X1    g084(.A(G148gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(G141gat), .ZN(new_n287));
  INV_X1    g086(.A(G141gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(G148gat), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n287), .A2(new_n289), .A3(KEYINPUT77), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n282), .B1(new_n285), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT3), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n288), .A2(KEYINPUT78), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT78), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(G141gat), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n294), .A2(new_n296), .A3(G148gat), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT79), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n298), .B1(new_n288), .B2(G148gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n286), .A2(KEYINPUT79), .A3(G141gat), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n297), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n279), .A2(new_n283), .ZN(new_n302));
  AND2_X1   g101(.A1(G155gat), .A2(G162gat), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n292), .A2(new_n293), .A3(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT29), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n278), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(G228gat), .A2(G233gat), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n277), .A2(new_n271), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT3), .B1(new_n313), .B2(new_n308), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT77), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n288), .A2(G148gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n286), .A2(G141gat), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n318), .A2(new_n283), .A3(new_n290), .ZN(new_n319));
  AOI22_X1  g118(.A1(new_n319), .A2(new_n282), .B1(new_n301), .B2(new_n305), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n310), .B(new_n312), .C1(new_n314), .C2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(G22gat), .ZN(new_n322));
  AOI22_X1  g121(.A1(new_n269), .A2(new_n270), .B1(new_n268), .B2(new_n267), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n293), .B1(new_n323), .B2(KEYINPUT29), .ZN(new_n324));
  INV_X1    g123(.A(new_n320), .ZN(new_n325));
  AOI22_X1  g124(.A1(new_n324), .A2(new_n325), .B1(new_n278), .B2(new_n309), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n321), .B(new_n322), .C1(new_n312), .C2(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G78gat), .B(G106gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(KEYINPUT31), .B(G50gat), .ZN(new_n329));
  XOR2_X1   g128(.A(new_n328), .B(new_n329), .Z(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n324), .A2(new_n325), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(new_n310), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(new_n311), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n322), .B1(new_n335), .B2(new_n321), .ZN(new_n336));
  OAI21_X1  g135(.A(KEYINPUT85), .B1(new_n332), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n321), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n326), .A2(new_n312), .ZN(new_n339));
  OAI21_X1  g138(.A(G22gat), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT85), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n340), .A2(new_n341), .A3(new_n331), .A4(new_n327), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n337), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT84), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n327), .A2(new_n344), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n335), .A2(KEYINPUT84), .A3(new_n322), .A4(new_n321), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(new_n340), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(new_n330), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT83), .ZN(new_n350));
  XOR2_X1   g149(.A(G1gat), .B(G29gat), .Z(new_n351));
  XNOR2_X1  g150(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n351), .B(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(G57gat), .B(G85gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n353), .B(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT76), .B1(new_n303), .B2(new_n279), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT76), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n358), .B1(G155gat), .B2(G162gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n287), .A2(new_n289), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT2), .B1(new_n361), .B2(new_n315), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n360), .B1(new_n362), .B2(new_n290), .ZN(new_n363));
  AND2_X1   g162(.A1(new_n299), .A2(new_n300), .ZN(new_n364));
  AOI22_X1  g163(.A1(new_n364), .A2(new_n297), .B1(new_n304), .B2(new_n302), .ZN(new_n365));
  OAI21_X1  g164(.A(KEYINPUT3), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(G134gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(G127gat), .ZN(new_n368));
  OR2_X1    g167(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n369));
  INV_X1    g168(.A(G127gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(G134gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n372));
  AND4_X1   g171(.A1(new_n368), .A2(new_n369), .A3(new_n371), .A4(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(G113gat), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT67), .B1(new_n374), .B2(G120gat), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT68), .ZN(new_n376));
  INV_X1    g175(.A(G120gat), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n376), .B1(new_n377), .B2(G113gat), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT67), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n379), .A2(new_n377), .A3(G113gat), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n374), .A2(KEYINPUT68), .A3(G120gat), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n375), .A2(new_n378), .A3(new_n380), .A4(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n373), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n377), .A2(G113gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n374), .A2(G120gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT1), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n370), .A2(G134gat), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n367), .A2(G127gat), .ZN(new_n390));
  OAI21_X1  g189(.A(KEYINPUT66), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT66), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n368), .A2(new_n371), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n388), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n383), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n366), .A2(new_n307), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(G225gat), .A2(G233gat), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n292), .A2(new_n306), .A3(new_n383), .A4(new_n394), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT4), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT1), .B1(new_n384), .B2(new_n385), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n392), .B1(new_n368), .B2(new_n371), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI22_X1  g202(.A1(new_n403), .A2(new_n393), .B1(new_n382), .B2(new_n373), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n320), .A2(new_n404), .A3(KEYINPUT4), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n396), .A2(new_n397), .A3(new_n400), .A4(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT5), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n395), .B1(new_n363), .B2(new_n365), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n398), .ZN(new_n409));
  INV_X1    g208(.A(new_n397), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n407), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  AND2_X1   g210(.A1(new_n406), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n406), .A2(KEYINPUT5), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n356), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT6), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT81), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n406), .A2(new_n411), .ZN(new_n418));
  AND3_X1   g217(.A1(new_n320), .A2(new_n404), .A3(KEYINPUT4), .ZN(new_n419));
  AOI21_X1  g218(.A(KEYINPUT4), .B1(new_n320), .B2(new_n404), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n421), .A2(new_n407), .A3(new_n397), .A4(new_n396), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n418), .A2(new_n422), .A3(new_n355), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n417), .B1(new_n423), .B2(new_n415), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT82), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n418), .A2(new_n422), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n425), .B1(new_n426), .B2(new_n356), .ZN(new_n427));
  AOI211_X1 g226(.A(KEYINPUT82), .B(new_n355), .C1(new_n418), .C2(new_n422), .ZN(new_n428));
  NOR3_X1   g227(.A1(new_n424), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n423), .A2(new_n417), .A3(new_n415), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n416), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT75), .ZN(new_n432));
  NAND2_X1  g231(.A1(G226gat), .A2(G233gat), .ZN(new_n433));
  NOR2_X1   g232(.A1(G169gat), .A2(G176gat), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT26), .ZN(new_n436));
  NAND2_X1  g235(.A1(G169gat), .A2(G176gat), .ZN(new_n437));
  AND3_X1   g236(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(G183gat), .A2(G190gat), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n439), .B1(new_n435), .B2(new_n436), .ZN(new_n440));
  XNOR2_X1  g239(.A(KEYINPUT27), .B(G183gat), .ZN(new_n441));
  INV_X1    g240(.A(G190gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT28), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n441), .A2(KEYINPUT28), .A3(new_n442), .ZN(new_n446));
  AOI211_X1 g245(.A(new_n438), .B(new_n440), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(G169gat), .ZN(new_n448));
  INV_X1    g247(.A(G176gat), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(new_n449), .A3(KEYINPUT23), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT24), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n451), .A2(G183gat), .A3(G190gat), .ZN(new_n452));
  AND3_X1   g251(.A1(new_n450), .A2(new_n452), .A3(new_n437), .ZN(new_n453));
  OAI21_X1  g252(.A(KEYINPUT64), .B1(new_n434), .B2(KEYINPUT23), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT64), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT23), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n455), .B(new_n456), .C1(G169gat), .C2(G176gat), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  OR2_X1    g257(.A1(G183gat), .A2(G190gat), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n459), .A2(KEYINPUT24), .A3(new_n439), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n453), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT65), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT25), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n462), .A2(KEYINPUT25), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT25), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n461), .A2(KEYINPUT65), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n447), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n433), .B1(new_n470), .B2(KEYINPUT29), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n445), .A2(new_n446), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n438), .A2(new_n440), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n461), .A2(KEYINPUT65), .A3(new_n468), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n465), .B1(new_n461), .B2(new_n463), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n433), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n432), .B1(new_n471), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n478), .B1(new_n477), .B2(new_n308), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n481), .A2(KEYINPUT75), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n278), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n469), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n433), .B1(new_n484), .B2(new_n474), .ZN(new_n485));
  NOR3_X1   g284(.A1(new_n481), .A2(new_n485), .A3(new_n278), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  XNOR2_X1  g286(.A(G8gat), .B(G36gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(G64gat), .B(G92gat), .ZN(new_n489));
  XOR2_X1   g288(.A(new_n488), .B(new_n489), .Z(new_n490));
  NAND3_X1  g289(.A1(new_n483), .A2(new_n487), .A3(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT30), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n490), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT75), .B1(new_n481), .B2(new_n485), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n471), .A2(new_n432), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n313), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n494), .B1(new_n497), .B2(new_n486), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n483), .A2(KEYINPUT30), .A3(new_n487), .A4(new_n490), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n493), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n350), .B1(new_n431), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n499), .A2(new_n498), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n495), .A2(new_n496), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n486), .B1(new_n503), .B2(new_n278), .ZN(new_n504));
  AOI21_X1  g303(.A(KEYINPUT30), .B1(new_n504), .B2(new_n490), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n423), .A2(new_n415), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT81), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n414), .A2(KEYINPUT82), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n426), .A2(new_n425), .A3(new_n356), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n508), .A2(new_n430), .A3(new_n509), .A4(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n416), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n506), .A2(new_n513), .A3(KEYINPUT83), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n349), .B1(new_n501), .B2(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(G15gat), .B(G43gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(KEYINPUT70), .ZN(new_n517));
  XNOR2_X1  g316(.A(G71gat), .B(G99gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n517), .B(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n470), .A2(new_n395), .ZN(new_n520));
  INV_X1    g319(.A(G227gat), .ZN(new_n521));
  INV_X1    g320(.A(G233gat), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n477), .A2(new_n404), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n520), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT33), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n519), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n525), .A2(KEYINPUT32), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n525), .B(KEYINPUT32), .C1(new_n526), .C2(new_n519), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n523), .B1(new_n520), .B2(new_n524), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT34), .ZN(new_n533));
  OR2_X1    g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n533), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n531), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n532), .B(KEYINPUT34), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n538), .A2(new_n529), .A3(new_n530), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT36), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT71), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g343(.A(KEYINPUT71), .B1(new_n531), .B2(new_n536), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n542), .B1(new_n546), .B2(new_n541), .ZN(new_n547));
  OAI21_X1  g346(.A(KEYINPUT86), .B1(new_n515), .B2(new_n547), .ZN(new_n548));
  AOI22_X1  g347(.A1(new_n337), .A2(new_n342), .B1(new_n347), .B2(new_n330), .ZN(new_n549));
  AND3_X1   g348(.A1(new_n506), .A2(new_n513), .A3(KEYINPUT83), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT83), .B1(new_n506), .B2(new_n513), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT86), .ZN(new_n553));
  INV_X1    g352(.A(new_n542), .ZN(new_n554));
  INV_X1    g353(.A(new_n545), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n555), .B1(new_n540), .B2(new_n543), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n554), .B1(new_n556), .B2(KEYINPUT36), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n552), .A2(new_n553), .A3(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT87), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n500), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n396), .A2(new_n400), .A3(new_n405), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(new_n410), .ZN(new_n562));
  OR2_X1    g361(.A1(new_n562), .A2(KEYINPUT39), .ZN(new_n563));
  OAI211_X1 g362(.A(new_n562), .B(KEYINPUT39), .C1(new_n410), .C2(new_n409), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n563), .A2(new_n564), .A3(new_n355), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT40), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(new_n414), .ZN(new_n568));
  OR3_X1    g367(.A1(new_n565), .A2(KEYINPUT88), .A3(new_n566), .ZN(new_n569));
  OAI21_X1  g368(.A(KEYINPUT88), .B1(new_n565), .B2(new_n566), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n493), .A2(KEYINPUT87), .A3(new_n498), .A4(new_n499), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n560), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT89), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n483), .A2(new_n487), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n494), .B1(new_n576), .B2(KEYINPUT37), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT38), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n278), .B1(new_n495), .B2(new_n496), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n471), .A2(new_n479), .A3(new_n278), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(KEYINPUT37), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n578), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n577), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n414), .A2(new_n415), .A3(new_n423), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n512), .A2(new_n491), .A3(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  AND2_X1   g385(.A1(new_n576), .A2(KEYINPUT37), .ZN(new_n587));
  OAI21_X1  g386(.A(KEYINPUT38), .B1(new_n587), .B2(new_n577), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n549), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n560), .A2(new_n571), .A3(KEYINPUT89), .A4(new_n572), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n575), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n548), .A2(new_n558), .A3(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n549), .A2(new_n540), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n501), .A2(new_n514), .ZN(new_n595));
  OAI21_X1  g394(.A(KEYINPUT35), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n560), .A2(new_n572), .ZN(new_n597));
  XOR2_X1   g396(.A(KEYINPUT90), .B(KEYINPUT35), .Z(new_n598));
  AOI21_X1  g397(.A(new_n598), .B1(new_n512), .B2(new_n584), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n597), .A2(new_n556), .A3(new_n349), .A4(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n262), .B1(new_n592), .B2(new_n601), .ZN(new_n602));
  XOR2_X1   g401(.A(G57gat), .B(G64gat), .Z(new_n603));
  INV_X1    g402(.A(KEYINPUT9), .ZN(new_n604));
  INV_X1    g403(.A(G71gat), .ZN(new_n605));
  INV_X1    g404(.A(G78gat), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(G71gat), .B(G78gat), .Z(new_n609));
  OR2_X1    g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n608), .A2(new_n609), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT21), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n241), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT96), .ZN(new_n616));
  XNOR2_X1  g415(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(G155gat), .ZN(new_n618));
  OR2_X1    g417(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n616), .A2(new_n618), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n612), .A2(new_n613), .ZN(new_n622));
  NAND2_X1  g421(.A1(G231gat), .A2(G233gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(new_n370), .ZN(new_n625));
  XNOR2_X1  g424(.A(G183gat), .B(G211gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n621), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n619), .A2(new_n627), .A3(new_n620), .ZN(new_n630));
  AND2_X1   g429(.A1(G232gat), .A2(G233gat), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n631), .A2(KEYINPUT41), .ZN(new_n632));
  XNOR2_X1  g431(.A(G134gat), .B(G162gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(G85gat), .A2(G92gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT7), .ZN(new_n637));
  NAND2_X1  g436(.A1(G99gat), .A2(G106gat), .ZN(new_n638));
  INV_X1    g437(.A(G85gat), .ZN(new_n639));
  INV_X1    g438(.A(G92gat), .ZN(new_n640));
  AOI22_X1  g439(.A1(KEYINPUT8), .A2(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(G99gat), .B(G106gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n226), .A2(new_n236), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g445(.A(G190gat), .B(G218gat), .Z(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  AOI22_X1  g447(.A1(new_n242), .A2(new_n644), .B1(KEYINPUT41), .B2(new_n631), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n646), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n648), .B1(new_n646), .B2(new_n649), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n635), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n652), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n654), .A2(new_n634), .A3(new_n650), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n629), .A2(new_n630), .A3(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT97), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND4_X1  g458(.A1(new_n629), .A2(KEYINPUT97), .A3(new_n630), .A4(new_n656), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n644), .B(new_n612), .ZN(new_n661));
  NAND2_X1  g460(.A1(G230gat), .A2(G233gat), .ZN(new_n662));
  OR3_X1    g461(.A1(new_n661), .A2(KEYINPUT98), .A3(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(KEYINPUT98), .B1(new_n661), .B2(new_n662), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(G120gat), .B(G148gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(G176gat), .B(G204gat), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n667), .B(new_n668), .Z(new_n669));
  INV_X1    g468(.A(KEYINPUT10), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n661), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n644), .A2(KEYINPUT10), .A3(new_n611), .A4(new_n610), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(new_n662), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n666), .A2(new_n669), .A3(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n669), .ZN(new_n676));
  INV_X1    g475(.A(new_n662), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n677), .B1(new_n671), .B2(new_n672), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n676), .B1(new_n665), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT99), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n675), .A2(KEYINPUT99), .A3(new_n679), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n659), .A2(new_n660), .A3(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n513), .B(KEYINPUT100), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n602), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g488(.A1(new_n685), .A2(new_n597), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n602), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  XOR2_X1   g491(.A(KEYINPUT16), .B(G8gat), .Z(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n694), .B1(new_n692), .B2(new_n231), .ZN(new_n695));
  MUX2_X1   g494(.A(new_n694), .B(new_n695), .S(KEYINPUT42), .Z(G1325gat));
  NAND2_X1  g495(.A1(new_n602), .A2(new_n686), .ZN(new_n697));
  OAI21_X1  g496(.A(G15gat), .B1(new_n697), .B2(new_n557), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n546), .A2(G15gat), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n698), .B1(new_n697), .B2(new_n699), .ZN(G1326gat));
  NOR2_X1   g499(.A1(new_n697), .A2(new_n349), .ZN(new_n701));
  XOR2_X1   g500(.A(KEYINPUT43), .B(G22gat), .Z(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(G1327gat));
  AOI21_X1  g502(.A(new_n656), .B1(new_n592), .B2(new_n601), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n629), .A2(new_n630), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n684), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n706), .A2(new_n262), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n704), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n710), .A2(new_n215), .A3(new_n687), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT45), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n592), .A2(new_n601), .ZN(new_n714));
  INV_X1    g513(.A(new_n656), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n515), .A2(new_n547), .ZN(new_n717));
  AOI22_X1  g516(.A1(new_n596), .A2(new_n600), .B1(new_n717), .B2(new_n591), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT102), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n656), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n653), .A2(new_n655), .A3(KEYINPUT102), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n718), .A2(KEYINPUT44), .A3(new_n723), .ZN(new_n724));
  OR2_X1    g523(.A1(new_n716), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n708), .B(KEYINPUT101), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n687), .ZN(new_n728));
  OAI21_X1  g527(.A(G29gat), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n712), .A2(new_n729), .ZN(G1328gat));
  NOR3_X1   g529(.A1(new_n709), .A2(G36gat), .A3(new_n597), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT46), .ZN(new_n732));
  OAI21_X1  g531(.A(G36gat), .B1(new_n727), .B2(new_n597), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(G1329gat));
  OAI211_X1 g533(.A(new_n547), .B(new_n726), .C1(new_n716), .C2(new_n724), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(G43gat), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n710), .A2(new_n203), .A3(new_n556), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT47), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n738), .B(new_n739), .ZN(G1330gat));
  OAI211_X1 g539(.A(new_n549), .B(new_n726), .C1(new_n716), .C2(new_n724), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(G50gat), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n710), .A2(new_n205), .A3(new_n549), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT48), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n744), .B(new_n745), .ZN(G1331gat));
  NAND2_X1  g545(.A1(new_n717), .A2(new_n591), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n601), .A2(new_n747), .ZN(new_n748));
  AND4_X1   g547(.A1(new_n262), .A2(new_n659), .A3(new_n660), .A4(new_n707), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(new_n687), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(G57gat), .ZN(G1332gat));
  INV_X1    g551(.A(new_n597), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n755));
  XOR2_X1   g554(.A(KEYINPUT49), .B(G64gat), .Z(new_n756));
  OAI21_X1  g555(.A(new_n755), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  XOR2_X1   g556(.A(new_n757), .B(KEYINPUT103), .Z(G1333gat));
  INV_X1    g557(.A(new_n750), .ZN(new_n759));
  OAI21_X1  g558(.A(G71gat), .B1(new_n759), .B2(new_n557), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n750), .A2(new_n605), .A3(new_n556), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  XOR2_X1   g561(.A(new_n762), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g562(.A1(new_n750), .A2(new_n549), .ZN(new_n764));
  XNOR2_X1  g563(.A(KEYINPUT104), .B(G78gat), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n764), .B(new_n765), .ZN(G1335gat));
  NOR3_X1   g565(.A1(new_n706), .A2(new_n261), .A3(new_n684), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n725), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(G85gat), .B1(new_n768), .B2(new_n728), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n706), .A2(new_n261), .ZN(new_n770));
  NOR2_X1   g569(.A1(KEYINPUT105), .A2(KEYINPUT51), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n656), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  OAI211_X1 g572(.A(KEYINPUT105), .B(KEYINPUT51), .C1(new_n718), .C2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(KEYINPUT105), .A2(KEYINPUT51), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n748), .A2(new_n770), .A3(new_n775), .A4(new_n772), .ZN(new_n776));
  AND2_X1   g575(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n687), .A2(new_n639), .A3(new_n707), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(KEYINPUT106), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n769), .A2(new_n780), .ZN(G1336gat));
  NAND3_X1  g580(.A1(new_n725), .A2(new_n753), .A3(new_n767), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(G92gat), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n597), .A2(G92gat), .A3(new_n684), .ZN(new_n784));
  AOI21_X1  g583(.A(KEYINPUT52), .B1(new_n777), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n784), .B(KEYINPUT107), .ZN(new_n787));
  AOI22_X1  g586(.A1(new_n782), .A2(G92gat), .B1(new_n777), .B2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n786), .B1(new_n788), .B2(new_n789), .ZN(G1337gat));
  OAI21_X1  g589(.A(G99gat), .B1(new_n768), .B2(new_n557), .ZN(new_n791));
  INV_X1    g590(.A(G99gat), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n546), .A2(new_n684), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n777), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n791), .A2(new_n794), .ZN(G1338gat));
  INV_X1    g594(.A(KEYINPUT110), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n549), .B(new_n767), .C1(new_n716), .C2(new_n724), .ZN(new_n798));
  XNOR2_X1  g597(.A(KEYINPUT108), .B(G106gat), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n349), .A2(new_n684), .A3(G106gat), .ZN(new_n801));
  XOR2_X1   g600(.A(new_n801), .B(KEYINPUT109), .Z(new_n802));
  NAND2_X1  g601(.A1(new_n777), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n797), .B1(new_n800), .B2(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n774), .A2(new_n776), .A3(new_n801), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(new_n797), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n806), .B1(new_n798), .B2(new_n799), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n796), .B1(new_n804), .B2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n806), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n800), .ZN(new_n810));
  AOI22_X1  g609(.A1(new_n798), .A2(new_n799), .B1(new_n777), .B2(new_n802), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n810), .B(KEYINPUT110), .C1(new_n811), .C2(new_n797), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n808), .A2(new_n812), .ZN(G1339gat));
  NAND3_X1  g612(.A1(new_n671), .A2(new_n677), .A3(new_n672), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n674), .A2(KEYINPUT54), .A3(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n669), .B1(new_n678), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n815), .A2(KEYINPUT55), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n675), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT111), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n818), .A2(new_n675), .A3(KEYINPUT111), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n815), .A2(new_n817), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT55), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n821), .A2(new_n261), .A3(new_n822), .A4(new_n825), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n249), .A2(new_n250), .A3(new_n248), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n238), .B1(new_n237), .B2(new_n243), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n256), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n260), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n830), .A2(new_n682), .A3(new_n683), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n722), .B1(new_n826), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n821), .A2(new_n822), .A3(new_n825), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n720), .A2(new_n830), .A3(new_n721), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n705), .B1(new_n832), .B2(new_n835), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n659), .A2(new_n262), .A3(new_n660), .A4(new_n684), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(KEYINPUT112), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT112), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n836), .A2(new_n837), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n842), .A2(new_n728), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n594), .A2(new_n753), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n261), .A2(new_n374), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n847), .B(KEYINPUT114), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n842), .A2(new_n549), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n850), .A2(new_n597), .A3(new_n556), .A4(new_n687), .ZN(new_n851));
  OAI21_X1  g650(.A(G113gat), .B1(new_n851), .B2(new_n262), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT113), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  OAI211_X1 g653(.A(KEYINPUT113), .B(G113gat), .C1(new_n851), .C2(new_n262), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n849), .B1(new_n854), .B2(new_n856), .ZN(G1340gat));
  NAND3_X1  g656(.A1(new_n846), .A2(new_n377), .A3(new_n707), .ZN(new_n858));
  OAI21_X1  g657(.A(G120gat), .B1(new_n851), .B2(new_n684), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT115), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI211_X1 g660(.A(KEYINPUT115), .B(G120gat), .C1(new_n851), .C2(new_n684), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n858), .B1(new_n861), .B2(new_n863), .ZN(G1341gat));
  NOR3_X1   g663(.A1(new_n851), .A2(new_n370), .A3(new_n705), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n845), .A2(KEYINPUT116), .A3(new_n705), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n866), .A2(G127gat), .ZN(new_n867));
  OAI21_X1  g666(.A(KEYINPUT116), .B1(new_n845), .B2(new_n705), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n865), .B1(new_n867), .B2(new_n868), .ZN(G1342gat));
  NOR3_X1   g668(.A1(new_n845), .A2(G134gat), .A3(new_n656), .ZN(new_n870));
  XOR2_X1   g669(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n871));
  OR2_X1    g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(G134gat), .B1(new_n851), .B2(new_n656), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n870), .A2(new_n871), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(G1343gat));
  INV_X1    g674(.A(new_n837), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n831), .A2(KEYINPUT118), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT118), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n830), .A2(new_n682), .A3(new_n878), .A4(new_n683), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n261), .A2(new_n675), .A3(new_n818), .A4(new_n825), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n877), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n656), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n882), .B1(new_n833), .B2(new_n834), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n876), .B1(new_n883), .B2(new_n705), .ZN(new_n884));
  OAI21_X1  g683(.A(KEYINPUT57), .B1(new_n884), .B2(new_n349), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT57), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n839), .A2(new_n886), .A3(new_n549), .A4(new_n841), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n728), .A2(new_n547), .A3(new_n753), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n885), .A2(new_n261), .A3(new_n887), .A4(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n294), .A2(new_n296), .ZN(new_n890));
  AOI21_X1  g689(.A(KEYINPUT120), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n547), .A2(new_n349), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n597), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n839), .A2(new_n687), .A3(new_n841), .A4(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n261), .A2(new_n288), .ZN(new_n896));
  XOR2_X1   g695(.A(new_n896), .B(KEYINPUT119), .Z(new_n897));
  NOR2_X1   g696(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n898), .B1(new_n889), .B2(new_n890), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n891), .A2(new_n899), .A3(KEYINPUT58), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT58), .ZN(new_n901));
  AOI221_X4 g700(.A(new_n898), .B1(KEYINPUT120), .B2(new_n901), .C1(new_n889), .C2(new_n890), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n900), .A2(new_n902), .ZN(G1344gat));
  NAND3_X1  g702(.A1(new_n839), .A2(new_n549), .A3(new_n841), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(KEYINPUT57), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT122), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n833), .A2(new_n906), .A3(new_n656), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n906), .B1(new_n833), .B2(new_n656), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n830), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n882), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(new_n705), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(new_n837), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n349), .A2(KEYINPUT57), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT123), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT121), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n888), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n888), .A2(new_n916), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n917), .A2(new_n918), .A3(new_n684), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n905), .A2(new_n914), .A3(new_n915), .A4(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(G148gat), .ZN(new_n921));
  AOI22_X1  g720(.A1(new_n904), .A2(KEYINPUT57), .B1(new_n912), .B2(new_n913), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n915), .B1(new_n922), .B2(new_n919), .ZN(new_n923));
  OAI21_X1  g722(.A(KEYINPUT59), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n286), .A2(KEYINPUT59), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n885), .A2(new_n887), .A3(new_n888), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n925), .B1(new_n926), .B2(new_n684), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(new_n895), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n929), .A2(new_n286), .A3(new_n707), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(G1345gat));
  OAI21_X1  g730(.A(G155gat), .B1(new_n926), .B2(new_n705), .ZN(new_n932));
  OR3_X1    g731(.A1(new_n895), .A2(G155gat), .A3(new_n705), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT124), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n932), .A2(KEYINPUT124), .A3(new_n933), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(G1346gat));
  INV_X1    g737(.A(G162gat), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n926), .A2(new_n939), .A3(new_n723), .ZN(new_n940));
  AOI21_X1  g739(.A(G162gat), .B1(new_n929), .B2(new_n715), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n940), .A2(new_n941), .ZN(G1347gat));
  NOR2_X1   g741(.A1(new_n687), .A2(new_n597), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n850), .A2(new_n943), .ZN(new_n944));
  AND4_X1   g743(.A1(G169gat), .A2(new_n944), .A3(new_n261), .A4(new_n556), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n839), .A2(new_n728), .A3(new_n841), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT125), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n597), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n839), .A2(KEYINPUT125), .A3(new_n728), .A4(new_n841), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n950), .A2(new_n261), .A3(new_n593), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n945), .B1(new_n448), .B2(new_n951), .ZN(G1348gat));
  NAND4_X1  g751(.A1(new_n948), .A2(new_n593), .A3(new_n707), .A4(new_n949), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(new_n449), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n944), .A2(G176gat), .A3(new_n793), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT126), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n954), .A2(new_n955), .A3(KEYINPUT126), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(G1349gat));
  NAND4_X1  g759(.A1(new_n850), .A2(new_n556), .A3(new_n706), .A4(new_n943), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(G183gat), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n706), .A2(new_n441), .ZN(new_n963));
  INV_X1    g762(.A(new_n963), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n948), .A2(new_n593), .A3(new_n949), .A4(new_n964), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n966), .B(KEYINPUT60), .ZN(G1350gat));
  NAND4_X1  g766(.A1(new_n950), .A2(new_n442), .A3(new_n593), .A4(new_n722), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n944), .A2(new_n556), .A3(new_n715), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT61), .ZN(new_n970));
  AND3_X1   g769(.A1(new_n969), .A2(new_n970), .A3(G190gat), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n970), .B1(new_n969), .B2(G190gat), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n968), .B1(new_n971), .B2(new_n972), .ZN(G1351gat));
  NAND3_X1  g772(.A1(new_n950), .A2(new_n261), .A3(new_n892), .ZN(new_n974));
  INV_X1    g773(.A(G197gat), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n943), .A2(new_n557), .ZN(new_n976));
  INV_X1    g775(.A(new_n976), .ZN(new_n977));
  AND2_X1   g776(.A1(new_n922), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n262), .A2(new_n975), .ZN(new_n979));
  AOI22_X1  g778(.A1(new_n974), .A2(new_n975), .B1(new_n978), .B2(new_n979), .ZN(G1352gat));
  XOR2_X1   g779(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n981));
  INV_X1    g780(.A(new_n981), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n950), .A2(new_n892), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n684), .A2(G204gat), .ZN(new_n984));
  INV_X1    g783(.A(new_n984), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n982), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n978), .A2(new_n707), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n987), .A2(G204gat), .ZN(new_n988));
  NAND4_X1  g787(.A1(new_n950), .A2(new_n892), .A3(new_n984), .A4(new_n981), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n986), .A2(new_n988), .A3(new_n989), .ZN(G1353gat));
  NAND3_X1  g789(.A1(new_n922), .A2(new_n706), .A3(new_n977), .ZN(new_n991));
  AND3_X1   g790(.A1(new_n991), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n992));
  AOI21_X1  g791(.A(KEYINPUT63), .B1(new_n991), .B2(G211gat), .ZN(new_n993));
  OR2_X1    g792(.A1(new_n705), .A2(G211gat), .ZN(new_n994));
  OAI22_X1  g793(.A1(new_n992), .A2(new_n993), .B1(new_n983), .B2(new_n994), .ZN(G1354gat));
  NAND2_X1  g794(.A1(new_n978), .A2(new_n715), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n996), .A2(G218gat), .ZN(new_n997));
  OR2_X1    g796(.A1(new_n723), .A2(G218gat), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n997), .B1(new_n983), .B2(new_n998), .ZN(G1355gat));
endmodule


