

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589;

  XNOR2_X1 U322 ( .A(KEYINPUT117), .B(KEYINPUT45), .ZN(n464) );
  XNOR2_X1 U323 ( .A(n465), .B(n464), .ZN(n466) );
  INV_X1 U324 ( .A(KEYINPUT109), .ZN(n433) );
  NOR2_X1 U325 ( .A1(n494), .A2(n527), .ZN(n454) );
  NOR2_X1 U326 ( .A1(n480), .A2(n479), .ZN(n568) );
  XOR2_X1 U327 ( .A(KEYINPUT82), .B(n565), .Z(n549) );
  XNOR2_X1 U328 ( .A(n422), .B(n421), .ZN(n573) );
  XOR2_X1 U329 ( .A(n360), .B(n359), .Z(n529) );
  XNOR2_X1 U330 ( .A(n484), .B(G190GAT), .ZN(n485) );
  XNOR2_X1 U331 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U332 ( .A(n486), .B(n485), .ZN(G1351GAT) );
  XNOR2_X1 U333 ( .A(n458), .B(n457), .ZN(G1330GAT) );
  INV_X1 U334 ( .A(KEYINPUT8), .ZN(n293) );
  XOR2_X1 U335 ( .A(KEYINPUT7), .B(G50GAT), .Z(n291) );
  XNOR2_X1 U336 ( .A(G43GAT), .B(G29GAT), .ZN(n290) );
  XNOR2_X1 U337 ( .A(n291), .B(n290), .ZN(n292) );
  XNOR2_X1 U338 ( .A(n293), .B(n292), .ZN(n435) );
  XOR2_X1 U339 ( .A(G169GAT), .B(G8GAT), .Z(n343) );
  XOR2_X1 U340 ( .A(G15GAT), .B(G1GAT), .Z(n335) );
  XOR2_X1 U341 ( .A(n343), .B(n335), .Z(n295) );
  NAND2_X1 U342 ( .A1(G229GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U343 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U344 ( .A(G141GAT), .B(G22GAT), .Z(n375) );
  XOR2_X1 U345 ( .A(n296), .B(n375), .Z(n304) );
  XOR2_X1 U346 ( .A(KEYINPUT30), .B(G113GAT), .Z(n298) );
  XNOR2_X1 U347 ( .A(G36GAT), .B(G197GAT), .ZN(n297) );
  XNOR2_X1 U348 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U349 ( .A(KEYINPUT70), .B(KEYINPUT29), .Z(n300) );
  XNOR2_X1 U350 ( .A(KEYINPUT69), .B(KEYINPUT68), .ZN(n299) );
  XNOR2_X1 U351 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U352 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U353 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U354 ( .A(n435), .B(n305), .ZN(n576) );
  XNOR2_X1 U355 ( .A(KEYINPUT71), .B(n576), .ZN(n567) );
  XOR2_X1 U356 ( .A(KEYINPUT72), .B(G92GAT), .Z(n307) );
  XOR2_X1 U357 ( .A(G148GAT), .B(G78GAT), .Z(n365) );
  XOR2_X1 U358 ( .A(G57GAT), .B(KEYINPUT13), .Z(n334) );
  XNOR2_X1 U359 ( .A(n365), .B(n334), .ZN(n306) );
  XNOR2_X1 U360 ( .A(n307), .B(n306), .ZN(n313) );
  XOR2_X1 U361 ( .A(G64GAT), .B(KEYINPUT76), .Z(n309) );
  XNOR2_X1 U362 ( .A(G176GAT), .B(G204GAT), .ZN(n308) );
  XNOR2_X1 U363 ( .A(n309), .B(n308), .ZN(n352) );
  XOR2_X1 U364 ( .A(KEYINPUT31), .B(n352), .Z(n311) );
  NAND2_X1 U365 ( .A1(G230GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U366 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U367 ( .A(n313), .B(n312), .Z(n318) );
  XOR2_X1 U368 ( .A(G120GAT), .B(G71GAT), .Z(n388) );
  XOR2_X1 U369 ( .A(KEYINPUT75), .B(KEYINPUT32), .Z(n315) );
  XNOR2_X1 U370 ( .A(KEYINPUT33), .B(KEYINPUT77), .ZN(n314) );
  XNOR2_X1 U371 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U372 ( .A(n388), .B(n316), .ZN(n317) );
  XNOR2_X1 U373 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U374 ( .A(KEYINPUT74), .B(KEYINPUT73), .Z(n320) );
  XNOR2_X1 U375 ( .A(G106GAT), .B(G85GAT), .ZN(n319) );
  XNOR2_X1 U376 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U377 ( .A(G99GAT), .B(n321), .ZN(n450) );
  XOR2_X1 U378 ( .A(n322), .B(n450), .Z(n579) );
  NAND2_X1 U379 ( .A1(n567), .A2(n579), .ZN(n494) );
  XOR2_X1 U380 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n324) );
  NAND2_X1 U381 ( .A1(G231GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U382 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U383 ( .A(G183GAT), .B(KEYINPUT83), .Z(n342) );
  XOR2_X1 U384 ( .A(n325), .B(n342), .Z(n333) );
  XOR2_X1 U385 ( .A(G64GAT), .B(G71GAT), .Z(n327) );
  XNOR2_X1 U386 ( .A(G8GAT), .B(G127GAT), .ZN(n326) );
  XNOR2_X1 U387 ( .A(n327), .B(n326), .ZN(n331) );
  XOR2_X1 U388 ( .A(KEYINPUT86), .B(KEYINPUT84), .Z(n329) );
  XNOR2_X1 U389 ( .A(KEYINPUT85), .B(KEYINPUT15), .ZN(n328) );
  XNOR2_X1 U390 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U391 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U392 ( .A(n333), .B(n332), .ZN(n339) );
  XOR2_X1 U393 ( .A(n334), .B(G211GAT), .Z(n337) );
  XNOR2_X1 U394 ( .A(n335), .B(G155GAT), .ZN(n336) );
  XNOR2_X1 U395 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U396 ( .A(n339), .B(n338), .Z(n341) );
  XNOR2_X1 U397 ( .A(G22GAT), .B(G78GAT), .ZN(n340) );
  XNOR2_X1 U398 ( .A(n341), .B(n340), .ZN(n545) );
  XNOR2_X1 U399 ( .A(n343), .B(n342), .ZN(n360) );
  INV_X1 U400 ( .A(G218GAT), .ZN(n344) );
  NAND2_X1 U401 ( .A1(G92GAT), .A2(n344), .ZN(n347) );
  INV_X1 U402 ( .A(G92GAT), .ZN(n345) );
  NAND2_X1 U403 ( .A1(n345), .A2(G218GAT), .ZN(n346) );
  NAND2_X1 U404 ( .A1(n347), .A2(n346), .ZN(n349) );
  XNOR2_X1 U405 ( .A(G36GAT), .B(G190GAT), .ZN(n348) );
  XNOR2_X1 U406 ( .A(n349), .B(n348), .ZN(n443) );
  XOR2_X1 U407 ( .A(KEYINPUT101), .B(n443), .Z(n351) );
  NAND2_X1 U408 ( .A1(G226GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U409 ( .A(n351), .B(n350), .ZN(n353) );
  XOR2_X1 U410 ( .A(n353), .B(n352), .Z(n358) );
  XOR2_X1 U411 ( .A(KEYINPUT19), .B(KEYINPUT90), .Z(n355) );
  XNOR2_X1 U412 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n354) );
  XNOR2_X1 U413 ( .A(n355), .B(n354), .ZN(n397) );
  XNOR2_X1 U414 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n356) );
  XNOR2_X1 U415 ( .A(n356), .B(G211GAT), .ZN(n376) );
  XNOR2_X1 U416 ( .A(n397), .B(n376), .ZN(n357) );
  XNOR2_X1 U417 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U418 ( .A(n529), .B(KEYINPUT27), .Z(n361) );
  XNOR2_X1 U419 ( .A(n361), .B(KEYINPUT102), .ZN(n428) );
  XOR2_X1 U420 ( .A(KEYINPUT23), .B(KEYINPUT95), .Z(n363) );
  XNOR2_X1 U421 ( .A(G218GAT), .B(G162GAT), .ZN(n362) );
  XNOR2_X1 U422 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U423 ( .A(n364), .B(G106GAT), .Z(n367) );
  XNOR2_X1 U424 ( .A(G50GAT), .B(n365), .ZN(n366) );
  XNOR2_X1 U425 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U426 ( .A(n368), .B(G204GAT), .Z(n372) );
  XOR2_X1 U427 ( .A(G155GAT), .B(KEYINPUT3), .Z(n370) );
  XNOR2_X1 U428 ( .A(KEYINPUT93), .B(KEYINPUT2), .ZN(n369) );
  XNOR2_X1 U429 ( .A(n370), .B(n369), .ZN(n418) );
  XNOR2_X1 U430 ( .A(n418), .B(KEYINPUT96), .ZN(n371) );
  XNOR2_X1 U431 ( .A(n372), .B(n371), .ZN(n382) );
  XOR2_X1 U432 ( .A(KEYINPUT22), .B(KEYINPUT92), .Z(n374) );
  XNOR2_X1 U433 ( .A(KEYINPUT24), .B(KEYINPUT94), .ZN(n373) );
  XNOR2_X1 U434 ( .A(n374), .B(n373), .ZN(n380) );
  XOR2_X1 U435 ( .A(n376), .B(n375), .Z(n378) );
  NAND2_X1 U436 ( .A1(G228GAT), .A2(G233GAT), .ZN(n377) );
  XNOR2_X1 U437 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U438 ( .A(n380), .B(n379), .Z(n381) );
  XNOR2_X1 U439 ( .A(n382), .B(n381), .ZN(n474) );
  XOR2_X1 U440 ( .A(KEYINPUT28), .B(n474), .Z(n532) );
  NOR2_X1 U441 ( .A1(n428), .A2(n532), .ZN(n539) );
  XOR2_X1 U442 ( .A(KEYINPUT89), .B(KEYINPUT20), .Z(n384) );
  XNOR2_X1 U443 ( .A(KEYINPUT91), .B(KEYINPUT87), .ZN(n383) );
  XNOR2_X1 U444 ( .A(n384), .B(n383), .ZN(n392) );
  XOR2_X1 U445 ( .A(KEYINPUT88), .B(G99GAT), .Z(n386) );
  XNOR2_X1 U446 ( .A(G15GAT), .B(G190GAT), .ZN(n385) );
  XNOR2_X1 U447 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U448 ( .A(n387), .B(G134GAT), .Z(n390) );
  XNOR2_X1 U449 ( .A(G43GAT), .B(n388), .ZN(n389) );
  XNOR2_X1 U450 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U451 ( .A(n392), .B(n391), .ZN(n401) );
  XOR2_X1 U452 ( .A(G176GAT), .B(G183GAT), .Z(n394) );
  NAND2_X1 U453 ( .A1(G227GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U454 ( .A(n394), .B(n393), .ZN(n396) );
  XNOR2_X1 U455 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n395) );
  XNOR2_X1 U456 ( .A(n395), .B(G127GAT), .ZN(n413) );
  XOR2_X1 U457 ( .A(n396), .B(n413), .Z(n399) );
  XNOR2_X1 U458 ( .A(G169GAT), .B(n397), .ZN(n398) );
  XNOR2_X1 U459 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U460 ( .A(n401), .B(n400), .ZN(n480) );
  NAND2_X1 U461 ( .A1(n539), .A2(n480), .ZN(n423) );
  XOR2_X1 U462 ( .A(KEYINPUT6), .B(G57GAT), .Z(n403) );
  XNOR2_X1 U463 ( .A(G1GAT), .B(G120GAT), .ZN(n402) );
  XNOR2_X1 U464 ( .A(n403), .B(n402), .ZN(n407) );
  XOR2_X1 U465 ( .A(KEYINPUT97), .B(KEYINPUT5), .Z(n405) );
  XNOR2_X1 U466 ( .A(KEYINPUT4), .B(KEYINPUT1), .ZN(n404) );
  XNOR2_X1 U467 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U468 ( .A(n407), .B(n406), .Z(n412) );
  XOR2_X1 U469 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n409) );
  NAND2_X1 U470 ( .A1(G225GAT), .A2(G233GAT), .ZN(n408) );
  XNOR2_X1 U471 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U472 ( .A(KEYINPUT100), .B(n410), .ZN(n411) );
  XNOR2_X1 U473 ( .A(n412), .B(n411), .ZN(n422) );
  XOR2_X1 U474 ( .A(G85GAT), .B(G148GAT), .Z(n415) );
  XNOR2_X1 U475 ( .A(G29GAT), .B(n413), .ZN(n414) );
  XNOR2_X1 U476 ( .A(n415), .B(n414), .ZN(n417) );
  XNOR2_X1 U477 ( .A(G134GAT), .B(G162GAT), .ZN(n416) );
  XNOR2_X1 U478 ( .A(n416), .B(KEYINPUT80), .ZN(n436) );
  XOR2_X1 U479 ( .A(n417), .B(n436), .Z(n420) );
  XNOR2_X1 U480 ( .A(G141GAT), .B(n418), .ZN(n419) );
  XNOR2_X1 U481 ( .A(n420), .B(n419), .ZN(n421) );
  NAND2_X1 U482 ( .A1(n423), .A2(n573), .ZN(n432) );
  INV_X1 U483 ( .A(n480), .ZN(n537) );
  NAND2_X1 U484 ( .A1(n537), .A2(n529), .ZN(n424) );
  NAND2_X1 U485 ( .A1(n474), .A2(n424), .ZN(n425) );
  XNOR2_X1 U486 ( .A(KEYINPUT25), .B(n425), .ZN(n426) );
  NOR2_X1 U487 ( .A1(n573), .A2(n426), .ZN(n430) );
  NOR2_X1 U488 ( .A1(n474), .A2(n537), .ZN(n427) );
  XNOR2_X1 U489 ( .A(n427), .B(KEYINPUT26), .ZN(n574) );
  INV_X1 U490 ( .A(n428), .ZN(n429) );
  NAND2_X1 U491 ( .A1(n574), .A2(n429), .ZN(n553) );
  NAND2_X1 U492 ( .A1(n430), .A2(n553), .ZN(n431) );
  NAND2_X1 U493 ( .A1(n432), .A2(n431), .ZN(n491) );
  NOR2_X1 U494 ( .A1(n545), .A2(n491), .ZN(n434) );
  XNOR2_X1 U495 ( .A(n434), .B(n433), .ZN(n452) );
  XOR2_X1 U496 ( .A(n435), .B(KEYINPUT81), .Z(n440) );
  XOR2_X1 U497 ( .A(n436), .B(KEYINPUT11), .Z(n438) );
  NAND2_X1 U498 ( .A1(G232GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U499 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U500 ( .A(n440), .B(n439), .ZN(n449) );
  XOR2_X1 U501 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n442) );
  XNOR2_X1 U502 ( .A(KEYINPUT66), .B(KEYINPUT65), .ZN(n441) );
  XNOR2_X1 U503 ( .A(n442), .B(n441), .ZN(n447) );
  XNOR2_X1 U504 ( .A(KEYINPUT79), .B(n443), .ZN(n445) );
  XOR2_X1 U505 ( .A(KEYINPUT67), .B(KEYINPUT78), .Z(n444) );
  XNOR2_X1 U506 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U507 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U508 ( .A(n449), .B(n448), .ZN(n451) );
  XNOR2_X1 U509 ( .A(n451), .B(n450), .ZN(n565) );
  XNOR2_X1 U510 ( .A(KEYINPUT36), .B(n549), .ZN(n586) );
  NAND2_X1 U511 ( .A1(n452), .A2(n586), .ZN(n453) );
  XOR2_X1 U512 ( .A(KEYINPUT37), .B(n453), .Z(n527) );
  XNOR2_X1 U513 ( .A(n454), .B(KEYINPUT38), .ZN(n513) );
  NAND2_X1 U514 ( .A1(n513), .A2(n537), .ZN(n458) );
  XOR2_X1 U515 ( .A(KEYINPUT40), .B(KEYINPUT112), .Z(n456) );
  INV_X1 U516 ( .A(G43GAT), .ZN(n455) );
  XNOR2_X1 U517 ( .A(KEYINPUT55), .B(KEYINPUT122), .ZN(n478) );
  XOR2_X1 U518 ( .A(n579), .B(KEYINPUT64), .Z(n459) );
  XNOR2_X1 U519 ( .A(n459), .B(KEYINPUT41), .ZN(n557) );
  NOR2_X1 U520 ( .A1(n557), .A2(n576), .ZN(n460) );
  XNOR2_X1 U521 ( .A(n460), .B(KEYINPUT46), .ZN(n461) );
  NOR2_X1 U522 ( .A1(n545), .A2(n461), .ZN(n462) );
  NAND2_X1 U523 ( .A1(n462), .A2(n565), .ZN(n463) );
  XNOR2_X1 U524 ( .A(n463), .B(KEYINPUT47), .ZN(n469) );
  NAND2_X1 U525 ( .A1(n545), .A2(n586), .ZN(n465) );
  NAND2_X1 U526 ( .A1(n466), .A2(n579), .ZN(n467) );
  NOR2_X1 U527 ( .A1(n467), .A2(n567), .ZN(n468) );
  NOR2_X1 U528 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U529 ( .A(n470), .B(KEYINPUT48), .ZN(n554) );
  XNOR2_X1 U530 ( .A(KEYINPUT121), .B(n529), .ZN(n471) );
  NOR2_X1 U531 ( .A1(n554), .A2(n471), .ZN(n473) );
  INV_X1 U532 ( .A(KEYINPUT54), .ZN(n472) );
  XNOR2_X1 U533 ( .A(n473), .B(n472), .ZN(n572) );
  INV_X1 U534 ( .A(n573), .ZN(n475) );
  NAND2_X1 U535 ( .A1(n475), .A2(n474), .ZN(n476) );
  NOR2_X1 U536 ( .A1(n572), .A2(n476), .ZN(n477) );
  XNOR2_X1 U537 ( .A(n478), .B(n477), .ZN(n479) );
  INV_X1 U538 ( .A(n557), .ZN(n542) );
  NAND2_X1 U539 ( .A1(n568), .A2(n542), .ZN(n483) );
  XOR2_X1 U540 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n481) );
  XNOR2_X1 U541 ( .A(n481), .B(G176GAT), .ZN(n482) );
  XNOR2_X1 U542 ( .A(n483), .B(n482), .ZN(G1349GAT) );
  NAND2_X1 U543 ( .A1(n568), .A2(n549), .ZN(n486) );
  XOR2_X1 U544 ( .A(KEYINPUT58), .B(KEYINPUT125), .Z(n484) );
  NAND2_X1 U545 ( .A1(n568), .A2(n545), .ZN(n489) );
  XOR2_X1 U546 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n487) );
  XNOR2_X1 U547 ( .A(n487), .B(G183GAT), .ZN(n488) );
  XNOR2_X1 U548 ( .A(n489), .B(n488), .ZN(G1350GAT) );
  XNOR2_X1 U549 ( .A(KEYINPUT104), .B(KEYINPUT34), .ZN(n499) );
  XOR2_X1 U550 ( .A(G1GAT), .B(KEYINPUT105), .Z(n497) );
  INV_X1 U551 ( .A(n545), .ZN(n582) );
  NOR2_X1 U552 ( .A1(n549), .A2(n582), .ZN(n490) );
  XNOR2_X1 U553 ( .A(KEYINPUT16), .B(n490), .ZN(n493) );
  INV_X1 U554 ( .A(n491), .ZN(n492) );
  NAND2_X1 U555 ( .A1(n493), .A2(n492), .ZN(n515) );
  NOR2_X1 U556 ( .A1(n494), .A2(n515), .ZN(n495) );
  XOR2_X1 U557 ( .A(KEYINPUT103), .B(n495), .Z(n504) );
  NAND2_X1 U558 ( .A1(n504), .A2(n573), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U560 ( .A(n499), .B(n498), .ZN(G1324GAT) );
  NAND2_X1 U561 ( .A1(n529), .A2(n504), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n500), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U563 ( .A(KEYINPUT106), .B(KEYINPUT35), .Z(n502) );
  NAND2_X1 U564 ( .A1(n504), .A2(n537), .ZN(n501) );
  XNOR2_X1 U565 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U566 ( .A(G15GAT), .B(n503), .ZN(G1326GAT) );
  XOR2_X1 U567 ( .A(G22GAT), .B(KEYINPUT107), .Z(n506) );
  NAND2_X1 U568 ( .A1(n504), .A2(n532), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n506), .B(n505), .ZN(G1327GAT) );
  XNOR2_X1 U570 ( .A(KEYINPUT108), .B(KEYINPUT39), .ZN(n510) );
  XOR2_X1 U571 ( .A(G29GAT), .B(KEYINPUT110), .Z(n508) );
  NAND2_X1 U572 ( .A1(n513), .A2(n573), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U574 ( .A(n510), .B(n509), .ZN(G1328GAT) );
  XOR2_X1 U575 ( .A(G36GAT), .B(KEYINPUT111), .Z(n512) );
  NAND2_X1 U576 ( .A1(n513), .A2(n529), .ZN(n511) );
  XNOR2_X1 U577 ( .A(n512), .B(n511), .ZN(G1329GAT) );
  NAND2_X1 U578 ( .A1(n513), .A2(n532), .ZN(n514) );
  XNOR2_X1 U579 ( .A(n514), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT113), .B(KEYINPUT42), .Z(n517) );
  NAND2_X1 U581 ( .A1(n576), .A2(n542), .ZN(n526) );
  NOR2_X1 U582 ( .A1(n526), .A2(n515), .ZN(n522) );
  NAND2_X1 U583 ( .A1(n522), .A2(n573), .ZN(n516) );
  XNOR2_X1 U584 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U585 ( .A(G57GAT), .B(n518), .ZN(G1332GAT) );
  NAND2_X1 U586 ( .A1(n529), .A2(n522), .ZN(n519) );
  XNOR2_X1 U587 ( .A(n519), .B(KEYINPUT114), .ZN(n520) );
  XNOR2_X1 U588 ( .A(G64GAT), .B(n520), .ZN(G1333GAT) );
  NAND2_X1 U589 ( .A1(n537), .A2(n522), .ZN(n521) );
  XNOR2_X1 U590 ( .A(n521), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT43), .B(KEYINPUT115), .Z(n524) );
  NAND2_X1 U592 ( .A1(n522), .A2(n532), .ZN(n523) );
  XNOR2_X1 U593 ( .A(n524), .B(n523), .ZN(n525) );
  XOR2_X1 U594 ( .A(G78GAT), .B(n525), .Z(G1335GAT) );
  NOR2_X1 U595 ( .A1(n527), .A2(n526), .ZN(n533) );
  NAND2_X1 U596 ( .A1(n533), .A2(n573), .ZN(n528) );
  XNOR2_X1 U597 ( .A(G85GAT), .B(n528), .ZN(G1336GAT) );
  NAND2_X1 U598 ( .A1(n529), .A2(n533), .ZN(n530) );
  XNOR2_X1 U599 ( .A(n530), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U600 ( .A1(n537), .A2(n533), .ZN(n531) );
  XNOR2_X1 U601 ( .A(n531), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT116), .B(KEYINPUT44), .Z(n535) );
  NAND2_X1 U603 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U604 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U605 ( .A(G106GAT), .B(n536), .Z(G1339GAT) );
  AND2_X1 U606 ( .A1(n537), .A2(n573), .ZN(n538) );
  NAND2_X1 U607 ( .A1(n539), .A2(n538), .ZN(n540) );
  NOR2_X1 U608 ( .A1(n554), .A2(n540), .ZN(n550) );
  NAND2_X1 U609 ( .A1(n567), .A2(n550), .ZN(n541) );
  XNOR2_X1 U610 ( .A(G113GAT), .B(n541), .ZN(G1340GAT) );
  XOR2_X1 U611 ( .A(G120GAT), .B(KEYINPUT49), .Z(n544) );
  NAND2_X1 U612 ( .A1(n550), .A2(n542), .ZN(n543) );
  XNOR2_X1 U613 ( .A(n544), .B(n543), .ZN(G1341GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n547) );
  NAND2_X1 U615 ( .A1(n550), .A2(n545), .ZN(n546) );
  XNOR2_X1 U616 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U617 ( .A(G127GAT), .B(n548), .Z(G1342GAT) );
  XOR2_X1 U618 ( .A(G134GAT), .B(KEYINPUT51), .Z(n552) );
  NAND2_X1 U619 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U620 ( .A(n552), .B(n551), .ZN(G1343GAT) );
  NOR2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n555) );
  NAND2_X1 U622 ( .A1(n555), .A2(n573), .ZN(n564) );
  NOR2_X1 U623 ( .A1(n576), .A2(n564), .ZN(n556) );
  XOR2_X1 U624 ( .A(G141GAT), .B(n556), .Z(G1344GAT) );
  NOR2_X1 U625 ( .A1(n564), .A2(n557), .ZN(n561) );
  XOR2_X1 U626 ( .A(KEYINPUT53), .B(KEYINPUT119), .Z(n559) );
  XNOR2_X1 U627 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n558) );
  XNOR2_X1 U628 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U629 ( .A(n561), .B(n560), .ZN(G1345GAT) );
  NOR2_X1 U630 ( .A1(n582), .A2(n564), .ZN(n562) );
  XOR2_X1 U631 ( .A(KEYINPUT120), .B(n562), .Z(n563) );
  XNOR2_X1 U632 ( .A(G155GAT), .B(n563), .ZN(G1346GAT) );
  NOR2_X1 U633 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U634 ( .A(G162GAT), .B(n566), .Z(G1347GAT) );
  NAND2_X1 U635 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n569), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n571) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n570) );
  XNOR2_X1 U639 ( .A(n571), .B(n570), .ZN(n578) );
  NOR2_X1 U640 ( .A1(n573), .A2(n572), .ZN(n575) );
  NAND2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n585) );
  NOR2_X1 U642 ( .A1(n576), .A2(n585), .ZN(n577) );
  XOR2_X1 U643 ( .A(n578), .B(n577), .Z(G1352GAT) );
  NOR2_X1 U644 ( .A1(n579), .A2(n585), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1353GAT) );
  NOR2_X1 U647 ( .A1(n582), .A2(n585), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G211GAT), .B(KEYINPUT127), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1354GAT) );
  INV_X1 U650 ( .A(n585), .ZN(n587) );
  NAND2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U652 ( .A(n588), .B(KEYINPUT62), .ZN(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

