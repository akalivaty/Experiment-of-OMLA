//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 1 0 1 1 0 1 0 0 0 0 0 1 1 0 0 0 0 0 1 1 1 1 1 0 0 0 0 0 0 1 0 1 1 0 1 1 0 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:28 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n434, new_n437, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n569, new_n570, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n623,
    new_n624, new_n627, new_n629, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n840, new_n841, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT66), .B(G44), .Z(new_n434));
  INV_X1    g009(.A(new_n434), .ZN(G218));
  INV_X1    g010(.A(G132), .ZN(G219));
  XOR2_X1   g011(.A(KEYINPUT0), .B(G82), .Z(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT67), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n434), .A2(new_n437), .A3(G96), .A4(G132), .ZN(new_n453));
  INV_X1    g028(.A(KEYINPUT2), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(new_n455), .ZN(new_n459));
  INV_X1    g034(.A(new_n456), .ZN(new_n460));
  AOI22_X1  g035(.A1(new_n459), .A2(G2106), .B1(G567), .B2(new_n460), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT68), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  OAI211_X1 g041(.A(G137), .B(new_n464), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n464), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g045(.A(G125), .B1(new_n465), .B2(new_n466), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(KEYINPUT69), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n473));
  OAI211_X1 g048(.A(new_n473), .B(G125), .C1(new_n465), .C2(new_n466), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n472), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n470), .B1(new_n476), .B2(G2105), .ZN(G160));
  OR2_X1    g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n464), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n484), .B1(G112), .B2(new_n464), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT70), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n465), .A2(new_n466), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(new_n464), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  AOI211_X1 g065(.A(new_n482), .B(new_n486), .C1(G136), .C2(new_n490), .ZN(G162));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n493), .B1(new_n465), .B2(new_n466), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT72), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n493), .B(KEYINPUT72), .C1(new_n466), .C2(new_n465), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n496), .A2(KEYINPUT4), .A3(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT71), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT71), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G114), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G2105), .ZN(new_n504));
  OAI21_X1  g079(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n504), .A2(new_n506), .B1(new_n480), .B2(G126), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT4), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n494), .A2(new_n495), .A3(new_n508), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n498), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(G164));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT73), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g090(.A1(KEYINPUT73), .A2(KEYINPUT6), .A3(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n518), .B1(new_n519), .B2(KEYINPUT74), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT74), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n521), .A2(KEYINPUT5), .A3(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n517), .A2(G88), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n517), .A2(G50), .A3(G543), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT75), .ZN(new_n526));
  AND3_X1   g101(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n526), .B1(new_n524), .B2(new_n525), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n523), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n529));
  OAI22_X1  g104(.A1(new_n527), .A2(new_n528), .B1(new_n514), .B2(new_n529), .ZN(G303));
  INV_X1    g105(.A(G303), .ZN(G166));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n517), .A2(new_n523), .ZN(new_n534));
  INV_X1    g109(.A(G89), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT78), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n523), .A2(G63), .A3(G651), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n517), .A2(KEYINPUT76), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT76), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n515), .A2(new_n540), .A3(new_n516), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n539), .A2(G543), .A3(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(G51), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n538), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT77), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI211_X1 g121(.A(KEYINPUT77), .B(new_n538), .C1(new_n542), .C2(new_n543), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n537), .A2(new_n546), .A3(new_n547), .ZN(G286));
  INV_X1    g123(.A(G286), .ZN(G168));
  NOR2_X1   g124(.A1(KEYINPUT79), .A2(G52), .ZN(new_n550));
  AND2_X1   g125(.A1(KEYINPUT79), .A2(G52), .ZN(new_n551));
  NOR3_X1   g126(.A1(new_n542), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n523), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G90), .ZN(new_n554));
  OAI22_X1  g129(.A1(new_n553), .A2(new_n514), .B1(new_n534), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n552), .A2(new_n555), .ZN(G171));
  NAND2_X1  g131(.A1(G68), .A2(G543), .ZN(new_n557));
  AND2_X1   g132(.A1(new_n520), .A2(new_n522), .ZN(new_n558));
  INV_X1    g133(.A(G56), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G651), .ZN(new_n561));
  AND2_X1   g136(.A1(new_n517), .A2(new_n523), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G81), .ZN(new_n563));
  INV_X1    g138(.A(G43), .ZN(new_n564));
  OAI211_X1 g139(.A(new_n561), .B(new_n563), .C1(new_n564), .C2(new_n542), .ZN(new_n565));
  INV_X1    g140(.A(G860), .ZN(new_n566));
  OR2_X1    g141(.A1(new_n565), .A2(new_n566), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND4_X1  g145(.A1(G319), .A2(G483), .A3(G661), .A4(new_n570), .ZN(G188));
  NAND4_X1  g146(.A1(new_n539), .A2(G53), .A3(G543), .A4(new_n541), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(KEYINPUT9), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n519), .B1(new_n517), .B2(KEYINPUT76), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n574), .A2(new_n575), .A3(G53), .A4(new_n541), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(G78), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(G65), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n558), .B2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n580), .A2(G651), .B1(new_n562), .B2(G91), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n577), .A2(new_n581), .ZN(G299));
  INV_X1    g157(.A(G171), .ZN(G301));
  OAI21_X1  g158(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n584));
  INV_X1    g159(.A(G87), .ZN(new_n585));
  INV_X1    g160(.A(G49), .ZN(new_n586));
  OAI221_X1 g161(.A(new_n584), .B1(new_n585), .B2(new_n534), .C1(new_n542), .C2(new_n586), .ZN(G288));
  AOI21_X1  g162(.A(new_n519), .B1(new_n515), .B2(new_n516), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(G48), .ZN(new_n589));
  INV_X1    g164(.A(G86), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n590), .B2(new_n534), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT80), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n523), .A2(new_n592), .A3(G61), .ZN(new_n593));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT81), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n592), .B1(new_n523), .B2(G61), .ZN(new_n597));
  OAI21_X1  g172(.A(G651), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT82), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n591), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  OAI211_X1 g175(.A(KEYINPUT82), .B(G651), .C1(new_n596), .C2(new_n597), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(G305));
  NAND2_X1  g177(.A1(new_n562), .A2(G85), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n604));
  INV_X1    g179(.A(G47), .ZN(new_n605));
  OAI221_X1 g180(.A(new_n603), .B1(new_n514), .B2(new_n604), .C1(new_n542), .C2(new_n605), .ZN(G290));
  NAND2_X1  g181(.A1(G301), .A2(G868), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT83), .ZN(new_n608));
  AND3_X1   g183(.A1(new_n562), .A2(KEYINPUT10), .A3(G92), .ZN(new_n609));
  AOI21_X1  g184(.A(KEYINPUT10), .B1(new_n562), .B2(G92), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(G54), .ZN(new_n612));
  XOR2_X1   g187(.A(KEYINPUT84), .B(G66), .Z(new_n613));
  AOI22_X1  g188(.A1(new_n613), .A2(new_n523), .B1(G79), .B2(G543), .ZN(new_n614));
  OAI22_X1  g189(.A1(new_n542), .A2(new_n612), .B1(new_n514), .B2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT85), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  OAI221_X1 g192(.A(KEYINPUT85), .B1(new_n614), .B2(new_n514), .C1(new_n542), .C2(new_n612), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n611), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n608), .B1(G868), .B2(new_n619), .ZN(G284));
  OAI21_X1  g195(.A(new_n608), .B1(G868), .B2(new_n619), .ZN(G321));
  INV_X1    g196(.A(G868), .ZN(new_n622));
  NOR2_X1   g197(.A1(G286), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(G299), .B(KEYINPUT86), .Z(new_n624));
  AOI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(new_n622), .ZN(G297));
  AOI21_X1  g200(.A(new_n623), .B1(new_n624), .B2(new_n622), .ZN(G280));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n619), .B1(new_n627), .B2(G860), .ZN(G148));
  AOI21_X1  g203(.A(new_n622), .B1(new_n619), .B2(new_n627), .ZN(new_n629));
  INV_X1    g204(.A(KEYINPUT87), .ZN(new_n630));
  AOI22_X1  g205(.A1(new_n629), .A2(new_n630), .B1(new_n622), .B2(new_n565), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(new_n630), .B2(new_n629), .ZN(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g208(.A1(new_n488), .A2(new_n468), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT12), .Z(new_n635));
  XOR2_X1   g210(.A(KEYINPUT88), .B(KEYINPUT13), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(G2100), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n480), .A2(G123), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n464), .A2(G111), .ZN(new_n642));
  OAI21_X1  g217(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n643));
  INV_X1    g218(.A(G135), .ZN(new_n644));
  OAI221_X1 g219(.A(new_n641), .B1(new_n642), .B2(new_n643), .C1(new_n489), .C2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(G2096), .Z(new_n646));
  NAND3_X1  g221(.A1(new_n639), .A2(new_n640), .A3(new_n646), .ZN(G156));
  INV_X1    g222(.A(KEYINPUT14), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2427), .B(G2438), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2430), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT15), .B(G2435), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n648), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n652), .B1(new_n651), .B2(new_n650), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2451), .B(G2454), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n653), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2443), .B(G2446), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n660), .A2(G14), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n658), .A2(new_n659), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n663), .A2(KEYINPUT89), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(KEYINPUT89), .ZN(new_n665));
  AND2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(G401));
  XOR2_X1   g241(.A(G2072), .B(G2078), .Z(new_n667));
  XOR2_X1   g242(.A(G2084), .B(G2090), .Z(new_n668));
  XNOR2_X1  g243(.A(G2067), .B(G2678), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n667), .B1(new_n670), .B2(KEYINPUT18), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT90), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2096), .B(G2100), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(KEYINPUT18), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n670), .A2(KEYINPUT17), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n668), .A2(new_n669), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n675), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT91), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n674), .B(new_n679), .ZN(G227));
  XOR2_X1   g255(.A(G1971), .B(G1976), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  XOR2_X1   g257(.A(G1956), .B(G2474), .Z(new_n683));
  XOR2_X1   g258(.A(G1961), .B(G1966), .Z(new_n684));
  AND2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT20), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n683), .A2(new_n684), .ZN(new_n688));
  NOR3_X1   g263(.A1(new_n682), .A2(new_n685), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(new_n682), .B2(new_n688), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(G1991), .B(G1996), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n693), .A2(new_n694), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n693), .A2(new_n694), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n699), .A2(new_n696), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(G229));
  INV_X1    g278(.A(G29), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G26), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT28), .ZN(new_n706));
  OAI21_X1  g281(.A(KEYINPUT95), .B1(G104), .B2(G2105), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  NOR3_X1   g283(.A1(KEYINPUT95), .A2(G104), .A3(G2105), .ZN(new_n709));
  OAI221_X1 g284(.A(G2104), .B1(G116), .B2(new_n464), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n480), .ZN(new_n711));
  INV_X1    g286(.A(G128), .ZN(new_n712));
  INV_X1    g287(.A(G140), .ZN(new_n713));
  OAI221_X1 g288(.A(new_n710), .B1(new_n711), .B2(new_n712), .C1(new_n489), .C2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n706), .B1(new_n715), .B2(new_n704), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT96), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(G2067), .ZN(new_n718));
  MUX2_X1   g293(.A(G19), .B(new_n565), .S(G16), .Z(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(G1341), .Z(new_n720));
  NAND2_X1  g295(.A1(new_n619), .A2(G16), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G4), .B2(G16), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT94), .B(G1348), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  OAI211_X1 g299(.A(new_n718), .B(new_n720), .C1(new_n722), .C2(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(new_n722), .B2(new_n724), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n726), .A2(KEYINPUT97), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(KEYINPUT97), .ZN(new_n728));
  INV_X1    g303(.A(G32), .ZN(new_n729));
  AOI21_X1  g304(.A(KEYINPUT99), .B1(new_n704), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n490), .A2(G141), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  AND2_X1   g307(.A1(new_n468), .A2(G105), .ZN(new_n733));
  NAND3_X1  g308(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT26), .Z(new_n735));
  INV_X1    g310(.A(G129), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n735), .B1(new_n711), .B2(new_n736), .ZN(new_n737));
  NOR3_X1   g312(.A1(new_n732), .A2(new_n733), .A3(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n730), .B1(new_n739), .B2(new_n704), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n738), .A2(KEYINPUT99), .A3(G29), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XOR2_X1   g317(.A(KEYINPUT27), .B(G1996), .Z(new_n743));
  NOR2_X1   g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT100), .Z(new_n745));
  NOR2_X1   g320(.A1(G29), .A2(G35), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(G162), .B2(G29), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT101), .B(KEYINPUT29), .Z(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G2090), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n747), .B(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(G16), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(G5), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G171), .B2(new_n751), .ZN(new_n753));
  INV_X1    g328(.A(G2072), .ZN(new_n754));
  NOR2_X1   g329(.A1(G29), .A2(G33), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT98), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT25), .ZN(new_n757));
  NAND2_X1  g332(.A1(G103), .A2(G2104), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n757), .B1(new_n758), .B2(G2105), .ZN(new_n759));
  NAND4_X1  g334(.A1(new_n464), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n760));
  AOI22_X1  g335(.A1(new_n490), .A2(G139), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n488), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n761), .B1(new_n464), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n756), .B1(new_n763), .B2(new_n704), .ZN(new_n764));
  OAI221_X1 g339(.A(new_n750), .B1(G1961), .B2(new_n753), .C1(new_n754), .C2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(G160), .A2(G29), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT24), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n767), .A2(G34), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n704), .B1(new_n767), .B2(G34), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n766), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(G2084), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n753), .A2(G1961), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(new_n771), .B2(new_n770), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT30), .B(G28), .ZN(new_n774));
  OR2_X1    g349(.A1(KEYINPUT31), .A2(G11), .ZN(new_n775));
  NAND2_X1  g350(.A1(KEYINPUT31), .A2(G11), .ZN(new_n776));
  AOI22_X1  g351(.A1(new_n774), .A2(new_n704), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n645), .B2(new_n704), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n764), .A2(new_n754), .ZN(new_n779));
  AOI211_X1 g354(.A(new_n778), .B(new_n779), .C1(new_n742), .C2(new_n743), .ZN(new_n780));
  NOR2_X1   g355(.A1(G27), .A2(G29), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G164), .B2(G29), .ZN(new_n782));
  INV_X1    g357(.A(G2078), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n780), .A2(new_n784), .ZN(new_n785));
  NOR4_X1   g360(.A1(new_n745), .A2(new_n765), .A3(new_n773), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n751), .A2(G21), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G168), .B2(new_n751), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G1966), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n751), .A2(G20), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT23), .Z(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G299), .B2(G16), .ZN(new_n792));
  INV_X1    g367(.A(G1956), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n789), .A2(new_n794), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n727), .A2(new_n728), .A3(new_n786), .A4(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT93), .ZN(new_n797));
  NAND2_X1  g372(.A1(G288), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n584), .B1(new_n534), .B2(new_n585), .ZN(new_n799));
  INV_X1    g374(.A(new_n542), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(G49), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n801), .A2(KEYINPUT93), .ZN(new_n802));
  AND2_X1   g377(.A1(new_n798), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n803), .A2(G16), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G16), .B2(G23), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT33), .B(G1976), .ZN(new_n806));
  AND2_X1   g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g382(.A1(G6), .A2(G16), .ZN(new_n808));
  INV_X1    g383(.A(G305), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n808), .B1(new_n809), .B2(G16), .ZN(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT32), .B(G1981), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n805), .A2(new_n806), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n751), .A2(G22), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(G166), .B2(new_n751), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(G1971), .ZN(new_n816));
  NOR4_X1   g391(.A1(new_n807), .A2(new_n812), .A3(new_n813), .A4(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT34), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n817), .A2(new_n818), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n480), .A2(G119), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n464), .A2(G107), .ZN(new_n822));
  OAI21_X1  g397(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n823));
  INV_X1    g398(.A(G131), .ZN(new_n824));
  OAI221_X1 g399(.A(new_n821), .B1(new_n822), .B2(new_n823), .C1(new_n489), .C2(new_n824), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT92), .Z(new_n826));
  MUX2_X1   g401(.A(G25), .B(new_n826), .S(G29), .Z(new_n827));
  XOR2_X1   g402(.A(KEYINPUT35), .B(G1991), .Z(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n827), .B(new_n829), .ZN(new_n830));
  MUX2_X1   g405(.A(G24), .B(G290), .S(G16), .Z(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(G1986), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n819), .A2(new_n820), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(KEYINPUT36), .ZN(new_n835));
  AND2_X1   g410(.A1(new_n820), .A2(new_n833), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT36), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n836), .A2(new_n837), .A3(new_n819), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n796), .B1(new_n835), .B2(new_n838), .ZN(G311));
  AND4_X1   g414(.A1(new_n727), .A2(new_n786), .A3(new_n728), .A4(new_n795), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n837), .B1(new_n836), .B2(new_n819), .ZN(new_n841));
  AND4_X1   g416(.A1(new_n837), .A2(new_n819), .A3(new_n820), .A4(new_n833), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n840), .B1(new_n841), .B2(new_n842), .ZN(G150));
  AND3_X1   g418(.A1(new_n574), .A2(G55), .A3(new_n541), .ZN(new_n844));
  AOI22_X1  g419(.A1(new_n523), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n845));
  INV_X1    g420(.A(G93), .ZN(new_n846));
  OAI22_X1  g421(.A1(new_n845), .A2(new_n514), .B1(new_n534), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n848), .A2(new_n566), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT37), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n619), .A2(G559), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT38), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n848), .B(new_n565), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n852), .B(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT39), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT102), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n855), .A2(new_n856), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(new_n566), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n850), .B1(new_n858), .B2(new_n860), .ZN(G145));
  XNOR2_X1  g436(.A(new_n714), .B(new_n510), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n763), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n863), .A2(new_n738), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n738), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n480), .A2(G130), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT103), .ZN(new_n869));
  OAI21_X1  g444(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n870));
  INV_X1    g445(.A(G118), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n870), .B1(new_n871), .B2(G2105), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n872), .B1(new_n490), .B2(G142), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT104), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(new_n635), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(new_n825), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n867), .A2(new_n877), .A3(KEYINPUT105), .ZN(new_n878));
  XOR2_X1   g453(.A(new_n645), .B(G160), .Z(new_n879));
  XOR2_X1   g454(.A(new_n879), .B(G162), .Z(new_n880));
  AND2_X1   g455(.A1(new_n876), .A2(new_n825), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n876), .A2(new_n825), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT105), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n883), .B1(new_n884), .B2(new_n866), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n867), .A2(KEYINPUT105), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n878), .B(new_n880), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(G37), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n866), .B1(new_n877), .B2(KEYINPUT106), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT106), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n883), .A2(new_n867), .A3(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n880), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n889), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n887), .A2(new_n888), .A3(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g470(.A1(new_n619), .A2(new_n627), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(new_n853), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(G299), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n619), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n619), .A2(new_n899), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n898), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(KEYINPUT41), .B1(new_n901), .B2(new_n902), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n617), .A2(new_n618), .ZN(new_n906));
  INV_X1    g481(.A(new_n611), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(G299), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT41), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n909), .A2(new_n910), .A3(new_n900), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n905), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(new_n897), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n904), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT108), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n904), .A2(KEYINPUT108), .A3(new_n913), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n798), .A2(new_n802), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n919), .B(G305), .ZN(new_n920));
  XNOR2_X1  g495(.A(G303), .B(G290), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n921), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n803), .A2(G305), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n809), .A2(new_n919), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n922), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(KEYINPUT107), .B(KEYINPUT42), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n927), .B(new_n928), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n918), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n929), .B1(new_n915), .B2(new_n914), .ZN(new_n931));
  OAI21_X1  g506(.A(G868), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n932), .B1(G868), .B2(new_n848), .ZN(G295));
  OAI21_X1  g508(.A(new_n932), .B1(G868), .B2(new_n848), .ZN(G331));
  NAND2_X1  g509(.A1(G286), .A2(G301), .ZN(new_n935));
  NAND4_X1  g510(.A1(G171), .A2(new_n537), .A3(new_n546), .A4(new_n547), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(new_n854), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n935), .A2(new_n853), .A3(new_n936), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n903), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT109), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n935), .A2(new_n853), .A3(KEYINPUT109), .A4(new_n936), .ZN(new_n943));
  AOI22_X1  g518(.A1(new_n942), .A2(new_n943), .B1(new_n854), .B2(new_n937), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n905), .A2(new_n911), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n927), .B(new_n940), .C1(new_n944), .C2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(new_n888), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n942), .A2(new_n943), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n938), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(new_n912), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n927), .B1(new_n950), .B2(new_n940), .ZN(new_n951));
  OAI21_X1  g526(.A(KEYINPUT43), .B1(new_n947), .B2(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n948), .A2(new_n903), .A3(new_n938), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n903), .A2(KEYINPUT110), .A3(new_n910), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n938), .A2(new_n939), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT110), .ZN(new_n957));
  AND3_X1   g532(.A1(new_n905), .A2(new_n957), .A3(new_n911), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n953), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n927), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT43), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n961), .A2(new_n962), .A3(new_n888), .A4(new_n946), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT44), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n952), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n955), .B(new_n954), .C1(new_n912), .C2(KEYINPUT110), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n927), .B1(new_n966), .B2(new_n953), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT43), .B1(new_n947), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(KEYINPUT111), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT111), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n970), .B(KEYINPUT43), .C1(new_n947), .C2(new_n967), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n946), .A2(new_n888), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n950), .A2(new_n940), .ZN(new_n973));
  OAI211_X1 g548(.A(new_n972), .B(new_n962), .C1(new_n927), .C2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n969), .A2(new_n971), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n965), .B1(new_n975), .B2(KEYINPUT44), .ZN(G397));
  NAND2_X1  g551(.A1(G303), .A2(G8), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT55), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n977), .B(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G1384), .ZN(new_n980));
  AND3_X1   g555(.A1(new_n496), .A2(KEYINPUT4), .A3(new_n497), .ZN(new_n981));
  XNOR2_X1  g556(.A(KEYINPUT71), .B(G114), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n506), .B1(new_n982), .B2(new_n464), .ZN(new_n983));
  OAI211_X1 g558(.A(G126), .B(G2105), .C1(new_n465), .C2(new_n466), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n509), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n980), .B1(new_n981), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT45), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT115), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n987), .A2(G1384), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n510), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G40), .ZN(new_n991));
  AOI211_X1 g566(.A(new_n991), .B(new_n470), .C1(new_n476), .C2(G2105), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n988), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n986), .A2(KEYINPUT115), .A3(new_n987), .ZN(new_n995));
  AOI21_X1  g570(.A(G1971), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  XNOR2_X1  g571(.A(KEYINPUT116), .B(KEYINPUT50), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n980), .B(new_n997), .C1(new_n981), .C2(new_n985), .ZN(new_n998));
  AND3_X1   g573(.A1(new_n494), .A2(new_n495), .A3(new_n508), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n464), .B1(new_n500), .B2(new_n502), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n984), .B1(new_n1000), .B2(new_n505), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(G1384), .B1(new_n1002), .B2(new_n498), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT50), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n992), .B(new_n998), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1005), .A2(G2090), .ZN(new_n1006));
  OAI211_X1 g581(.A(G8), .B(new_n979), .C1(new_n996), .C2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(KEYINPUT117), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT115), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1009), .B1(new_n1003), .B2(KEYINPUT45), .ZN(new_n1010));
  INV_X1    g585(.A(new_n989), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1011), .B1(new_n1002), .B2(new_n498), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n476), .A2(G2105), .ZN(new_n1013));
  INV_X1    g588(.A(new_n470), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1013), .A2(G40), .A3(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1010), .A2(new_n995), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G1971), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1019), .B1(G2090), .B2(new_n1005), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT117), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1020), .A2(new_n1021), .A3(G8), .A4(new_n979), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1008), .A2(new_n1022), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n510), .A2(G160), .A3(G40), .A4(new_n980), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(G8), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G1976), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT52), .B1(G288), .B2(new_n1027), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1026), .B(new_n1028), .C1(new_n919), .C2(new_n1027), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1025), .B1(new_n803), .B2(G1976), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1029), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n598), .A2(new_n599), .ZN(new_n1033));
  INV_X1    g608(.A(G1981), .ZN(new_n1034));
  INV_X1    g609(.A(new_n591), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1033), .A2(new_n1034), .A3(new_n601), .A4(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT118), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT118), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n600), .A2(new_n1038), .A3(new_n1034), .A4(new_n601), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(G305), .A2(G1981), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT49), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1025), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1040), .A2(KEYINPUT49), .A3(new_n1041), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1032), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(G8), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT119), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n990), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1012), .A2(KEYINPUT119), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT45), .B1(new_n510), .B2(new_n980), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1052), .A2(new_n1015), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(G1966), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1005), .A2(G2084), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  AOI211_X1 g633(.A(new_n1047), .B(G286), .C1(new_n1056), .C2(new_n1058), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1004), .B(new_n980), .C1(new_n981), .C2(new_n985), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n992), .B(new_n1060), .C1(new_n1003), .C2(new_n997), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1061), .A2(G2090), .ZN(new_n1062));
  OAI21_X1  g637(.A(G8), .B1(new_n996), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n979), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1023), .A2(new_n1046), .A3(new_n1059), .A4(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT63), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1006), .B1(new_n1018), .B2(new_n1017), .ZN(new_n1069));
  OAI21_X1  g644(.A(KEYINPUT120), .B1(new_n1069), .B2(new_n1047), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT120), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1071), .B(G8), .C1(new_n996), .C2(new_n1006), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1070), .A2(new_n1064), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1074), .A2(KEYINPUT63), .A3(G8), .A4(G168), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1023), .A2(new_n1046), .A3(new_n1073), .A4(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT121), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1075), .B1(new_n1008), .B2(new_n1022), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1080), .A2(KEYINPUT121), .A3(new_n1046), .A4(new_n1073), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1068), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1082));
  AOI211_X1 g657(.A(KEYINPUT60), .B(new_n611), .C1(new_n617), .C2(new_n618), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT122), .ZN(new_n1084));
  INV_X1    g659(.A(G2067), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1003), .A2(new_n992), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(G1348), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n998), .A2(new_n992), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1004), .B1(new_n510), .B2(new_n980), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1087), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT122), .B1(new_n1024), .B2(G2067), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1083), .A2(new_n1086), .A3(new_n1090), .A4(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(G1996), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1010), .A2(new_n1016), .A3(new_n1093), .A4(new_n995), .ZN(new_n1094));
  XOR2_X1   g669(.A(KEYINPUT58), .B(G1341), .Z(new_n1095));
  NAND2_X1  g670(.A1(new_n1024), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n565), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1092), .B1(new_n1097), .B2(KEYINPUT59), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT59), .ZN(new_n1099));
  AOI211_X1 g674(.A(new_n1099), .B(new_n565), .C1(new_n1094), .C2(new_n1096), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1090), .A2(new_n1086), .A3(new_n1091), .ZN(new_n1102));
  AND2_X1   g677(.A1(new_n1102), .A2(new_n619), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1102), .A2(new_n619), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT60), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g680(.A(KEYINPUT56), .B(G2072), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1010), .A2(new_n1016), .A3(new_n995), .A4(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1061), .A2(new_n793), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  OR2_X1    g684(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1110));
  NAND2_X1  g685(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1109), .A2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1107), .A2(new_n1110), .A3(new_n1108), .A4(new_n1111), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1113), .A2(KEYINPUT61), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT61), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1114), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n1107), .A2(new_n1108), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1116), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1101), .A2(new_n1105), .A3(new_n1115), .A4(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT123), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1102), .A2(new_n1121), .A3(new_n619), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(new_n1113), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1121), .B1(new_n1102), .B2(new_n619), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1114), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(KEYINPUT124), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT124), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1127), .B(new_n1114), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1120), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT54), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1010), .A2(new_n1016), .A3(new_n783), .A4(new_n995), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT53), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n1012), .A2(new_n1132), .A3(G2078), .ZN(new_n1134));
  INV_X1    g709(.A(G1961), .ZN(new_n1135));
  AOI22_X1  g710(.A1(new_n1053), .A2(new_n1134), .B1(new_n1005), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1133), .A2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1130), .B1(new_n1137), .B2(G171), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1005), .A2(new_n1135), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1051), .A2(new_n1053), .A3(KEYINPUT53), .A4(new_n783), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1133), .A2(G301), .A3(new_n1139), .A4(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT126), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  AND2_X1   g718(.A1(new_n1138), .A2(new_n1143), .ZN(new_n1144));
  OR2_X1    g719(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1056), .A2(G168), .A3(new_n1058), .ZN(new_n1146));
  AOI21_X1  g721(.A(G1966), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1147));
  OAI21_X1  g722(.A(G286), .B1(new_n1147), .B2(new_n1057), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1146), .A2(G8), .A3(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(KEYINPUT51), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT51), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1146), .A2(new_n1151), .A3(G8), .ZN(new_n1152));
  AOI22_X1  g727(.A1(new_n1144), .A2(new_n1145), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n1023), .A2(new_n1046), .A3(new_n1065), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1133), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(G171), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(KEYINPUT125), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT125), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1155), .A2(new_n1158), .A3(G171), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1133), .A2(new_n1136), .A3(G301), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1157), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(new_n1130), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1129), .A2(new_n1153), .A3(new_n1154), .A4(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(KEYINPUT62), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT62), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1150), .A2(new_n1167), .A3(new_n1152), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1165), .A2(new_n1154), .A3(new_n1166), .A4(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1170), .A2(new_n1027), .A3(new_n801), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1171), .A2(new_n1040), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1023), .ZN(new_n1173));
  AOI22_X1  g748(.A1(new_n1172), .A2(new_n1026), .B1(new_n1046), .B2(new_n1173), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1082), .A2(new_n1163), .A3(new_n1169), .A4(new_n1174), .ZN(new_n1175));
  OR3_X1    g750(.A1(G290), .A2(KEYINPUT112), .A3(G1986), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1052), .A2(new_n992), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1177), .ZN(new_n1178));
  OAI21_X1  g753(.A(KEYINPUT112), .B1(G290), .B2(G1986), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1176), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1178), .A2(G1986), .A3(G290), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  XOR2_X1   g757(.A(new_n1182), .B(KEYINPUT113), .Z(new_n1183));
  NAND3_X1  g758(.A1(new_n1178), .A2(new_n1093), .A3(new_n738), .ZN(new_n1184));
  XNOR2_X1  g759(.A(new_n1184), .B(KEYINPUT114), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n714), .B(new_n1085), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1186), .B1(new_n1093), .B2(new_n738), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1187), .A2(new_n1178), .ZN(new_n1188));
  XNOR2_X1  g763(.A(new_n825), .B(new_n828), .ZN(new_n1189));
  OAI211_X1 g764(.A(new_n1185), .B(new_n1188), .C1(new_n1177), .C2(new_n1189), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1183), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1175), .A2(new_n1191), .ZN(new_n1192));
  XOR2_X1   g767(.A(new_n1180), .B(KEYINPUT48), .Z(new_n1193));
  NOR2_X1   g768(.A1(new_n1190), .A2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n826), .A2(new_n829), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1185), .A2(new_n1188), .A3(new_n1195), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n715), .A2(new_n1085), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1177), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1177), .B1(new_n1186), .B2(new_n738), .ZN(new_n1199));
  OR3_X1    g774(.A1(new_n1177), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1200));
  OAI21_X1  g775(.A(KEYINPUT46), .B1(new_n1177), .B2(G1996), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n1199), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  XNOR2_X1  g777(.A(new_n1202), .B(KEYINPUT47), .ZN(new_n1203));
  NOR3_X1   g778(.A1(new_n1194), .A2(new_n1198), .A3(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1192), .A2(new_n1204), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g780(.A1(G227), .A2(new_n462), .ZN(new_n1207));
  AOI21_X1  g781(.A(new_n1207), .B1(new_n664), .B2(new_n665), .ZN(new_n1208));
  OAI21_X1  g782(.A(new_n702), .B1(KEYINPUT127), .B2(new_n1208), .ZN(new_n1209));
  AND2_X1   g783(.A1(new_n1208), .A2(KEYINPUT127), .ZN(new_n1210));
  NOR2_X1   g784(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g785(.A1(new_n952), .A2(new_n963), .ZN(new_n1212));
  NAND3_X1  g786(.A1(new_n1211), .A2(new_n894), .A3(new_n1212), .ZN(G225));
  INV_X1    g787(.A(G225), .ZN(G308));
endmodule


