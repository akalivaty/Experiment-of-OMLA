//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 0 1 1 1 0 1 1 0 0 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 0 0 1 1 0 1 1 0 0 1 1 1 0 1 1 0 1 0 0 1 0 0 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:25 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(KEYINPUT66), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G143), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(new_n187), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(KEYINPUT64), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT64), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G143), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(KEYINPUT66), .A3(G146), .ZN(new_n197));
  AND2_X1   g011(.A1(KEYINPUT0), .A2(G128), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n191), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n193), .A2(new_n195), .A3(new_n187), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT65), .B1(new_n187), .B2(G143), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT65), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(new_n192), .A3(G146), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n200), .A2(new_n201), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g018(.A1(KEYINPUT0), .A2(G128), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n198), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  AND2_X1   g021(.A1(new_n199), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G137), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n209), .A2(G134), .ZN(new_n210));
  INV_X1    g024(.A(G134), .ZN(new_n211));
  OAI21_X1  g025(.A(KEYINPUT11), .B1(new_n211), .B2(G137), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT11), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(new_n209), .A3(G134), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n210), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G131), .ZN(new_n216));
  OR2_X1    g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n212), .A2(new_n214), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n211), .A2(G137), .ZN(new_n219));
  AND4_X1   g033(.A1(KEYINPUT68), .A2(new_n218), .A3(new_n216), .A4(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(KEYINPUT68), .B1(new_n215), .B2(new_n216), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n217), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n208), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G128), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n224), .B1(new_n188), .B2(KEYINPUT1), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n191), .A2(new_n197), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n225), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n204), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n218), .A2(new_n216), .A3(new_n219), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n215), .A2(KEYINPUT68), .A3(new_n216), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(new_n219), .B(KEYINPUT69), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n211), .A2(G137), .ZN(new_n236));
  OAI21_X1  g050(.A(G131), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n229), .A2(new_n234), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT2), .ZN(new_n239));
  INV_X1    g053(.A(G113), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT70), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT70), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n242), .A2(KEYINPUT2), .A3(G113), .ZN(new_n243));
  AOI22_X1  g057(.A1(new_n241), .A2(new_n243), .B1(new_n239), .B2(new_n240), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT71), .ZN(new_n245));
  INV_X1    g059(.A(G119), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n245), .B1(new_n246), .B2(G116), .ZN(new_n247));
  INV_X1    g061(.A(G116), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n248), .A2(KEYINPUT71), .A3(G119), .ZN(new_n249));
  AOI22_X1  g063(.A1(new_n247), .A2(new_n249), .B1(G116), .B2(new_n246), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n244), .A2(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n244), .A2(new_n250), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n223), .A2(new_n238), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT28), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT28), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n223), .A2(new_n238), .A3(new_n256), .A4(new_n253), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n199), .A2(new_n207), .A3(KEYINPUT67), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n222), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(KEYINPUT67), .B1(new_n199), .B2(new_n207), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n238), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n253), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n258), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(G237), .ZN(new_n266));
  INV_X1    g080(.A(G953), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n266), .A2(new_n267), .A3(G210), .ZN(new_n268));
  INV_X1    g082(.A(G101), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n268), .B(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n270), .B(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n265), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n254), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n199), .A2(new_n207), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT67), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n277), .A2(new_n222), .A3(new_n259), .ZN(new_n278));
  AOI21_X1  g092(.A(KEYINPUT30), .B1(new_n278), .B2(new_n238), .ZN(new_n279));
  AND3_X1   g093(.A1(new_n223), .A2(KEYINPUT30), .A3(new_n238), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n274), .B1(new_n281), .B2(new_n263), .ZN(new_n282));
  INV_X1    g096(.A(new_n272), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT31), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT30), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n262), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n223), .A2(new_n238), .A3(KEYINPUT30), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(new_n263), .A3(new_n287), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n288), .A2(KEYINPUT31), .A3(new_n254), .A4(new_n283), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n273), .B1(new_n284), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G472), .ZN(new_n292));
  INV_X1    g106(.A(G902), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT32), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n283), .B1(new_n288), .B2(new_n254), .ZN(new_n297));
  AOI221_X4 g111(.A(new_n272), .B1(new_n262), .B2(new_n263), .C1(new_n255), .C2(new_n257), .ZN(new_n298));
  OAI21_X1  g112(.A(KEYINPUT72), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT29), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT72), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n301), .B1(new_n265), .B2(new_n272), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n299), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n253), .B1(new_n223), .B2(new_n238), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n304), .B1(new_n255), .B2(new_n257), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n305), .A2(KEYINPUT29), .A3(new_n283), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n293), .ZN(new_n307));
  OAI21_X1  g121(.A(G472), .B1(new_n303), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n288), .A2(new_n254), .A3(new_n283), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT31), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n289), .ZN(new_n312));
  AOI21_X1  g126(.A(G902), .B1(new_n312), .B2(new_n273), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n313), .A2(KEYINPUT32), .A3(new_n292), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n296), .A2(new_n308), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT73), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT73), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n296), .A2(new_n308), .A3(new_n317), .A4(new_n314), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G217), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n320), .B1(G234), .B2(new_n293), .ZN(new_n321));
  INV_X1    g135(.A(G140), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G125), .ZN(new_n323));
  INV_X1    g137(.A(G125), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G140), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT16), .ZN(new_n327));
  OR2_X1    g141(.A1(new_n323), .A2(KEYINPUT16), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n327), .A2(G146), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n326), .A2(new_n187), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n246), .A2(G128), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(KEYINPUT23), .B1(new_n224), .B2(G119), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n333), .B(KEYINPUT75), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT76), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n332), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT23), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n331), .B(new_n337), .C1(KEYINPUT75), .C2(KEYINPUT76), .ZN(new_n338));
  AOI21_X1  g152(.A(G110), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT74), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n224), .A2(G119), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n341), .A2(new_n340), .ZN(new_n342));
  MUX2_X1   g156(.A(new_n340), .B(new_n342), .S(new_n332), .Z(new_n343));
  XOR2_X1   g157(.A(KEYINPUT24), .B(G110), .Z(new_n344));
  NOR2_X1   g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n329), .B(new_n330), .C1(new_n339), .C2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n336), .A2(G110), .A3(new_n338), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n327), .A2(new_n328), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n187), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n329), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n343), .A2(new_n344), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n347), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(KEYINPUT22), .B(G137), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n267), .A2(G221), .A3(G234), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n353), .B(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n346), .A2(new_n352), .A3(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n346), .A2(new_n352), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(KEYINPUT77), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT77), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n346), .A2(new_n360), .A3(new_n352), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  XOR2_X1   g176(.A(new_n355), .B(KEYINPUT78), .Z(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n357), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(KEYINPUT25), .B1(new_n365), .B2(new_n293), .ZN(new_n366));
  INV_X1    g180(.A(new_n361), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n360), .B1(new_n346), .B2(new_n352), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n364), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  AND4_X1   g183(.A1(KEYINPUT25), .A2(new_n369), .A3(new_n293), .A4(new_n356), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n321), .B1(new_n366), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n365), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n321), .A2(G902), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n371), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  XOR2_X1   g190(.A(KEYINPUT9), .B(G234), .Z(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(G221), .B1(new_n378), .B2(G902), .ZN(new_n379));
  INV_X1    g193(.A(G469), .ZN(new_n380));
  XNOR2_X1  g194(.A(G110), .B(G140), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n267), .A2(G227), .ZN(new_n382));
  XOR2_X1   g196(.A(new_n381), .B(new_n382), .Z(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT82), .ZN(new_n385));
  INV_X1    g199(.A(G104), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n386), .A2(KEYINPUT3), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT80), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n388), .A2(G107), .ZN(new_n389));
  INV_X1    g203(.A(G107), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n390), .A2(KEYINPUT80), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n387), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n390), .A2(G104), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(KEYINPUT3), .B1(new_n386), .B2(G107), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(KEYINPUT79), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n390), .A2(G104), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT79), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n397), .A2(new_n398), .A3(KEYINPUT3), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n392), .A2(new_n394), .A3(new_n396), .A4(new_n399), .ZN(new_n400));
  XOR2_X1   g214(.A(KEYINPUT81), .B(G101), .Z(new_n401));
  OAI21_X1  g215(.A(new_n385), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  AND2_X1   g216(.A1(new_n396), .A2(new_n399), .ZN(new_n403));
  XOR2_X1   g217(.A(KEYINPUT80), .B(G107), .Z(new_n404));
  AOI21_X1  g218(.A(new_n393), .B1(new_n404), .B2(new_n387), .ZN(new_n405));
  INV_X1    g219(.A(new_n401), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n403), .A2(new_n405), .A3(KEYINPUT82), .A4(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n402), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n389), .A2(new_n391), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(new_n386), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n269), .B1(new_n410), .B2(new_n397), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n408), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n229), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n411), .B1(new_n402), .B2(new_n407), .ZN(new_n416));
  OR2_X1    g230(.A1(new_n226), .A2(KEYINPUT83), .ZN(new_n417));
  AND3_X1   g231(.A1(new_n196), .A2(KEYINPUT66), .A3(G146), .ZN(new_n418));
  AOI22_X1  g232(.A1(new_n196), .A2(G146), .B1(KEYINPUT66), .B2(new_n188), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT1), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n420), .B1(new_n190), .B2(new_n187), .ZN(new_n421));
  OAI22_X1  g235(.A1(new_n418), .A2(new_n419), .B1(new_n421), .B2(new_n224), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n422), .A2(KEYINPUT83), .A3(new_n226), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n416), .A2(new_n417), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n415), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(KEYINPUT12), .B1(new_n425), .B2(new_n222), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT12), .ZN(new_n427));
  INV_X1    g241(.A(new_n222), .ZN(new_n428));
  AOI211_X1 g242(.A(new_n427), .B(new_n428), .C1(new_n415), .C2(new_n424), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n269), .B1(new_n403), .B2(new_n405), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT4), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT4), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n433), .B1(new_n402), .B2(new_n407), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n432), .B1(new_n434), .B2(new_n431), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n208), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT10), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n424), .A2(new_n437), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n414), .A2(new_n437), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n416), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n436), .A2(new_n438), .A3(new_n428), .A4(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n384), .B1(new_n430), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n436), .A2(new_n438), .A3(new_n440), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n222), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n445), .A2(new_n441), .A3(new_n383), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT84), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n443), .A2(KEYINPUT84), .A3(new_n446), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n380), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  AOI22_X1  g265(.A1(new_n435), .A2(new_n208), .B1(new_n416), .B2(new_n439), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n428), .B1(new_n452), .B2(new_n438), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n384), .B1(new_n442), .B2(new_n453), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n441), .B(new_n383), .C1(new_n426), .C2(new_n429), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n456), .A2(new_n380), .A3(new_n293), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n380), .A2(new_n293), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n379), .B1(new_n451), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n266), .A2(new_n267), .A3(G143), .A4(G214), .ZN(new_n463));
  AND3_X1   g277(.A1(new_n266), .A2(new_n267), .A3(G214), .ZN(new_n464));
  OAI211_X1 g278(.A(KEYINPUT90), .B(new_n463), .C1(new_n190), .C2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT18), .ZN(new_n466));
  OAI21_X1  g280(.A(KEYINPUT91), .B1(new_n466), .B2(new_n216), .ZN(new_n467));
  OR2_X1    g281(.A1(new_n463), .A2(KEYINPUT90), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n465), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NOR3_X1   g283(.A1(new_n466), .A2(new_n216), .A3(KEYINPUT91), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n469), .B(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n323), .A2(new_n325), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(G146), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n330), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n329), .ZN(new_n475));
  XOR2_X1   g289(.A(KEYINPUT92), .B(KEYINPUT19), .Z(new_n476));
  NAND2_X1  g290(.A1(new_n326), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT92), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n472), .B1(new_n478), .B2(KEYINPUT19), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(KEYINPUT93), .B1(new_n480), .B2(G146), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT93), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n477), .A2(new_n479), .A3(new_n482), .A4(new_n187), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n475), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n465), .A2(new_n468), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n216), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n465), .A2(G131), .A3(new_n468), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AOI22_X1  g302(.A1(new_n471), .A2(new_n474), .B1(new_n484), .B2(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(G113), .B(G122), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n490), .B(new_n386), .ZN(new_n491));
  OAI21_X1  g305(.A(KEYINPUT94), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT95), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n493), .B1(new_n488), .B2(KEYINPUT17), .ZN(new_n494));
  INV_X1    g308(.A(new_n350), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT17), .ZN(new_n496));
  OR2_X1    g310(.A1(new_n487), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n486), .A2(KEYINPUT95), .A3(new_n496), .A4(new_n487), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n494), .A2(new_n495), .A3(new_n497), .A4(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n471), .A2(new_n474), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n499), .A2(new_n491), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n484), .A2(new_n488), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT94), .ZN(new_n504));
  INV_X1    g318(.A(new_n491), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n492), .A2(new_n501), .A3(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(G475), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n507), .A2(new_n508), .A3(new_n293), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(KEYINPUT20), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT20), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n507), .A2(new_n511), .A3(new_n508), .A4(new_n293), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n501), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n491), .B1(new_n499), .B2(new_n500), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n293), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(G475), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(KEYINPUT96), .B1(new_n190), .B2(new_n224), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT96), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n196), .A2(new_n521), .A3(G128), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n224), .A2(G143), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n520), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n524), .B(G134), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n248), .A2(KEYINPUT14), .A3(G122), .ZN(new_n526));
  XNOR2_X1  g340(.A(G116), .B(G122), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  OAI211_X1 g342(.A(G107), .B(new_n526), .C1(new_n528), .C2(KEYINPUT14), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n525), .B(new_n529), .C1(new_n409), .C2(new_n528), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT13), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n211), .B1(new_n523), .B2(new_n531), .ZN(new_n532));
  XOR2_X1   g346(.A(new_n524), .B(new_n532), .Z(new_n533));
  XNOR2_X1  g347(.A(new_n404), .B(new_n527), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  NOR3_X1   g350(.A1(new_n378), .A2(new_n320), .A3(G953), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n530), .A2(new_n535), .A3(new_n537), .ZN(new_n540));
  AOI21_X1  g354(.A(G902), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(G478), .ZN(new_n542));
  OAI22_X1  g356(.A1(new_n541), .A2(KEYINPUT97), .B1(KEYINPUT15), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n541), .B(KEYINPUT97), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n542), .A2(KEYINPUT15), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n267), .A2(G952), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n548), .B1(G234), .B2(G237), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  AOI211_X1 g364(.A(new_n293), .B(new_n267), .C1(G234), .C2(G237), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  XOR2_X1   g366(.A(KEYINPUT21), .B(G898), .Z(new_n553));
  OAI21_X1  g367(.A(new_n550), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n519), .A2(new_n547), .A3(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n432), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n408), .A2(KEYINPUT4), .ZN(new_n557));
  INV_X1    g371(.A(new_n431), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NOR3_X1   g373(.A1(new_n248), .A2(KEYINPUT5), .A3(G119), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n560), .B1(new_n250), .B2(KEYINPUT5), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n251), .B1(G113), .B2(new_n561), .ZN(new_n562));
  AND4_X1   g376(.A1(KEYINPUT85), .A2(new_n408), .A3(new_n412), .A4(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(KEYINPUT85), .B1(new_n416), .B2(new_n562), .ZN(new_n564));
  OAI22_X1  g378(.A1(new_n559), .A2(new_n253), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  XOR2_X1   g379(.A(G110), .B(G122), .Z(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n435), .A2(new_n263), .ZN(new_n568));
  INV_X1    g382(.A(new_n566), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n568), .B(new_n569), .C1(new_n564), .C2(new_n563), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n567), .A2(KEYINPUT6), .A3(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT6), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n565), .A2(new_n572), .A3(new_n566), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n275), .A2(G125), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(KEYINPUT86), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT86), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n275), .A2(new_n576), .A3(G125), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n414), .A2(new_n324), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n575), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(KEYINPUT87), .ZN(new_n580));
  AND2_X1   g394(.A1(new_n267), .A2(G224), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT87), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n575), .A2(new_n578), .A3(new_n582), .A4(new_n577), .ZN(new_n583));
  AND3_X1   g397(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n581), .B1(new_n580), .B2(new_n583), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n571), .A2(new_n573), .A3(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT7), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n581), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n575), .A2(new_n578), .A3(new_n577), .A4(new_n589), .ZN(new_n590));
  XOR2_X1   g404(.A(new_n590), .B(KEYINPUT89), .Z(new_n591));
  NOR2_X1   g405(.A1(new_n229), .A2(G125), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(KEYINPUT88), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n593), .A2(new_n577), .A3(new_n575), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n592), .A2(KEYINPUT88), .ZN(new_n595));
  OAI22_X1  g409(.A1(new_n594), .A2(new_n595), .B1(new_n588), .B2(new_n581), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n416), .B(new_n562), .ZN(new_n597));
  XOR2_X1   g411(.A(new_n566), .B(KEYINPUT8), .Z(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n591), .A2(new_n570), .A3(new_n596), .A4(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n587), .A2(new_n293), .A3(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(G210), .B1(G237), .B2(G902), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n587), .A2(new_n293), .A3(new_n602), .A4(new_n600), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(G214), .B1(G237), .B2(G902), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n555), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n319), .A2(new_n376), .A3(new_n462), .A4(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(new_n401), .ZN(G3));
  INV_X1    g425(.A(KEYINPUT98), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n539), .A2(new_n540), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT33), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n539), .A2(KEYINPUT33), .A3(new_n540), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n542), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n541), .A2(new_n542), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n542), .A2(new_n293), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n618), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n518), .A2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n607), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n625), .B1(new_n604), .B2(new_n605), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(KEYINPUT98), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n613), .A2(new_n554), .A3(new_n624), .A4(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(KEYINPUT99), .ZN(new_n629));
  AOI21_X1  g443(.A(KEYINPUT98), .B1(new_n606), .B2(new_n607), .ZN(new_n630));
  AOI211_X1 g444(.A(new_n612), .B(new_n625), .C1(new_n604), .C2(new_n605), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT99), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n632), .A2(new_n633), .A3(new_n554), .A4(new_n624), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n629), .A2(new_n634), .ZN(new_n635));
  AOI22_X1  g449(.A1(new_n311), .A2(new_n289), .B1(new_n265), .B2(new_n272), .ZN(new_n636));
  OAI21_X1  g450(.A(G472), .B1(new_n636), .B2(G902), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n294), .A2(new_n637), .ZN(new_n638));
  NOR3_X1   g452(.A1(new_n461), .A2(new_n375), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(new_n640), .B(KEYINPUT100), .Z(new_n641));
  XNOR2_X1  g455(.A(KEYINPUT34), .B(G104), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G6));
  XNOR2_X1  g457(.A(new_n512), .B(KEYINPUT101), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n547), .B1(new_n510), .B2(new_n644), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n632), .A2(new_n554), .A3(new_n517), .A4(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n639), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(KEYINPUT35), .B(G107), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G9));
  NOR2_X1   g464(.A1(new_n364), .A2(KEYINPUT36), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n362), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n373), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n371), .A2(new_n653), .ZN(new_n654));
  OAI211_X1 g468(.A(new_n379), .B(new_n654), .C1(new_n451), .C2(new_n460), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n656), .A2(new_n609), .A3(new_n294), .A4(new_n637), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT37), .B(G110), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G12));
  NAND2_X1  g473(.A1(new_n644), .A2(new_n510), .ZN(new_n660));
  INV_X1    g474(.A(new_n547), .ZN(new_n661));
  INV_X1    g475(.A(G900), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n549), .B1(new_n551), .B2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n517), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n660), .A2(new_n661), .A3(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n613), .A2(new_n627), .A3(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT102), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n613), .A2(new_n667), .A3(KEYINPUT102), .A4(new_n627), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n670), .A2(new_n319), .A3(new_n656), .A4(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G128), .ZN(G30));
  XNOR2_X1  g487(.A(new_n606), .B(KEYINPUT38), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n663), .B(KEYINPUT39), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n462), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n674), .B1(new_n677), .B2(KEYINPUT40), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  AOI21_X1  g493(.A(KEYINPUT32), .B1(new_n313), .B2(new_n292), .ZN(new_n680));
  NOR4_X1   g494(.A1(new_n636), .A2(new_n295), .A3(G472), .A4(G902), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n272), .B1(new_n274), .B2(new_n304), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n309), .A2(G472), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(G472), .A2(G902), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(new_n686), .B(KEYINPUT103), .Z(new_n687));
  AOI21_X1  g501(.A(new_n654), .B1(new_n682), .B2(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n625), .B1(new_n677), .B2(KEYINPUT40), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n519), .A2(new_n547), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n679), .A2(new_n688), .A3(new_n689), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(new_n190), .ZN(G45));
  NAND3_X1  g506(.A1(new_n518), .A2(new_n622), .A3(new_n664), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n319), .A2(new_n632), .A3(new_n656), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G146), .ZN(G48));
  INV_X1    g510(.A(KEYINPUT105), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT104), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n380), .B1(new_n456), .B2(new_n293), .ZN(new_n699));
  AOI211_X1 g513(.A(G469), .B(G902), .C1(new_n454), .C2(new_n455), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n698), .B1(new_n701), .B2(new_n379), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n441), .A2(new_n383), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n430), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n383), .B1(new_n445), .B2(new_n441), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n293), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(G469), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n707), .A2(new_n698), .A3(new_n379), .A4(new_n457), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n697), .B1(new_n702), .B2(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n707), .A2(new_n379), .A3(new_n457), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(KEYINPUT104), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n712), .A2(KEYINPUT105), .A3(new_n708), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n319), .A2(new_n710), .A3(new_n376), .A4(new_n713), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n714), .B1(new_n634), .B2(new_n629), .ZN(new_n715));
  XOR2_X1   g529(.A(KEYINPUT41), .B(G113), .Z(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(G15));
  NOR2_X1   g531(.A1(new_n714), .A2(new_n646), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(new_n248), .ZN(G18));
  NAND2_X1  g533(.A1(new_n712), .A2(new_n708), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n720), .A2(new_n630), .A3(new_n631), .ZN(new_n721));
  INV_X1    g535(.A(new_n555), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n721), .A2(new_n319), .A3(new_n722), .A4(new_n654), .ZN(new_n723));
  XOR2_X1   g537(.A(KEYINPUT106), .B(G119), .Z(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(G21));
  INV_X1    g539(.A(new_n713), .ZN(new_n726));
  AOI21_X1  g540(.A(KEYINPUT105), .B1(new_n712), .B2(new_n708), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n613), .A2(new_n627), .A3(new_n690), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT108), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n283), .B1(new_n305), .B2(KEYINPUT107), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n731), .B1(KEYINPUT107), .B2(new_n305), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n312), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n733), .A2(new_n292), .A3(new_n293), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n637), .ZN(new_n735));
  INV_X1    g549(.A(new_n554), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n375), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n728), .A2(new_n729), .A3(new_n730), .A4(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n710), .A2(new_n713), .A3(new_n737), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n632), .A2(new_n690), .ZN(new_n740));
  OAI21_X1  g554(.A(KEYINPUT108), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G122), .ZN(G24));
  NOR2_X1   g557(.A1(new_n702), .A2(new_n709), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n654), .A2(new_n637), .A3(new_n734), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(new_n693), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n744), .A2(new_n613), .A3(new_n627), .A4(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(KEYINPUT109), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT109), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n721), .A2(new_n749), .A3(new_n746), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G125), .ZN(G27));
  INV_X1    g566(.A(KEYINPUT110), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n443), .A2(G469), .A3(new_n446), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n457), .A2(new_n459), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n379), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n604), .A2(new_n607), .A3(new_n605), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n758), .A2(KEYINPUT42), .A3(new_n694), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n315), .A2(new_n376), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n753), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n760), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n756), .A2(new_n757), .A3(new_n693), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n762), .A2(new_n763), .A3(KEYINPUT110), .A4(KEYINPUT42), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n319), .A2(new_n376), .A3(new_n694), .A4(new_n758), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT42), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G131), .ZN(G33));
  NAND4_X1  g584(.A1(new_n319), .A2(new_n376), .A3(new_n667), .A4(new_n758), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G134), .ZN(G36));
  INV_X1    g586(.A(KEYINPUT45), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n449), .A2(new_n773), .A3(new_n450), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n774), .B(G469), .C1(new_n773), .C2(new_n447), .ZN(new_n775));
  AOI21_X1  g589(.A(KEYINPUT46), .B1(new_n775), .B2(new_n459), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n776), .A2(KEYINPUT111), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n775), .A2(KEYINPUT46), .A3(new_n459), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n776), .A2(KEYINPUT111), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n777), .A2(new_n457), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n379), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n781), .A2(new_n675), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n519), .A2(new_n622), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(KEYINPUT43), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n785), .A2(new_n638), .A3(new_n654), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT44), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n757), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n782), .B(new_n788), .C1(new_n787), .C2(new_n786), .ZN(new_n789));
  XNOR2_X1  g603(.A(KEYINPUT112), .B(G137), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n789), .B(new_n790), .ZN(G39));
  INV_X1    g605(.A(KEYINPUT47), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n792), .B1(new_n780), .B2(new_n379), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n780), .A2(new_n792), .A3(new_n379), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n794), .A2(new_n694), .A3(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n319), .ZN(new_n797));
  INV_X1    g611(.A(new_n757), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n796), .A2(new_n797), .A3(new_n375), .A4(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G140), .ZN(G42));
  INV_X1    g614(.A(new_n701), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n783), .B1(new_n801), .B2(KEYINPUT49), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n802), .A2(new_n376), .A3(new_n379), .A4(new_n607), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT113), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n674), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n803), .A2(new_n804), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n682), .A2(new_n687), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT49), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n808), .B1(new_n809), .B2(new_n701), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n805), .A2(new_n806), .A3(new_n807), .A4(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT118), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n801), .A2(new_n379), .ZN(new_n813));
  AOI22_X1  g627(.A1(new_n794), .A2(new_n795), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n814), .B1(new_n812), .B2(new_n813), .ZN(new_n815));
  NOR4_X1   g629(.A1(new_n784), .A2(new_n375), .A3(new_n550), .A4(new_n735), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(new_n798), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n816), .A2(new_n625), .A3(new_n806), .A4(new_n744), .ZN(new_n820));
  NOR2_X1   g634(.A1(KEYINPUT119), .A2(KEYINPUT50), .ZN(new_n821));
  AND2_X1   g635(.A1(KEYINPUT119), .A2(KEYINPUT50), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n820), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n823), .B1(new_n820), .B2(new_n821), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n824), .B1(KEYINPUT120), .B2(KEYINPUT51), .ZN(new_n825));
  OR2_X1    g639(.A1(new_n824), .A2(KEYINPUT120), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n720), .A2(new_n757), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n785), .A2(new_n549), .A3(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n828), .A2(new_n745), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n827), .A2(new_n376), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n830), .A2(new_n550), .A3(new_n808), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n518), .A2(new_n622), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n829), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n819), .A2(new_n825), .A3(new_n826), .A4(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n813), .B1(new_n794), .B2(new_n795), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n824), .B(new_n833), .C1(new_n835), .C2(new_n817), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT51), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n548), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n816), .A2(new_n744), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(new_n632), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n751), .A2(new_n672), .A3(new_n695), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT116), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n756), .A2(new_n663), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n688), .A2(new_n729), .A3(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n841), .A2(new_n842), .A3(KEYINPUT52), .A4(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n751), .A2(new_n672), .A3(new_n695), .A4(new_n844), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT52), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(KEYINPUT116), .B1(new_n846), .B2(new_n847), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n845), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n623), .B1(new_n547), .B2(new_n518), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n639), .A2(new_n626), .A3(new_n554), .A4(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n853), .A2(new_n610), .A3(new_n657), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n660), .A2(new_n666), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n604), .A2(new_n547), .A3(new_n607), .A4(new_n605), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT114), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n665), .B1(new_n644), .B2(new_n510), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT114), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n798), .A2(new_n858), .A3(new_n859), .A4(new_n547), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n319), .A2(new_n656), .A3(new_n857), .A4(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n746), .A2(new_n758), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n771), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(KEYINPUT115), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT115), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n771), .A2(new_n861), .A3(new_n865), .A4(new_n862), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n854), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n723), .B1(new_n646), .B2(new_n714), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n868), .A2(new_n715), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n867), .A2(new_n742), .A3(new_n769), .A4(new_n869), .ZN(new_n870));
  OR3_X1    g684(.A1(new_n851), .A2(KEYINPUT53), .A3(new_n870), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n846), .B(KEYINPUT52), .ZN(new_n872));
  OAI21_X1  g686(.A(KEYINPUT53), .B1(new_n872), .B2(new_n870), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n871), .A2(KEYINPUT54), .A3(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT53), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n875), .B1(new_n872), .B2(new_n870), .ZN(new_n876));
  INV_X1    g690(.A(new_n868), .ZN(new_n877));
  INV_X1    g691(.A(new_n715), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n877), .A2(new_n878), .A3(new_n742), .A4(new_n769), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(KEYINPUT117), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT117), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n869), .A2(new_n881), .A3(new_n742), .A4(new_n769), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n880), .A2(KEYINPUT53), .A3(new_n867), .A4(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n876), .B1(new_n851), .B2(new_n883), .ZN(new_n884));
  OR2_X1    g698(.A1(new_n884), .A2(KEYINPUT54), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n838), .A2(new_n840), .A3(new_n874), .A4(new_n885), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n831), .A2(new_n624), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n828), .A2(new_n760), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT48), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n886), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(G952), .A2(G953), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n811), .B1(new_n890), .B2(new_n891), .ZN(G75));
  AND2_X1   g706(.A1(new_n882), .A2(KEYINPUT53), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n864), .A2(new_n866), .ZN(new_n894));
  INV_X1    g708(.A(new_n854), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n896), .B1(KEYINPUT117), .B2(new_n879), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n893), .A2(new_n897), .A3(new_n850), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n293), .B1(new_n898), .B2(new_n876), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT56), .B1(new_n899), .B2(G210), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n571), .A2(new_n573), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(new_n586), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT55), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n900), .B(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n267), .A2(G952), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n904), .A2(new_n905), .ZN(G51));
  NAND2_X1  g720(.A1(new_n884), .A2(KEYINPUT54), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n885), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n459), .A2(KEYINPUT57), .ZN(new_n909));
  OR2_X1    g723(.A1(new_n459), .A2(KEYINPUT57), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(new_n456), .ZN(new_n912));
  INV_X1    g726(.A(new_n899), .ZN(new_n913));
  OR2_X1    g727(.A1(new_n913), .A2(new_n775), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n905), .B1(new_n912), .B2(new_n914), .ZN(G54));
  NAND3_X1  g729(.A1(new_n899), .A2(KEYINPUT58), .A3(G475), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(new_n507), .Z(new_n917));
  NOR2_X1   g731(.A1(new_n917), .A2(new_n905), .ZN(G60));
  INV_X1    g732(.A(new_n905), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n621), .B(KEYINPUT59), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n920), .B1(new_n874), .B2(new_n885), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n616), .A2(new_n617), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n919), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n920), .B1(new_n907), .B2(new_n885), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n924), .B1(new_n925), .B2(new_n923), .ZN(G63));
  NAND2_X1  g740(.A1(G217), .A2(G902), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT60), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n928), .B1(new_n898), .B2(new_n876), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n929), .A2(KEYINPUT124), .A3(new_n365), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT61), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n928), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n884), .A2(new_n652), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(KEYINPUT122), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT122), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n929), .A2(new_n936), .A3(new_n652), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(KEYINPUT124), .B1(new_n929), .B2(new_n365), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n932), .A2(new_n938), .A3(new_n919), .A4(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n919), .B1(new_n929), .B2(new_n365), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n941), .B1(new_n935), .B2(new_n937), .ZN(new_n942));
  XNOR2_X1  g756(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n942), .A2(KEYINPUT123), .A3(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT123), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n884), .A2(new_n933), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n905), .B1(new_n946), .B2(new_n372), .ZN(new_n947));
  AND4_X1   g761(.A1(new_n936), .A2(new_n884), .A3(new_n652), .A4(new_n933), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n936), .B1(new_n929), .B2(new_n652), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n943), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n945), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n940), .B1(new_n944), .B2(new_n952), .ZN(G66));
  AOI21_X1  g767(.A(new_n267), .B1(new_n553), .B2(G224), .ZN(new_n954));
  INV_X1    g768(.A(new_n742), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n955), .A2(new_n715), .A3(new_n868), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(new_n895), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n954), .B1(new_n957), .B2(new_n267), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n901), .B1(G898), .B2(new_n267), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n958), .B(new_n959), .Z(G69));
  NAND2_X1  g774(.A1(G227), .A2(G900), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n267), .A2(G900), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n780), .A2(new_n379), .A3(new_n676), .A4(new_n729), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n963), .A2(new_n760), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT125), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n964), .B(new_n965), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n841), .A2(new_n769), .A3(new_n771), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n799), .A2(new_n966), .A3(new_n789), .A4(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n962), .B1(new_n968), .B2(new_n267), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT126), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n281), .B(new_n480), .Z(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  OAI211_X1 g787(.A(G953), .B(new_n961), .C1(new_n971), .C2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n968), .A2(new_n267), .ZN(new_n975));
  INV_X1    g789(.A(new_n962), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n970), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  AOI211_X1 g791(.A(KEYINPUT126), .B(new_n962), .C1(new_n968), .C2(new_n267), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n972), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n961), .A2(G953), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n841), .A2(new_n691), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(KEYINPUT62), .Z(new_n982));
  NOR2_X1   g796(.A1(new_n677), .A2(new_n757), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n983), .A2(new_n319), .A3(new_n376), .A4(new_n852), .ZN(new_n984));
  AND4_X1   g798(.A1(new_n789), .A2(new_n982), .A3(new_n799), .A4(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n973), .B1(new_n985), .B2(G953), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n979), .A2(new_n980), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n974), .A2(new_n987), .ZN(G72));
  NOR2_X1   g802(.A1(new_n282), .A2(new_n272), .ZN(new_n989));
  INV_X1    g803(.A(new_n957), .ZN(new_n990));
  AND2_X1   g804(.A1(new_n985), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n685), .B(KEYINPUT63), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n989), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n282), .A2(new_n272), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n994), .B(KEYINPUT127), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n968), .A2(new_n957), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n995), .B1(new_n996), .B2(new_n992), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n993), .A2(new_n919), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n871), .A2(new_n873), .ZN(new_n999));
  INV_X1    g813(.A(new_n994), .ZN(new_n1000));
  NOR4_X1   g814(.A1(new_n999), .A2(new_n992), .A3(new_n989), .A4(new_n1000), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n998), .A2(new_n1001), .ZN(G57));
endmodule


