//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 0 1 1 1 1 1 0 1 1 0 1 0 1 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 0 0 1 1 1 1 1 1 0 1 0 0 1 0 1 1 0 0 0 0 1 1 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n742, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n831, new_n832, new_n833, new_n835,
    new_n836, new_n837, new_n838, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975, new_n976, new_n977;
  INV_X1    g000(.A(KEYINPUT86), .ZN(new_n202));
  NAND2_X1  g001(.A1(G228gat), .A2(G233gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G141gat), .B(G148gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(KEYINPUT75), .B(KEYINPUT2), .ZN(new_n208));
  OAI211_X1 g007(.A(new_n204), .B(new_n206), .C1(new_n207), .C2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G141gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n210), .A2(G148gat), .ZN(new_n211));
  XNOR2_X1  g010(.A(KEYINPUT76), .B(G141gat), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n211), .B1(new_n212), .B2(G148gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n204), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT2), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n214), .B1(new_n215), .B2(new_n205), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n209), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(G211gat), .B(G218gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(G211gat), .A2(G218gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT22), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G197gat), .B(G204gat), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n219), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT78), .ZN(new_n225));
  AOI21_X1  g024(.A(KEYINPUT29), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NOR2_X1   g025(.A1(G197gat), .A2(G204gat), .ZN(new_n227));
  AND2_X1   g026(.A1(G197gat), .A2(G204gat), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n222), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  XOR2_X1   g028(.A(G211gat), .B(G218gat), .Z(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n219), .A2(new_n223), .A3(new_n222), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n226), .B1(new_n233), .B2(new_n225), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n218), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n209), .B(new_n235), .C1(new_n213), .C2(new_n216), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT29), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n233), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n203), .B1(new_n236), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n237), .A2(new_n238), .ZN(new_n241));
  INV_X1    g040(.A(new_n233), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n203), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(KEYINPUT29), .B1(new_n231), .B2(new_n232), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT79), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT3), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n229), .A2(new_n230), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n238), .B1(new_n247), .B2(new_n224), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(KEYINPUT79), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n218), .B1(new_n246), .B2(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n243), .B1(new_n250), .B2(KEYINPUT80), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT80), .ZN(new_n252));
  AOI211_X1 g051(.A(new_n252), .B(new_n218), .C1(new_n246), .C2(new_n249), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n240), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(G22gat), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT81), .ZN(new_n256));
  INV_X1    g055(.A(G22gat), .ZN(new_n257));
  OAI211_X1 g056(.A(new_n240), .B(new_n257), .C1(new_n251), .C2(new_n253), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n255), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT82), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT82), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n255), .A2(new_n256), .A3(new_n261), .A4(new_n258), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n255), .A2(new_n258), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(KEYINPUT81), .ZN(new_n265));
  XNOR2_X1  g064(.A(G78gat), .B(G106gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(KEYINPUT31), .B(G50gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n266), .B(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n263), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n268), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n271), .B1(new_n264), .B2(KEYINPUT81), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n272), .A2(new_n260), .A3(new_n262), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(G71gat), .B(G99gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n275), .B(KEYINPUT71), .ZN(new_n276));
  INV_X1    g075(.A(G15gat), .ZN(new_n277));
  OR2_X1    g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n277), .ZN(new_n279));
  AND3_X1   g078(.A1(new_n278), .A2(G43gat), .A3(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(G43gat), .B1(new_n278), .B2(new_n279), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(G227gat), .ZN(new_n283));
  INV_X1    g082(.A(G233gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G113gat), .B(G120gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT69), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT1), .ZN(new_n289));
  XNOR2_X1  g088(.A(G127gat), .B(G134gat), .ZN(new_n290));
  INV_X1    g089(.A(G120gat), .ZN(new_n291));
  OR3_X1    g090(.A1(new_n291), .A2(KEYINPUT69), .A3(G113gat), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n288), .A2(new_n289), .A3(new_n290), .A4(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n290), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n294), .B1(KEYINPUT1), .B2(new_n287), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT25), .ZN(new_n297));
  NOR2_X1   g096(.A1(G169gat), .A2(G176gat), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT23), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(G169gat), .ZN(new_n301));
  INV_X1    g100(.A(G176gat), .ZN(new_n302));
  OAI21_X1  g101(.A(KEYINPUT64), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT64), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n304), .A2(G169gat), .A3(G176gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n300), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(G183gat), .A2(G190gat), .ZN(new_n308));
  OR2_X1    g107(.A1(new_n308), .A2(KEYINPUT65), .ZN(new_n309));
  AOI21_X1  g108(.A(KEYINPUT24), .B1(new_n308), .B2(KEYINPUT65), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OR2_X1    g110(.A1(G183gat), .A2(G190gat), .ZN(new_n312));
  NAND3_X1  g111(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT66), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n307), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n312), .A2(new_n313), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n317), .B1(new_n309), .B2(new_n310), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT66), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n297), .B1(new_n316), .B2(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n321));
  OR2_X1    g120(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n322), .A2(new_n297), .A3(new_n306), .A4(new_n300), .ZN(new_n323));
  OAI21_X1  g122(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n324), .B(KEYINPUT68), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT26), .ZN(new_n326));
  AOI22_X1  g125(.A1(new_n303), .A2(new_n305), .B1(new_n326), .B2(new_n298), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(KEYINPUT27), .B(G183gat), .ZN(new_n330));
  INV_X1    g129(.A(G190gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AND2_X1   g131(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NOR2_X1   g133(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n336), .A2(new_n330), .A3(new_n331), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n334), .A2(new_n308), .A3(new_n337), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n323), .B1(new_n329), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n296), .B1(new_n320), .B2(new_n339), .ZN(new_n340));
  AND3_X1   g139(.A1(new_n334), .A2(new_n308), .A3(new_n337), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n307), .A2(KEYINPUT25), .ZN(new_n342));
  AOI22_X1  g141(.A1(new_n341), .A2(new_n328), .B1(new_n342), .B2(new_n322), .ZN(new_n343));
  INV_X1    g142(.A(new_n319), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n306), .B(new_n300), .C1(new_n318), .C2(KEYINPUT66), .ZN(new_n345));
  OAI21_X1  g144(.A(KEYINPUT25), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n296), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n343), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n286), .B1(new_n340), .B2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(KEYINPUT70), .B(KEYINPUT33), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n282), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT32), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n340), .A2(new_n348), .ZN(new_n356));
  AOI221_X4 g155(.A(new_n353), .B1(new_n282), .B2(new_n351), .C1(new_n356), .C2(new_n285), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n340), .A2(new_n348), .A3(new_n286), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT34), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n359), .B(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT72), .B1(new_n358), .B2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n359), .B(KEYINPUT34), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n363), .B1(new_n355), .B2(new_n357), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n356), .A2(new_n285), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT32), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n350), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n366), .A2(new_n367), .A3(new_n282), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n354), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n368), .A2(new_n361), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n364), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n362), .B1(KEYINPUT72), .B2(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(G8gat), .B(G36gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(G64gat), .B(G92gat), .ZN(new_n374));
  XOR2_X1   g173(.A(new_n373), .B(new_n374), .Z(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(G226gat), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n377), .A2(new_n284), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT73), .ZN(new_n379));
  NOR3_X1   g178(.A1(new_n320), .A2(new_n339), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT73), .B1(new_n343), .B2(new_n346), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n378), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n378), .A2(KEYINPUT29), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n383), .B1(new_n320), .B2(new_n339), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n242), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n379), .B1(new_n320), .B2(new_n339), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n343), .A2(new_n346), .A3(KEYINPUT73), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n386), .A2(new_n387), .A3(new_n383), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n343), .A2(new_n346), .A3(new_n378), .ZN(new_n389));
  AND3_X1   g188(.A1(new_n388), .A2(new_n242), .A3(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n376), .B1(new_n385), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT74), .ZN(new_n392));
  INV_X1    g191(.A(new_n378), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n393), .B1(new_n386), .B2(new_n387), .ZN(new_n394));
  INV_X1    g193(.A(new_n384), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n233), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n388), .A2(new_n242), .A3(new_n389), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n375), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT74), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n396), .A2(new_n397), .A3(new_n375), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(KEYINPUT30), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT30), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n396), .A2(new_n397), .A3(new_n403), .A4(new_n375), .ZN(new_n404));
  AOI22_X1  g203(.A1(new_n392), .A2(new_n400), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT5), .ZN(new_n406));
  OR2_X1    g205(.A1(new_n213), .A2(new_n216), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n407), .A2(new_n209), .A3(new_n295), .A4(new_n293), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n296), .A2(new_n217), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(G225gat), .A2(G233gat), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n406), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n217), .A2(KEYINPUT3), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n415), .A2(new_n237), .A3(new_n296), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n347), .A2(new_n218), .A3(KEYINPUT4), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT4), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n418), .B1(new_n296), .B2(new_n217), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n416), .A2(new_n417), .A3(new_n411), .A4(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n414), .A2(new_n420), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n416), .A2(new_n417), .A3(new_n419), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n422), .A2(KEYINPUT5), .A3(new_n411), .ZN(new_n423));
  XOR2_X1   g222(.A(G1gat), .B(G29gat), .Z(new_n424));
  XNOR2_X1  g223(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n424), .B(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(G57gat), .B(G85gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n426), .B(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n421), .A2(new_n423), .A3(KEYINPUT6), .A4(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT84), .ZN(new_n431));
  AND2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n413), .B1(new_n422), .B2(new_n411), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n420), .A2(new_n406), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n428), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT6), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n421), .A2(new_n423), .A3(new_n429), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n430), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n432), .B1(new_n439), .B2(KEYINPUT84), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n440), .A2(KEYINPUT35), .ZN(new_n441));
  AND4_X1   g240(.A1(new_n274), .A2(new_n372), .A3(new_n405), .A4(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n371), .ZN(new_n443));
  AND3_X1   g242(.A1(new_n272), .A2(new_n260), .A3(new_n262), .ZN(new_n444));
  AOI22_X1  g243(.A1(new_n260), .A2(new_n262), .B1(new_n265), .B2(new_n268), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT85), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n402), .A2(new_n404), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n398), .A2(new_n399), .ZN(new_n450));
  AOI211_X1 g249(.A(KEYINPUT74), .B(new_n375), .C1(new_n396), .C2(new_n397), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n439), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n274), .A2(KEYINPUT85), .A3(new_n443), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n448), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n442), .B1(new_n456), .B2(KEYINPUT35), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n416), .A2(new_n417), .A3(new_n419), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n412), .ZN(new_n459));
  OR2_X1    g258(.A1(new_n459), .A2(KEYINPUT39), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n459), .B(KEYINPUT39), .C1(new_n412), .C2(new_n410), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(new_n461), .A3(new_n428), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT40), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n460), .A2(new_n461), .A3(KEYINPUT40), .A4(new_n428), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n464), .A2(new_n437), .A3(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT83), .B1(new_n405), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT37), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n375), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n398), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n468), .B1(new_n396), .B2(new_n397), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT38), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n242), .B1(new_n394), .B2(new_n395), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n388), .A2(new_n233), .A3(new_n389), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n473), .A2(KEYINPUT37), .A3(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT38), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n475), .B(new_n476), .C1(new_n398), .C2(new_n469), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n440), .A2(new_n472), .A3(new_n477), .A4(new_n401), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT83), .ZN(new_n479));
  INV_X1    g278(.A(new_n466), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n452), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  AND4_X1   g280(.A1(new_n274), .A2(new_n467), .A3(new_n478), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n371), .A2(KEYINPUT72), .ZN(new_n483));
  INV_X1    g282(.A(new_n362), .ZN(new_n484));
  AOI21_X1  g283(.A(KEYINPUT36), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n443), .A2(KEYINPUT36), .ZN(new_n486));
  OAI22_X1  g285(.A1(new_n485), .A2(new_n486), .B1(new_n454), .B2(new_n274), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n482), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n457), .A2(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(G15gat), .B(G22gat), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT16), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n490), .B1(new_n491), .B2(G1gat), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n492), .B1(G1gat), .B2(new_n490), .ZN(new_n493));
  XOR2_X1   g292(.A(new_n493), .B(G8gat), .Z(new_n494));
  XOR2_X1   g293(.A(G43gat), .B(G50gat), .Z(new_n495));
  INV_X1    g294(.A(G36gat), .ZN(new_n496));
  AND2_X1   g295(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n497));
  NOR2_X1   g296(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(G29gat), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n500), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n495), .B1(new_n502), .B2(KEYINPUT15), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n503), .B1(KEYINPUT15), .B2(new_n502), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n502), .A2(KEYINPUT15), .A3(new_n495), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AND2_X1   g305(.A1(new_n506), .A2(KEYINPUT17), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n506), .A2(KEYINPUT17), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n494), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(G229gat), .A2(G233gat), .ZN(new_n510));
  INV_X1    g309(.A(new_n506), .ZN(new_n511));
  OR2_X1    g310(.A1(new_n511), .A2(new_n494), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n509), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT18), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n509), .A2(KEYINPUT18), .A3(new_n510), .A4(new_n512), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n511), .A2(new_n494), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n512), .A2(new_n517), .ZN(new_n518));
  XOR2_X1   g317(.A(new_n510), .B(KEYINPUT13), .Z(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n515), .A2(new_n516), .A3(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(G113gat), .B(G141gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(G197gat), .ZN(new_n523));
  XOR2_X1   g322(.A(KEYINPUT11), .B(G169gat), .Z(new_n524));
  XNOR2_X1  g323(.A(new_n523), .B(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(KEYINPUT12), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n521), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n515), .A2(new_n526), .A3(new_n516), .A4(new_n520), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n202), .B1(new_n489), .B2(new_n531), .ZN(new_n532));
  OAI211_X1 g331(.A(KEYINPUT86), .B(new_n530), .C1(new_n457), .C2(new_n488), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT87), .ZN(new_n535));
  AOI22_X1  g334(.A1(new_n535), .A2(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n536), .B1(G71gat), .B2(G78gat), .ZN(new_n537));
  AOI21_X1  g336(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n538));
  AND2_X1   g337(.A1(G57gat), .A2(G64gat), .ZN(new_n539));
  NOR2_X1   g338(.A1(G57gat), .A2(G64gat), .ZN(new_n540));
  NOR3_X1   g339(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n537), .B(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT21), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(new_n544), .B(KEYINPUT88), .Z(new_n545));
  XOR2_X1   g344(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G183gat), .B(G211gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n494), .B1(new_n543), .B2(new_n542), .ZN(new_n550));
  XNOR2_X1  g349(.A(G127gat), .B(G155gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(G231gat), .A2(G233gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n550), .B(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n549), .B(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G190gat), .B(G218gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(G134gat), .B(G162gat), .ZN(new_n558));
  XOR2_X1   g357(.A(new_n557), .B(new_n558), .Z(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(G85gat), .A2(G92gat), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT90), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(KEYINPUT90), .A2(G85gat), .A3(G92gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT89), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT7), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n563), .A2(new_n566), .A3(KEYINPUT7), .A4(new_n564), .ZN(new_n569));
  NAND2_X1  g368(.A1(G99gat), .A2(G106gat), .ZN(new_n570));
  INV_X1    g369(.A(G85gat), .ZN(new_n571));
  INV_X1    g370(.A(G92gat), .ZN(new_n572));
  AOI22_X1  g371(.A1(KEYINPUT8), .A2(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n568), .A2(new_n569), .A3(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G99gat), .B(G106gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(KEYINPUT91), .ZN(new_n576));
  OR2_X1    g375(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n574), .A2(new_n576), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(new_n506), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT92), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT41), .ZN(new_n582));
  INV_X1    g381(.A(G232gat), .ZN(new_n583));
  NOR3_X1   g382(.A1(new_n582), .A2(new_n583), .A3(new_n284), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n580), .A2(new_n581), .A3(new_n585), .ZN(new_n586));
  AOI22_X1  g385(.A1(new_n577), .A2(new_n578), .B1(new_n504), .B2(new_n505), .ZN(new_n587));
  OAI21_X1  g386(.A(KEYINPUT92), .B1(new_n587), .B2(new_n584), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  OAI211_X1 g388(.A(new_n577), .B(new_n578), .C1(new_n507), .C2(new_n508), .ZN(new_n590));
  AOI21_X1  g389(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n589), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n592), .B1(new_n589), .B2(new_n590), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n560), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n595), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n597), .A2(new_n593), .A3(new_n559), .ZN(new_n598));
  AND2_X1   g397(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n556), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(G230gat), .A2(G233gat), .ZN(new_n602));
  INV_X1    g401(.A(new_n542), .ZN(new_n603));
  AND2_X1   g402(.A1(new_n574), .A2(new_n576), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n574), .A2(new_n576), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n577), .A2(new_n542), .A3(new_n578), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT10), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT93), .ZN(new_n610));
  AND2_X1   g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n606), .A2(new_n607), .A3(KEYINPUT93), .A4(new_n608), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n579), .A2(KEYINPUT10), .A3(new_n603), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n602), .B1(new_n611), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n606), .A2(new_n607), .ZN(new_n616));
  INV_X1    g415(.A(new_n602), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G120gat), .B(G148gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(G176gat), .B(G204gat), .ZN(new_n621));
  XOR2_X1   g420(.A(new_n620), .B(new_n621), .Z(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n615), .A2(new_n618), .A3(new_n622), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT94), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n624), .A2(KEYINPUT94), .A3(new_n625), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n601), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n534), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n633), .A2(new_n439), .ZN(new_n634));
  XNOR2_X1  g433(.A(KEYINPUT95), .B(G1gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(G1324gat));
  INV_X1    g435(.A(KEYINPUT42), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n633), .A2(new_n405), .ZN(new_n638));
  XOR2_X1   g437(.A(KEYINPUT16), .B(G8gat), .Z(new_n639));
  AOI21_X1  g438(.A(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(G8gat), .B1(new_n633), .B2(new_n405), .ZN(new_n641));
  NOR2_X1   g440(.A1(KEYINPUT96), .A2(KEYINPUT42), .ZN(new_n642));
  MUX2_X1   g441(.A(KEYINPUT96), .B(new_n642), .S(new_n639), .Z(new_n643));
  AOI22_X1  g442(.A1(new_n640), .A2(new_n641), .B1(new_n638), .B2(new_n643), .ZN(G1325gat));
  INV_X1    g443(.A(new_n485), .ZN(new_n645));
  INV_X1    g444(.A(new_n486), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NOR3_X1   g446(.A1(new_n633), .A2(new_n277), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n483), .A2(new_n484), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n277), .B1(new_n633), .B2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT97), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  OAI211_X1 g451(.A(KEYINPUT97), .B(new_n277), .C1(new_n633), .C2(new_n649), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n648), .B1(new_n652), .B2(new_n653), .ZN(G1326gat));
  NOR2_X1   g453(.A1(new_n633), .A2(new_n274), .ZN(new_n655));
  XOR2_X1   g454(.A(KEYINPUT43), .B(G22gat), .Z(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(G1327gat));
  NAND3_X1  g456(.A1(new_n555), .A2(new_n630), .A3(new_n599), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT98), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n660), .B1(new_n532), .B2(new_n533), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n661), .A2(new_n500), .A3(new_n453), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT45), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n662), .A2(new_n663), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n599), .B1(new_n457), .B2(new_n488), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OAI211_X1 g467(.A(KEYINPUT44), .B(new_n599), .C1(new_n457), .C2(new_n488), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n631), .A2(new_n556), .A3(new_n531), .ZN(new_n671));
  AND3_X1   g470(.A1(new_n670), .A2(new_n453), .A3(new_n671), .ZN(new_n672));
  OAI211_X1 g471(.A(new_n664), .B(new_n665), .C1(new_n500), .C2(new_n672), .ZN(G1328gat));
  INV_X1    g472(.A(new_n661), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n452), .A2(new_n496), .ZN(new_n675));
  OAI21_X1  g474(.A(KEYINPUT46), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  OR3_X1    g475(.A1(new_n674), .A2(KEYINPUT46), .A3(new_n675), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n670), .A2(new_n452), .A3(new_n671), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(KEYINPUT99), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(G36gat), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n678), .A2(KEYINPUT99), .ZN(new_n681));
  OAI211_X1 g480(.A(new_n676), .B(new_n677), .C1(new_n680), .C2(new_n681), .ZN(G1329gat));
  INV_X1    g481(.A(new_n647), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n683), .A2(G43gat), .ZN(new_n684));
  AND3_X1   g483(.A1(new_n670), .A2(new_n671), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(G43gat), .B1(new_n661), .B2(new_n372), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT47), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(KEYINPUT47), .B1(new_n685), .B2(new_n686), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(G1330gat));
  NOR2_X1   g490(.A1(new_n274), .A2(G50gat), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT101), .ZN(new_n693));
  INV_X1    g492(.A(new_n274), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n694), .B1(new_n453), .B2(new_n452), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n478), .A2(new_n274), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n467), .A2(new_n481), .ZN(new_n697));
  OAI211_X1 g496(.A(new_n647), .B(new_n695), .C1(new_n696), .C2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT35), .ZN(new_n699));
  AOI21_X1  g498(.A(KEYINPUT85), .B1(new_n274), .B2(new_n443), .ZN(new_n700));
  AOI211_X1 g499(.A(new_n447), .B(new_n371), .C1(new_n270), .C2(new_n273), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n699), .B1(new_n702), .B2(new_n454), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n698), .B1(new_n703), .B2(new_n442), .ZN(new_n704));
  AOI21_X1  g503(.A(KEYINPUT86), .B1(new_n704), .B2(new_n530), .ZN(new_n705));
  INV_X1    g504(.A(new_n533), .ZN(new_n706));
  OAI211_X1 g505(.A(new_n659), .B(new_n693), .C1(new_n705), .C2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT102), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n668), .A2(new_n694), .A3(new_n669), .A4(new_n671), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n710), .A2(KEYINPUT100), .A3(G50gat), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n661), .A2(KEYINPUT102), .A3(new_n693), .ZN(new_n712));
  AND3_X1   g511(.A1(new_n709), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT48), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT103), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n707), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n661), .A2(KEYINPUT103), .A3(new_n693), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n714), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n710), .A2(G50gat), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT100), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n719), .B1(new_n720), .B2(KEYINPUT48), .ZN(new_n721));
  OAI22_X1  g520(.A1(new_n713), .A2(KEYINPUT48), .B1(new_n718), .B2(new_n721), .ZN(G1331gat));
  NOR3_X1   g521(.A1(new_n489), .A2(new_n530), .A3(new_n601), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(new_n631), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n724), .A2(new_n439), .ZN(new_n725));
  XOR2_X1   g524(.A(KEYINPUT104), .B(G57gat), .Z(new_n726));
  XNOR2_X1  g525(.A(new_n725), .B(new_n726), .ZN(G1332gat));
  NOR2_X1   g526(.A1(new_n630), .A2(new_n405), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n729), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n723), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT105), .ZN(new_n732));
  OR2_X1    g531(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n732), .B(new_n733), .ZN(G1333gat));
  OR3_X1    g533(.A1(new_n724), .A2(G71gat), .A3(new_n649), .ZN(new_n735));
  OAI21_X1  g534(.A(G71gat), .B1(new_n724), .B2(new_n647), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT50), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n735), .A2(KEYINPUT50), .A3(new_n736), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(G1334gat));
  NOR2_X1   g540(.A1(new_n724), .A2(new_n274), .ZN(new_n742));
  XOR2_X1   g541(.A(new_n742), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g542(.A1(new_n556), .A2(new_n530), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n745), .A2(new_n630), .ZN(new_n746));
  AND3_X1   g545(.A1(new_n670), .A2(new_n453), .A3(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT51), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n748), .B1(new_n666), .B2(new_n745), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n704), .A2(KEYINPUT51), .A3(new_n599), .A4(new_n744), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT106), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n752), .B1(new_n751), .B2(new_n749), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n631), .A2(new_n571), .A3(new_n453), .ZN(new_n754));
  OAI22_X1  g553(.A1(new_n747), .A2(new_n571), .B1(new_n753), .B2(new_n754), .ZN(G1336gat));
  NAND4_X1  g554(.A1(new_n668), .A2(new_n452), .A3(new_n669), .A4(new_n746), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(G92gat), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n749), .A2(new_n750), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n729), .A2(G92gat), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n757), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(KEYINPUT52), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT107), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n756), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n756), .A2(new_n763), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n764), .A2(new_n765), .A3(new_n572), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n767), .B1(new_n753), .B2(new_n760), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n762), .B1(new_n766), .B2(new_n768), .ZN(G1337gat));
  NAND3_X1  g568(.A1(new_n670), .A2(new_n683), .A3(new_n746), .ZN(new_n770));
  XOR2_X1   g569(.A(KEYINPUT108), .B(G99gat), .Z(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  OR3_X1    g571(.A1(new_n649), .A2(new_n630), .A3(new_n771), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n772), .B1(new_n753), .B2(new_n773), .ZN(G1338gat));
  NAND4_X1  g573(.A1(new_n668), .A2(new_n694), .A3(new_n669), .A4(new_n746), .ZN(new_n775));
  AOI21_X1  g574(.A(KEYINPUT53), .B1(new_n775), .B2(G106gat), .ZN(new_n776));
  OR3_X1    g575(.A1(new_n274), .A2(new_n630), .A3(G106gat), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n776), .B1(new_n753), .B2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT109), .ZN(new_n779));
  AND3_X1   g578(.A1(new_n775), .A2(new_n779), .A3(G106gat), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n779), .B1(new_n775), .B2(G106gat), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n777), .B1(new_n749), .B2(new_n750), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT53), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n778), .B1(new_n783), .B2(new_n784), .ZN(G1339gat));
  AND2_X1   g584(.A1(new_n612), .A2(new_n613), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n609), .A2(new_n610), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n617), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT54), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n622), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n786), .A2(new_n617), .A3(new_n787), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n791), .A2(new_n615), .A3(KEYINPUT54), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n790), .A2(KEYINPUT55), .A3(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT110), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n790), .A2(KEYINPUT110), .A3(new_n792), .A4(KEYINPUT55), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n795), .A2(new_n625), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n790), .A2(new_n792), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT55), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n518), .A2(new_n519), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n510), .B1(new_n509), .B2(new_n512), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n525), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n529), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n599), .A2(new_n800), .A3(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(KEYINPUT111), .B1(new_n797), .B2(new_n805), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n596), .A2(new_n598), .A3(new_n529), .A4(new_n803), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT55), .B1(new_n790), .B2(new_n792), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n796), .A2(new_n625), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT111), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n809), .A2(new_n810), .A3(new_n811), .A4(new_n795), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n806), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n810), .A2(new_n530), .A3(new_n800), .A4(new_n795), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n628), .A2(new_n629), .A3(new_n804), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n599), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n555), .B1(new_n813), .B2(new_n816), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n556), .A2(new_n531), .A3(new_n630), .A4(new_n600), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n439), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n702), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n820), .A2(new_n452), .ZN(new_n821));
  AOI21_X1  g620(.A(G113gat), .B1(new_n821), .B2(new_n530), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n694), .B1(new_n817), .B2(new_n818), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n452), .A2(new_n439), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n824), .A2(new_n372), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n530), .A2(G113gat), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n822), .B1(new_n826), .B2(new_n827), .ZN(G1340gat));
  NAND3_X1  g627(.A1(new_n821), .A2(new_n291), .A3(new_n631), .ZN(new_n829));
  INV_X1    g628(.A(new_n826), .ZN(new_n830));
  OAI21_X1  g629(.A(G120gat), .B1(new_n830), .B2(new_n630), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n831), .A2(KEYINPUT112), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n831), .A2(KEYINPUT112), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n829), .B1(new_n832), .B2(new_n833), .ZN(G1341gat));
  NOR3_X1   g633(.A1(new_n820), .A2(new_n452), .A3(new_n555), .ZN(new_n835));
  OR2_X1    g634(.A1(new_n835), .A2(KEYINPUT113), .ZN(new_n836));
  AOI21_X1  g635(.A(G127gat), .B1(new_n835), .B2(KEYINPUT113), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n556), .A2(G127gat), .ZN(new_n838));
  AOI22_X1  g637(.A1(new_n836), .A2(new_n837), .B1(new_n826), .B2(new_n838), .ZN(G1342gat));
  NAND2_X1  g638(.A1(new_n405), .A2(new_n599), .ZN(new_n840));
  XOR2_X1   g639(.A(new_n840), .B(KEYINPUT114), .Z(new_n841));
  OR3_X1    g640(.A1(new_n820), .A2(G134gat), .A3(new_n841), .ZN(new_n842));
  OR2_X1    g641(.A1(new_n842), .A2(KEYINPUT56), .ZN(new_n843));
  OAI21_X1  g642(.A(G134gat), .B1(new_n830), .B2(new_n600), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n842), .A2(KEYINPUT56), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(G1343gat));
  INV_X1    g645(.A(new_n212), .ZN(new_n847));
  INV_X1    g646(.A(new_n818), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n808), .B(new_n849), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n795), .A2(new_n530), .A3(new_n625), .A4(new_n796), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n815), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n600), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n853), .A2(new_n806), .A3(new_n812), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n848), .B1(new_n854), .B2(new_n555), .ZN(new_n855));
  OAI21_X1  g654(.A(KEYINPUT57), .B1(new_n855), .B2(new_n274), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n274), .B1(new_n817), .B2(new_n818), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n647), .A2(new_n824), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n860), .B(KEYINPUT115), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n856), .A2(new_n859), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n847), .B1(new_n862), .B2(new_n531), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n647), .A2(new_n694), .ZN(new_n864));
  AOI211_X1 g663(.A(new_n439), .B(new_n864), .C1(new_n817), .C2(new_n818), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n865), .A2(new_n405), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n866), .A2(new_n210), .A3(new_n530), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(KEYINPUT58), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT58), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n863), .A2(new_n870), .A3(new_n867), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n869), .A2(new_n871), .ZN(G1344gat));
  INV_X1    g671(.A(G148gat), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n866), .A2(new_n873), .A3(new_n631), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n862), .A2(new_n630), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n875), .A2(KEYINPUT59), .A3(new_n873), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT59), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n817), .A2(new_n818), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n858), .B1(new_n878), .B2(new_n694), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n274), .A2(KEYINPUT57), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n809), .A2(new_n810), .A3(new_n795), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n853), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n555), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n881), .B1(new_n884), .B2(new_n818), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n879), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(new_n631), .A3(new_n861), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n877), .B1(new_n887), .B2(G148gat), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n874), .B1(new_n876), .B2(new_n888), .ZN(G1345gat));
  OAI21_X1  g688(.A(G155gat), .B1(new_n862), .B2(new_n555), .ZN(new_n890));
  INV_X1    g689(.A(G155gat), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n866), .A2(new_n891), .A3(new_n556), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT117), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n890), .A2(KEYINPUT117), .A3(new_n892), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(G1346gat));
  OAI21_X1  g696(.A(G162gat), .B1(new_n862), .B2(new_n600), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n841), .A2(G162gat), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n865), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(KEYINPUT118), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT118), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n898), .A2(new_n903), .A3(new_n900), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n902), .A2(new_n904), .ZN(G1347gat));
  NOR2_X1   g704(.A1(new_n405), .A2(new_n453), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n372), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n823), .A2(new_n907), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n908), .A2(new_n301), .A3(new_n531), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n453), .B1(new_n817), .B2(new_n818), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n702), .A2(new_n452), .ZN(new_n911));
  OR2_X1    g710(.A1(new_n911), .A2(KEYINPUT119), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(KEYINPUT119), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n910), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(new_n530), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n909), .B1(new_n916), .B2(new_n301), .ZN(G1348gat));
  OAI21_X1  g716(.A(G176gat), .B1(new_n908), .B2(new_n630), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n631), .A2(new_n302), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n918), .B1(new_n914), .B2(new_n919), .ZN(G1349gat));
  OAI21_X1  g719(.A(G183gat), .B1(new_n908), .B2(new_n555), .ZN(new_n921));
  NAND2_X1  g720(.A1(KEYINPUT120), .A2(KEYINPUT60), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n556), .A2(new_n330), .ZN(new_n923));
  OAI211_X1 g722(.A(new_n921), .B(new_n922), .C1(new_n914), .C2(new_n923), .ZN(new_n924));
  NOR2_X1   g723(.A1(KEYINPUT120), .A2(KEYINPUT60), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT121), .ZN(new_n926));
  XOR2_X1   g725(.A(new_n924), .B(new_n926), .Z(G1350gat));
  NAND3_X1  g726(.A1(new_n915), .A2(new_n331), .A3(new_n599), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n823), .A2(new_n599), .A3(new_n907), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT61), .ZN(new_n930));
  AND3_X1   g729(.A1(new_n929), .A2(new_n930), .A3(G190gat), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n930), .B1(new_n929), .B2(G190gat), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n928), .B1(new_n931), .B2(new_n932), .ZN(G1351gat));
  NOR2_X1   g732(.A1(new_n864), .A2(new_n405), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n910), .A2(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(G197gat), .B1(new_n936), .B2(new_n530), .ZN(new_n937));
  OAI21_X1  g736(.A(KEYINPUT122), .B1(new_n879), .B2(new_n885), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n556), .B1(new_n853), .B2(new_n882), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n880), .B1(new_n939), .B2(new_n848), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT122), .ZN(new_n941));
  OAI211_X1 g740(.A(new_n940), .B(new_n941), .C1(new_n857), .C2(new_n858), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n938), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n647), .A2(new_n906), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT123), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n944), .B(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  AND3_X1   g746(.A1(new_n947), .A2(G197gat), .A3(new_n530), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n937), .B1(new_n943), .B2(new_n948), .ZN(G1352gat));
  INV_X1    g748(.A(G204gat), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n910), .A2(new_n950), .A3(new_n631), .A4(new_n934), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT62), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n951), .B(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n947), .A2(new_n631), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n954), .B1(new_n938), .B2(new_n942), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n953), .B1(new_n955), .B2(new_n950), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(KEYINPUT124), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT124), .ZN(new_n958));
  OAI211_X1 g757(.A(new_n953), .B(new_n958), .C1(new_n955), .C2(new_n950), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n957), .A2(new_n959), .ZN(G1353gat));
  INV_X1    g759(.A(new_n879), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n946), .A2(new_n555), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n961), .A2(new_n962), .A3(new_n940), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(KEYINPUT126), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT126), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n886), .A2(new_n965), .A3(new_n962), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n964), .A2(G211gat), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(KEYINPUT63), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n935), .A2(G211gat), .A3(new_n555), .ZN(new_n969));
  XOR2_X1   g768(.A(new_n969), .B(KEYINPUT125), .Z(new_n970));
  INV_X1    g769(.A(KEYINPUT63), .ZN(new_n971));
  NAND4_X1  g770(.A1(new_n964), .A2(new_n971), .A3(G211gat), .A4(new_n966), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n968), .A2(new_n970), .A3(new_n972), .ZN(G1354gat));
  AOI21_X1  g772(.A(G218gat), .B1(new_n936), .B2(new_n599), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n599), .A2(G218gat), .ZN(new_n975));
  XNOR2_X1  g774(.A(new_n975), .B(KEYINPUT127), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n946), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n974), .B1(new_n943), .B2(new_n977), .ZN(G1355gat));
endmodule


