

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U545 ( .A1(n611), .A2(G2105), .ZN(n909) );
  XOR2_X1 U546 ( .A(KEYINPUT1), .B(n552), .Z(n807) );
  XNOR2_X2 U547 ( .A(KEYINPUT65), .B(G2104), .ZN(n611) );
  NOR2_X1 U548 ( .A1(n650), .A2(n966), .ZN(n628) );
  XNOR2_X2 U549 ( .A(n626), .B(KEYINPUT64), .ZN(n650) );
  INV_X1 U550 ( .A(KEYINPUT95), .ZN(n658) );
  NAND2_X1 U551 ( .A1(n516), .A2(G299), .ZN(n515) );
  NOR2_X1 U552 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U553 ( .A1(n522), .A2(n519), .ZN(n523) );
  AND2_X1 U554 ( .A1(n524), .A2(n520), .ZN(n519) );
  OR2_X1 U555 ( .A1(n696), .A2(n528), .ZN(n522) );
  AND2_X1 U556 ( .A1(n525), .A2(G8), .ZN(n524) );
  XNOR2_X1 U557 ( .A(n718), .B(n617), .ZN(n625) );
  INV_X1 U558 ( .A(KEYINPUT40), .ZN(n539) );
  NAND2_X1 U559 ( .A1(n538), .A2(n535), .ZN(n534) );
  NAND2_X1 U560 ( .A1(n777), .A2(n536), .ZN(n535) );
  NAND2_X1 U561 ( .A1(n540), .A2(n539), .ZN(n538) );
  NAND2_X1 U562 ( .A1(n537), .A2(n539), .ZN(n536) );
  NOR2_X1 U563 ( .A1(n655), .A2(n1031), .ZN(n649) );
  XNOR2_X1 U564 ( .A(n515), .B(KEYINPUT28), .ZN(n514) );
  NOR2_X1 U565 ( .A1(n679), .A2(n678), .ZN(n680) );
  NAND2_X1 U566 ( .A1(n526), .A2(KEYINPUT99), .ZN(n525) );
  INV_X1 U567 ( .A(n689), .ZN(n526) );
  NAND2_X1 U568 ( .A1(n689), .A2(n530), .ZN(n528) );
  NAND2_X1 U569 ( .A1(n527), .A2(n521), .ZN(n520) );
  INV_X1 U570 ( .A(n528), .ZN(n527) );
  INV_X1 U571 ( .A(G286), .ZN(n521) );
  NAND2_X1 U572 ( .A1(n616), .A2(n615), .ZN(n718) );
  NOR2_X1 U573 ( .A1(n529), .A2(n523), .ZN(n691) );
  INV_X1 U574 ( .A(n763), .ZN(n537) );
  INV_X1 U575 ( .A(n777), .ZN(n540) );
  NAND2_X1 U576 ( .A1(n545), .A2(n544), .ZN(n543) );
  INV_X1 U577 ( .A(G2105), .ZN(n545) );
  INV_X1 U578 ( .A(G2104), .ZN(n544) );
  NOR2_X1 U579 ( .A1(n636), .A2(n635), .ZN(n638) );
  AND2_X1 U580 ( .A1(n541), .A2(n534), .ZN(n533) );
  NAND2_X1 U581 ( .A1(n777), .A2(n539), .ZN(n532) );
  AND2_X1 U582 ( .A1(G286), .A2(KEYINPUT99), .ZN(n509) );
  NOR2_X1 U583 ( .A1(G164), .A2(G1384), .ZN(n717) );
  XOR2_X1 U584 ( .A(n621), .B(KEYINPUT84), .Z(n510) );
  AND2_X1 U585 ( .A1(n650), .A2(G1341), .ZN(n511) );
  AND2_X1 U586 ( .A1(n546), .A2(n510), .ZN(G164) );
  INV_X1 U587 ( .A(KEYINPUT99), .ZN(n530) );
  AND2_X1 U588 ( .A1(n763), .A2(KEYINPUT40), .ZN(n512) );
  XNOR2_X1 U589 ( .A(n513), .B(KEYINPUT29), .ZN(n672) );
  NAND2_X1 U590 ( .A1(n517), .A2(n514), .ZN(n513) );
  INV_X1 U591 ( .A(n665), .ZN(n516) );
  NAND2_X1 U592 ( .A1(n518), .A2(n663), .ZN(n517) );
  XNOR2_X1 U593 ( .A(n659), .B(n658), .ZN(n518) );
  AND2_X1 U594 ( .A1(n696), .A2(n509), .ZN(n529) );
  NAND2_X1 U595 ( .A1(n533), .A2(n531), .ZN(G329) );
  OR2_X1 U596 ( .A1(n542), .A2(n532), .ZN(n531) );
  NAND2_X1 U597 ( .A1(n542), .A2(n512), .ZN(n541) );
  XNOR2_X1 U598 ( .A(n762), .B(KEYINPUT100), .ZN(n542) );
  XNOR2_X2 U599 ( .A(n543), .B(KEYINPUT17), .ZN(n904) );
  NAND2_X1 U600 ( .A1(n625), .A2(n717), .ZN(n626) );
  XNOR2_X1 U601 ( .A(n624), .B(KEYINPUT85), .ZN(n546) );
  XNOR2_X1 U602 ( .A(n628), .B(n627), .ZN(n639) );
  NOR2_X1 U603 ( .A1(n1018), .A2(n511), .ZN(n547) );
  NOR2_X1 U604 ( .A1(n746), .A2(n738), .ZN(n548) );
  AND2_X1 U605 ( .A1(n761), .A2(n760), .ZN(n549) );
  AND2_X1 U606 ( .A1(n742), .A2(n741), .ZN(n550) );
  XNOR2_X1 U607 ( .A(KEYINPUT96), .B(KEYINPUT30), .ZN(n674) );
  INV_X1 U608 ( .A(KEYINPUT88), .ZN(n617) );
  INV_X1 U609 ( .A(G40), .ZN(n614) );
  INV_X1 U610 ( .A(n787), .ZN(n616) );
  INV_X1 U611 ( .A(KEYINPUT13), .ZN(n633) );
  NOR2_X1 U612 ( .A1(G543), .A2(n553), .ZN(n552) );
  NOR2_X1 U613 ( .A1(n590), .A2(n553), .ZN(n812) );
  NOR2_X1 U614 ( .A1(G543), .A2(G651), .ZN(n811) );
  AND2_X2 U615 ( .A1(G2105), .A2(G2104), .ZN(n908) );
  NOR2_X1 U616 ( .A1(n590), .A2(G651), .ZN(n808) );
  NAND2_X1 U617 ( .A1(n638), .A2(n637), .ZN(n1018) );
  XOR2_X1 U618 ( .A(KEYINPUT0), .B(G543), .Z(n590) );
  NAND2_X1 U619 ( .A1(G53), .A2(n808), .ZN(n551) );
  XNOR2_X1 U620 ( .A(n551), .B(KEYINPUT70), .ZN(n560) );
  INV_X1 U621 ( .A(G651), .ZN(n553) );
  NAND2_X1 U622 ( .A1(G65), .A2(n807), .ZN(n555) );
  NAND2_X1 U623 ( .A1(G78), .A2(n812), .ZN(n554) );
  NAND2_X1 U624 ( .A1(n555), .A2(n554), .ZN(n558) );
  NAND2_X1 U625 ( .A1(G91), .A2(n811), .ZN(n556) );
  XNOR2_X1 U626 ( .A(KEYINPUT69), .B(n556), .ZN(n557) );
  NOR2_X1 U627 ( .A1(n558), .A2(n557), .ZN(n559) );
  NAND2_X1 U628 ( .A1(n560), .A2(n559), .ZN(G299) );
  NAND2_X1 U629 ( .A1(G64), .A2(n807), .ZN(n562) );
  NAND2_X1 U630 ( .A1(G52), .A2(n808), .ZN(n561) );
  NAND2_X1 U631 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U632 ( .A(KEYINPUT68), .B(n563), .ZN(n568) );
  NAND2_X1 U633 ( .A1(G90), .A2(n811), .ZN(n565) );
  NAND2_X1 U634 ( .A1(G77), .A2(n812), .ZN(n564) );
  NAND2_X1 U635 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U636 ( .A(KEYINPUT9), .B(n566), .Z(n567) );
  NOR2_X1 U637 ( .A1(n568), .A2(n567), .ZN(G171) );
  NAND2_X1 U638 ( .A1(G63), .A2(n807), .ZN(n570) );
  NAND2_X1 U639 ( .A1(G51), .A2(n808), .ZN(n569) );
  NAND2_X1 U640 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U641 ( .A(KEYINPUT6), .B(n571), .ZN(n577) );
  NAND2_X1 U642 ( .A1(n811), .A2(G89), .ZN(n572) );
  XNOR2_X1 U643 ( .A(n572), .B(KEYINPUT4), .ZN(n574) );
  NAND2_X1 U644 ( .A1(G76), .A2(n812), .ZN(n573) );
  NAND2_X1 U645 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U646 ( .A(n575), .B(KEYINPUT5), .Z(n576) );
  NOR2_X1 U647 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U648 ( .A(KEYINPUT7), .B(n578), .Z(n579) );
  XOR2_X1 U649 ( .A(KEYINPUT73), .B(n579), .Z(G168) );
  XOR2_X1 U650 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U651 ( .A1(n807), .A2(G62), .ZN(n582) );
  NAND2_X1 U652 ( .A1(G50), .A2(n808), .ZN(n580) );
  XOR2_X1 U653 ( .A(KEYINPUT77), .B(n580), .Z(n581) );
  NAND2_X1 U654 ( .A1(n582), .A2(n581), .ZN(n586) );
  NAND2_X1 U655 ( .A1(G88), .A2(n811), .ZN(n584) );
  NAND2_X1 U656 ( .A1(G75), .A2(n812), .ZN(n583) );
  NAND2_X1 U657 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U658 ( .A1(n586), .A2(n585), .ZN(G166) );
  INV_X1 U659 ( .A(G166), .ZN(G303) );
  NAND2_X1 U660 ( .A1(G49), .A2(n808), .ZN(n588) );
  NAND2_X1 U661 ( .A1(G74), .A2(G651), .ZN(n587) );
  NAND2_X1 U662 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U663 ( .A1(n807), .A2(n589), .ZN(n592) );
  NAND2_X1 U664 ( .A1(n590), .A2(G87), .ZN(n591) );
  NAND2_X1 U665 ( .A1(n592), .A2(n591), .ZN(G288) );
  NAND2_X1 U666 ( .A1(G61), .A2(n807), .ZN(n594) );
  NAND2_X1 U667 ( .A1(G86), .A2(n811), .ZN(n593) );
  NAND2_X1 U668 ( .A1(n594), .A2(n593), .ZN(n597) );
  NAND2_X1 U669 ( .A1(n812), .A2(G73), .ZN(n595) );
  XOR2_X1 U670 ( .A(KEYINPUT2), .B(n595), .Z(n596) );
  NOR2_X1 U671 ( .A1(n597), .A2(n596), .ZN(n599) );
  NAND2_X1 U672 ( .A1(n808), .A2(G48), .ZN(n598) );
  NAND2_X1 U673 ( .A1(n599), .A2(n598), .ZN(G305) );
  NAND2_X1 U674 ( .A1(G60), .A2(n807), .ZN(n601) );
  NAND2_X1 U675 ( .A1(G47), .A2(n808), .ZN(n600) );
  NAND2_X1 U676 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U677 ( .A(KEYINPUT67), .B(n602), .ZN(n606) );
  NAND2_X1 U678 ( .A1(G85), .A2(n811), .ZN(n604) );
  NAND2_X1 U679 ( .A1(G72), .A2(n812), .ZN(n603) );
  AND2_X1 U680 ( .A1(n604), .A2(n603), .ZN(n605) );
  NAND2_X1 U681 ( .A1(n606), .A2(n605), .ZN(G290) );
  NOR2_X2 U682 ( .A1(n611), .A2(G2105), .ZN(n705) );
  NAND2_X1 U683 ( .A1(G101), .A2(n705), .ZN(n608) );
  XOR2_X1 U684 ( .A(KEYINPUT23), .B(KEYINPUT66), .Z(n607) );
  XNOR2_X1 U685 ( .A(n608), .B(n607), .ZN(n610) );
  NAND2_X1 U686 ( .A1(n908), .A2(G113), .ZN(n609) );
  NAND2_X1 U687 ( .A1(n610), .A2(n609), .ZN(n787) );
  NAND2_X1 U688 ( .A1(G137), .A2(n904), .ZN(n613) );
  NAND2_X1 U689 ( .A1(G125), .A2(n909), .ZN(n612) );
  NAND2_X1 U690 ( .A1(n613), .A2(n612), .ZN(n788) );
  NOR2_X1 U691 ( .A1(n788), .A2(n614), .ZN(n615) );
  NAND2_X1 U692 ( .A1(n908), .A2(G114), .ZN(n618) );
  XOR2_X1 U693 ( .A(KEYINPUT83), .B(n618), .Z(n620) );
  NAND2_X1 U694 ( .A1(n909), .A2(G126), .ZN(n619) );
  NAND2_X1 U695 ( .A1(n620), .A2(n619), .ZN(n621) );
  NAND2_X1 U696 ( .A1(G138), .A2(n904), .ZN(n623) );
  NAND2_X1 U697 ( .A1(G102), .A2(n705), .ZN(n622) );
  NAND2_X1 U698 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U699 ( .A(G1996), .B(KEYINPUT93), .ZN(n966) );
  INV_X1 U700 ( .A(KEYINPUT26), .ZN(n627) );
  NAND2_X1 U701 ( .A1(G56), .A2(n807), .ZN(n629) );
  XOR2_X1 U702 ( .A(KEYINPUT14), .B(n629), .Z(n636) );
  NAND2_X1 U703 ( .A1(G68), .A2(n812), .ZN(n632) );
  NAND2_X1 U704 ( .A1(n811), .A2(G81), .ZN(n630) );
  XNOR2_X1 U705 ( .A(n630), .B(KEYINPUT12), .ZN(n631) );
  NAND2_X1 U706 ( .A1(n632), .A2(n631), .ZN(n634) );
  XNOR2_X1 U707 ( .A(n634), .B(n633), .ZN(n635) );
  NAND2_X1 U708 ( .A1(n808), .A2(G43), .ZN(n637) );
  NAND2_X1 U709 ( .A1(n639), .A2(n547), .ZN(n655) );
  NAND2_X1 U710 ( .A1(G54), .A2(n808), .ZN(n641) );
  NAND2_X1 U711 ( .A1(G79), .A2(n812), .ZN(n640) );
  NAND2_X1 U712 ( .A1(n641), .A2(n640), .ZN(n646) );
  NAND2_X1 U713 ( .A1(G66), .A2(n807), .ZN(n643) );
  NAND2_X1 U714 ( .A1(G92), .A2(n811), .ZN(n642) );
  NAND2_X1 U715 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U716 ( .A(KEYINPUT72), .B(n644), .ZN(n645) );
  NOR2_X1 U717 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U718 ( .A(n647), .B(KEYINPUT15), .ZN(n1031) );
  INV_X1 U719 ( .A(KEYINPUT94), .ZN(n648) );
  XNOR2_X1 U720 ( .A(n649), .B(n648), .ZN(n654) );
  INV_X1 U721 ( .A(n650), .ZN(n666) );
  NOR2_X1 U722 ( .A1(G1348), .A2(n666), .ZN(n652) );
  INV_X1 U723 ( .A(n666), .ZN(n684) );
  NOR2_X1 U724 ( .A1(n684), .A2(G2067), .ZN(n651) );
  NOR2_X1 U725 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U726 ( .A1(n654), .A2(n653), .ZN(n657) );
  NAND2_X1 U727 ( .A1(n655), .A2(n1031), .ZN(n656) );
  NAND2_X1 U728 ( .A1(n657), .A2(n656), .ZN(n659) );
  NAND2_X1 U729 ( .A1(G2072), .A2(n666), .ZN(n660) );
  XNOR2_X1 U730 ( .A(n660), .B(KEYINPUT27), .ZN(n662) );
  AND2_X1 U731 ( .A1(n684), .A2(G1956), .ZN(n661) );
  NOR2_X1 U732 ( .A1(n662), .A2(n661), .ZN(n665) );
  INV_X1 U733 ( .A(G299), .ZN(n664) );
  NAND2_X1 U734 ( .A1(n665), .A2(n664), .ZN(n663) );
  NOR2_X1 U735 ( .A1(G1961), .A2(n666), .ZN(n668) );
  XOR2_X1 U736 ( .A(G2078), .B(KEYINPUT25), .Z(n967) );
  NOR2_X1 U737 ( .A1(n684), .A2(n967), .ZN(n667) );
  NOR2_X1 U738 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U739 ( .A(KEYINPUT91), .B(n669), .ZN(n677) );
  AND2_X1 U740 ( .A1(n677), .A2(G171), .ZN(n670) );
  XNOR2_X1 U741 ( .A(n670), .B(KEYINPUT92), .ZN(n671) );
  NOR2_X1 U742 ( .A1(n672), .A2(n671), .ZN(n682) );
  NAND2_X1 U743 ( .A1(n650), .A2(G8), .ZN(n746) );
  NOR2_X1 U744 ( .A1(G1966), .A2(n746), .ZN(n695) );
  NOR2_X1 U745 ( .A1(n684), .A2(G2084), .ZN(n692) );
  NOR2_X1 U746 ( .A1(n695), .A2(n692), .ZN(n673) );
  NAND2_X1 U747 ( .A1(G8), .A2(n673), .ZN(n675) );
  XNOR2_X1 U748 ( .A(n675), .B(n674), .ZN(n676) );
  NOR2_X1 U749 ( .A1(G168), .A2(n676), .ZN(n679) );
  NOR2_X1 U750 ( .A1(G171), .A2(n677), .ZN(n678) );
  XNOR2_X1 U751 ( .A(n680), .B(KEYINPUT31), .ZN(n681) );
  XNOR2_X1 U752 ( .A(n683), .B(KEYINPUT97), .ZN(n696) );
  NOR2_X1 U753 ( .A1(n684), .A2(G2090), .ZN(n685) );
  XNOR2_X1 U754 ( .A(n685), .B(KEYINPUT98), .ZN(n687) );
  NOR2_X1 U755 ( .A1(n746), .A2(G1971), .ZN(n686) );
  NOR2_X1 U756 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U757 ( .A1(n688), .A2(G303), .ZN(n689) );
  INV_X1 U758 ( .A(KEYINPUT32), .ZN(n690) );
  XNOR2_X1 U759 ( .A(n691), .B(n690), .ZN(n753) );
  NAND2_X1 U760 ( .A1(G8), .A2(n692), .ZN(n693) );
  XOR2_X1 U761 ( .A(KEYINPUT90), .B(n693), .Z(n694) );
  NOR2_X1 U762 ( .A1(n695), .A2(n694), .ZN(n697) );
  NAND2_X1 U763 ( .A1(n697), .A2(n696), .ZN(n751) );
  NAND2_X1 U764 ( .A1(G1976), .A2(G288), .ZN(n1022) );
  AND2_X1 U765 ( .A1(n751), .A2(n1022), .ZN(n733) );
  NOR2_X1 U766 ( .A1(G1976), .A2(G288), .ZN(n736) );
  NAND2_X1 U767 ( .A1(n736), .A2(KEYINPUT33), .ZN(n698) );
  OR2_X1 U768 ( .A1(n698), .A2(n746), .ZN(n699) );
  XOR2_X1 U769 ( .A(G1981), .B(G305), .Z(n1015) );
  NAND2_X1 U770 ( .A1(n699), .A2(n1015), .ZN(n731) );
  NAND2_X1 U771 ( .A1(G131), .A2(n904), .ZN(n701) );
  NAND2_X1 U772 ( .A1(G119), .A2(n909), .ZN(n700) );
  NAND2_X1 U773 ( .A1(n701), .A2(n700), .ZN(n704) );
  NAND2_X1 U774 ( .A1(G107), .A2(n908), .ZN(n702) );
  XNOR2_X1 U775 ( .A(KEYINPUT87), .B(n702), .ZN(n703) );
  NOR2_X1 U776 ( .A1(n704), .A2(n703), .ZN(n707) );
  NAND2_X1 U777 ( .A1(n705), .A2(G95), .ZN(n706) );
  NAND2_X1 U778 ( .A1(n707), .A2(n706), .ZN(n918) );
  AND2_X1 U779 ( .A1(n918), .A2(G1991), .ZN(n716) );
  NAND2_X1 U780 ( .A1(G141), .A2(n904), .ZN(n709) );
  NAND2_X1 U781 ( .A1(G117), .A2(n908), .ZN(n708) );
  NAND2_X1 U782 ( .A1(n709), .A2(n708), .ZN(n712) );
  NAND2_X1 U783 ( .A1(n705), .A2(G105), .ZN(n710) );
  XOR2_X1 U784 ( .A(KEYINPUT38), .B(n710), .Z(n711) );
  NOR2_X1 U785 ( .A1(n712), .A2(n711), .ZN(n714) );
  NAND2_X1 U786 ( .A1(n909), .A2(G129), .ZN(n713) );
  NAND2_X1 U787 ( .A1(n714), .A2(n713), .ZN(n919) );
  AND2_X1 U788 ( .A1(n919), .A2(G1996), .ZN(n715) );
  NOR2_X1 U789 ( .A1(n716), .A2(n715), .ZN(n991) );
  NOR2_X1 U790 ( .A1(n718), .A2(n717), .ZN(n775) );
  INV_X1 U791 ( .A(n775), .ZN(n719) );
  NOR2_X1 U792 ( .A1(n991), .A2(n719), .ZN(n767) );
  INV_X1 U793 ( .A(n767), .ZN(n730) );
  XNOR2_X1 U794 ( .A(G2067), .B(KEYINPUT37), .ZN(n772) );
  XNOR2_X1 U795 ( .A(KEYINPUT86), .B(KEYINPUT34), .ZN(n723) );
  NAND2_X1 U796 ( .A1(G140), .A2(n904), .ZN(n721) );
  NAND2_X1 U797 ( .A1(G104), .A2(n705), .ZN(n720) );
  NAND2_X1 U798 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U799 ( .A(n723), .B(n722), .ZN(n728) );
  NAND2_X1 U800 ( .A1(G116), .A2(n908), .ZN(n725) );
  NAND2_X1 U801 ( .A1(G128), .A2(n909), .ZN(n724) );
  NAND2_X1 U802 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U803 ( .A(KEYINPUT35), .B(n726), .Z(n727) );
  NOR2_X1 U804 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U805 ( .A(KEYINPUT36), .B(n729), .ZN(n926) );
  NOR2_X1 U806 ( .A1(n772), .A2(n926), .ZN(n1004) );
  NAND2_X1 U807 ( .A1(n775), .A2(n1004), .ZN(n770) );
  NAND2_X1 U808 ( .A1(n730), .A2(n770), .ZN(n747) );
  OR2_X1 U809 ( .A1(n731), .A2(n747), .ZN(n740) );
  INV_X1 U810 ( .A(n740), .ZN(n732) );
  AND2_X1 U811 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U812 ( .A1(n753), .A2(n734), .ZN(n742) );
  INV_X1 U813 ( .A(n1022), .ZN(n737) );
  NOR2_X1 U814 ( .A1(G1971), .A2(G303), .ZN(n735) );
  NOR2_X1 U815 ( .A1(n736), .A2(n735), .ZN(n1026) );
  OR2_X1 U816 ( .A1(n737), .A2(n1026), .ZN(n738) );
  NOR2_X1 U817 ( .A1(KEYINPUT33), .A2(n548), .ZN(n739) );
  OR2_X1 U818 ( .A1(n740), .A2(n739), .ZN(n741) );
  NOR2_X1 U819 ( .A1(G1981), .A2(G305), .ZN(n743) );
  XOR2_X1 U820 ( .A(n743), .B(KEYINPUT24), .Z(n744) );
  NOR2_X1 U821 ( .A1(n746), .A2(n744), .ZN(n745) );
  XOR2_X1 U822 ( .A(KEYINPUT89), .B(n745), .Z(n755) );
  OR2_X1 U823 ( .A1(n755), .A2(n746), .ZN(n749) );
  INV_X1 U824 ( .A(n747), .ZN(n748) );
  NAND2_X1 U825 ( .A1(n749), .A2(n748), .ZN(n759) );
  INV_X1 U826 ( .A(n759), .ZN(n750) );
  AND2_X1 U827 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U828 ( .A1(n753), .A2(n752), .ZN(n761) );
  NOR2_X1 U829 ( .A1(G2090), .A2(G303), .ZN(n754) );
  NAND2_X1 U830 ( .A1(G8), .A2(n754), .ZN(n757) );
  INV_X1 U831 ( .A(n755), .ZN(n756) );
  AND2_X1 U832 ( .A1(n757), .A2(n756), .ZN(n758) );
  OR2_X1 U833 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U834 ( .A1(n550), .A2(n549), .ZN(n762) );
  XNOR2_X1 U835 ( .A(G1986), .B(G290), .ZN(n1020) );
  NAND2_X1 U836 ( .A1(n775), .A2(n1020), .ZN(n763) );
  NOR2_X1 U837 ( .A1(G1996), .A2(n919), .ZN(n1007) );
  NOR2_X1 U838 ( .A1(G1986), .A2(G290), .ZN(n765) );
  NOR2_X1 U839 ( .A1(G1991), .A2(n918), .ZN(n764) );
  XOR2_X1 U840 ( .A(KEYINPUT101), .B(n764), .Z(n1001) );
  NOR2_X1 U841 ( .A1(n765), .A2(n1001), .ZN(n766) );
  NOR2_X1 U842 ( .A1(n767), .A2(n766), .ZN(n768) );
  NOR2_X1 U843 ( .A1(n1007), .A2(n768), .ZN(n769) );
  XNOR2_X1 U844 ( .A(n769), .B(KEYINPUT39), .ZN(n771) );
  NAND2_X1 U845 ( .A1(n771), .A2(n770), .ZN(n773) );
  NAND2_X1 U846 ( .A1(n772), .A2(n926), .ZN(n990) );
  NAND2_X1 U847 ( .A1(n773), .A2(n990), .ZN(n774) );
  NAND2_X1 U848 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U849 ( .A(n776), .B(KEYINPUT102), .ZN(n777) );
  AND2_X1 U850 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U851 ( .A1(G135), .A2(n904), .ZN(n780) );
  NAND2_X1 U852 ( .A1(G111), .A2(n908), .ZN(n779) );
  NAND2_X1 U853 ( .A1(n780), .A2(n779), .ZN(n783) );
  NAND2_X1 U854 ( .A1(n909), .A2(G123), .ZN(n781) );
  XOR2_X1 U855 ( .A(KEYINPUT18), .B(n781), .Z(n782) );
  NOR2_X1 U856 ( .A1(n783), .A2(n782), .ZN(n785) );
  NAND2_X1 U857 ( .A1(n705), .A2(G99), .ZN(n784) );
  NAND2_X1 U858 ( .A1(n785), .A2(n784), .ZN(n998) );
  XNOR2_X1 U859 ( .A(G2096), .B(n998), .ZN(n786) );
  OR2_X1 U860 ( .A1(G2100), .A2(n786), .ZN(G156) );
  INV_X1 U861 ( .A(G132), .ZN(G219) );
  INV_X1 U862 ( .A(G120), .ZN(G236) );
  INV_X1 U863 ( .A(G69), .ZN(G235) );
  INV_X1 U864 ( .A(G108), .ZN(G238) );
  NOR2_X1 U865 ( .A1(n788), .A2(n787), .ZN(G160) );
  NAND2_X1 U866 ( .A1(G7), .A2(G661), .ZN(n789) );
  XNOR2_X1 U867 ( .A(n789), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U868 ( .A(G223), .ZN(n855) );
  NAND2_X1 U869 ( .A1(n855), .A2(G567), .ZN(n790) );
  XOR2_X1 U870 ( .A(KEYINPUT11), .B(n790), .Z(G234) );
  INV_X1 U871 ( .A(G860), .ZN(n795) );
  OR2_X1 U872 ( .A1(n1018), .A2(n795), .ZN(G153) );
  INV_X1 U873 ( .A(G171), .ZN(G301) );
  NAND2_X1 U874 ( .A1(G868), .A2(G301), .ZN(n792) );
  INV_X1 U875 ( .A(G868), .ZN(n798) );
  NAND2_X1 U876 ( .A1(n1031), .A2(n798), .ZN(n791) );
  NAND2_X1 U877 ( .A1(n792), .A2(n791), .ZN(G284) );
  NOR2_X1 U878 ( .A1(G286), .A2(n798), .ZN(n794) );
  NOR2_X1 U879 ( .A1(G868), .A2(G299), .ZN(n793) );
  NOR2_X1 U880 ( .A1(n794), .A2(n793), .ZN(G297) );
  NAND2_X1 U881 ( .A1(n795), .A2(G559), .ZN(n796) );
  INV_X1 U882 ( .A(n1031), .ZN(n803) );
  NAND2_X1 U883 ( .A1(n796), .A2(n803), .ZN(n797) );
  XNOR2_X1 U884 ( .A(n797), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U885 ( .A1(n1031), .A2(n798), .ZN(n799) );
  XOR2_X1 U886 ( .A(KEYINPUT74), .B(n799), .Z(n800) );
  NOR2_X1 U887 ( .A1(G559), .A2(n800), .ZN(n802) );
  NOR2_X1 U888 ( .A1(G868), .A2(n1018), .ZN(n801) );
  NOR2_X1 U889 ( .A1(n802), .A2(n801), .ZN(G282) );
  NAND2_X1 U890 ( .A1(G559), .A2(n803), .ZN(n804) );
  XNOR2_X1 U891 ( .A(n804), .B(n1018), .ZN(n818) );
  XOR2_X1 U892 ( .A(n818), .B(KEYINPUT75), .Z(n805) );
  NOR2_X1 U893 ( .A1(G860), .A2(n805), .ZN(n806) );
  XOR2_X1 U894 ( .A(KEYINPUT76), .B(n806), .Z(n817) );
  NAND2_X1 U895 ( .A1(G67), .A2(n807), .ZN(n810) );
  NAND2_X1 U896 ( .A1(G55), .A2(n808), .ZN(n809) );
  NAND2_X1 U897 ( .A1(n810), .A2(n809), .ZN(n816) );
  NAND2_X1 U898 ( .A1(G93), .A2(n811), .ZN(n814) );
  NAND2_X1 U899 ( .A1(G80), .A2(n812), .ZN(n813) );
  NAND2_X1 U900 ( .A1(n814), .A2(n813), .ZN(n815) );
  NOR2_X1 U901 ( .A1(n816), .A2(n815), .ZN(n828) );
  XOR2_X1 U902 ( .A(n817), .B(n828), .Z(G145) );
  XNOR2_X1 U903 ( .A(KEYINPUT80), .B(n818), .ZN(n826) );
  XNOR2_X1 U904 ( .A(KEYINPUT79), .B(KEYINPUT19), .ZN(n820) );
  XNOR2_X1 U905 ( .A(G288), .B(KEYINPUT78), .ZN(n819) );
  XNOR2_X1 U906 ( .A(n820), .B(n819), .ZN(n821) );
  XNOR2_X1 U907 ( .A(n828), .B(n821), .ZN(n823) );
  XNOR2_X1 U908 ( .A(G290), .B(G166), .ZN(n822) );
  XNOR2_X1 U909 ( .A(n823), .B(n822), .ZN(n824) );
  XNOR2_X1 U910 ( .A(n824), .B(G305), .ZN(n825) );
  XNOR2_X1 U911 ( .A(n825), .B(G299), .ZN(n864) );
  XNOR2_X1 U912 ( .A(n826), .B(n864), .ZN(n827) );
  NAND2_X1 U913 ( .A1(n827), .A2(G868), .ZN(n830) );
  OR2_X1 U914 ( .A1(n828), .A2(G868), .ZN(n829) );
  NAND2_X1 U915 ( .A1(n830), .A2(n829), .ZN(G295) );
  NAND2_X1 U916 ( .A1(G2078), .A2(G2084), .ZN(n831) );
  XOR2_X1 U917 ( .A(KEYINPUT20), .B(n831), .Z(n832) );
  NAND2_X1 U918 ( .A1(G2090), .A2(n832), .ZN(n833) );
  XNOR2_X1 U919 ( .A(KEYINPUT21), .B(n833), .ZN(n834) );
  NAND2_X1 U920 ( .A1(n834), .A2(G2072), .ZN(G158) );
  XOR2_X1 U921 ( .A(KEYINPUT81), .B(G44), .Z(n835) );
  XNOR2_X1 U922 ( .A(KEYINPUT3), .B(n835), .ZN(G218) );
  XNOR2_X1 U923 ( .A(KEYINPUT71), .B(G82), .ZN(G220) );
  NOR2_X1 U924 ( .A1(G235), .A2(G236), .ZN(n836) );
  XOR2_X1 U925 ( .A(KEYINPUT82), .B(n836), .Z(n837) );
  NOR2_X1 U926 ( .A1(G238), .A2(n837), .ZN(n838) );
  NAND2_X1 U927 ( .A1(G57), .A2(n838), .ZN(n861) );
  NAND2_X1 U928 ( .A1(n861), .A2(G567), .ZN(n843) );
  NOR2_X1 U929 ( .A1(G219), .A2(G220), .ZN(n839) );
  XOR2_X1 U930 ( .A(KEYINPUT22), .B(n839), .Z(n840) );
  NOR2_X1 U931 ( .A1(G218), .A2(n840), .ZN(n841) );
  NAND2_X1 U932 ( .A1(G96), .A2(n841), .ZN(n862) );
  NAND2_X1 U933 ( .A1(n862), .A2(G2106), .ZN(n842) );
  NAND2_X1 U934 ( .A1(n843), .A2(n842), .ZN(n869) );
  NAND2_X1 U935 ( .A1(G483), .A2(G661), .ZN(n844) );
  NOR2_X1 U936 ( .A1(n869), .A2(n844), .ZN(n860) );
  NAND2_X1 U937 ( .A1(n860), .A2(G36), .ZN(G176) );
  XOR2_X1 U938 ( .A(G2430), .B(G2451), .Z(n846) );
  XNOR2_X1 U939 ( .A(G2446), .B(G2427), .ZN(n845) );
  XNOR2_X1 U940 ( .A(n846), .B(n845), .ZN(n853) );
  XOR2_X1 U941 ( .A(G2438), .B(KEYINPUT103), .Z(n848) );
  XNOR2_X1 U942 ( .A(G2443), .B(G2454), .ZN(n847) );
  XNOR2_X1 U943 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U944 ( .A(n849), .B(G2435), .Z(n851) );
  XNOR2_X1 U945 ( .A(G1341), .B(G1348), .ZN(n850) );
  XNOR2_X1 U946 ( .A(n851), .B(n850), .ZN(n852) );
  XNOR2_X1 U947 ( .A(n853), .B(n852), .ZN(n854) );
  NAND2_X1 U948 ( .A1(n854), .A2(G14), .ZN(n929) );
  XOR2_X1 U949 ( .A(KEYINPUT104), .B(n929), .Z(G401) );
  NAND2_X1 U950 ( .A1(G2106), .A2(n855), .ZN(G217) );
  NAND2_X1 U951 ( .A1(G15), .A2(G2), .ZN(n857) );
  INV_X1 U952 ( .A(G661), .ZN(n856) );
  NOR2_X1 U953 ( .A1(n857), .A2(n856), .ZN(n858) );
  XNOR2_X1 U954 ( .A(n858), .B(KEYINPUT105), .ZN(G259) );
  NAND2_X1 U955 ( .A1(G3), .A2(G1), .ZN(n859) );
  NAND2_X1 U956 ( .A1(n860), .A2(n859), .ZN(G188) );
  INV_X1 U958 ( .A(G96), .ZN(G221) );
  NOR2_X1 U959 ( .A1(n862), .A2(n861), .ZN(G325) );
  INV_X1 U960 ( .A(G325), .ZN(G261) );
  XOR2_X1 U961 ( .A(n1031), .B(n1018), .Z(n863) );
  XOR2_X1 U962 ( .A(n863), .B(KEYINPUT110), .Z(n866) );
  XNOR2_X1 U963 ( .A(G171), .B(n864), .ZN(n865) );
  XNOR2_X1 U964 ( .A(n866), .B(n865), .ZN(n867) );
  XNOR2_X1 U965 ( .A(n867), .B(G286), .ZN(n868) );
  NOR2_X1 U966 ( .A1(G37), .A2(n868), .ZN(G397) );
  INV_X1 U967 ( .A(n869), .ZN(G319) );
  XOR2_X1 U968 ( .A(G2096), .B(KEYINPUT43), .Z(n871) );
  XNOR2_X1 U969 ( .A(G2072), .B(KEYINPUT42), .ZN(n870) );
  XNOR2_X1 U970 ( .A(n871), .B(n870), .ZN(n872) );
  XOR2_X1 U971 ( .A(n872), .B(G2678), .Z(n874) );
  XNOR2_X1 U972 ( .A(G2067), .B(G2090), .ZN(n873) );
  XNOR2_X1 U973 ( .A(n874), .B(n873), .ZN(n878) );
  XOR2_X1 U974 ( .A(KEYINPUT106), .B(G2100), .Z(n876) );
  XNOR2_X1 U975 ( .A(G2078), .B(G2084), .ZN(n875) );
  XNOR2_X1 U976 ( .A(n876), .B(n875), .ZN(n877) );
  XNOR2_X1 U977 ( .A(n878), .B(n877), .ZN(G227) );
  XOR2_X1 U978 ( .A(G1961), .B(G1971), .Z(n880) );
  XNOR2_X1 U979 ( .A(G1981), .B(G1976), .ZN(n879) );
  XNOR2_X1 U980 ( .A(n880), .B(n879), .ZN(n884) );
  XOR2_X1 U981 ( .A(G1991), .B(G1996), .Z(n882) );
  XNOR2_X1 U982 ( .A(G1966), .B(G1956), .ZN(n881) );
  XNOR2_X1 U983 ( .A(n882), .B(n881), .ZN(n883) );
  XOR2_X1 U984 ( .A(n884), .B(n883), .Z(n886) );
  XNOR2_X1 U985 ( .A(G2474), .B(KEYINPUT41), .ZN(n885) );
  XNOR2_X1 U986 ( .A(n886), .B(n885), .ZN(n888) );
  XOR2_X1 U987 ( .A(G1986), .B(KEYINPUT107), .Z(n887) );
  XNOR2_X1 U988 ( .A(n888), .B(n887), .ZN(G229) );
  NAND2_X1 U989 ( .A1(G124), .A2(n909), .ZN(n889) );
  XNOR2_X1 U990 ( .A(n889), .B(KEYINPUT44), .ZN(n891) );
  NAND2_X1 U991 ( .A1(n908), .A2(G112), .ZN(n890) );
  NAND2_X1 U992 ( .A1(n891), .A2(n890), .ZN(n895) );
  NAND2_X1 U993 ( .A1(G136), .A2(n904), .ZN(n893) );
  NAND2_X1 U994 ( .A1(G100), .A2(n705), .ZN(n892) );
  NAND2_X1 U995 ( .A1(n893), .A2(n892), .ZN(n894) );
  NOR2_X1 U996 ( .A1(n895), .A2(n894), .ZN(G162) );
  NAND2_X1 U997 ( .A1(G118), .A2(n908), .ZN(n897) );
  NAND2_X1 U998 ( .A1(G130), .A2(n909), .ZN(n896) );
  NAND2_X1 U999 ( .A1(n897), .A2(n896), .ZN(n902) );
  NAND2_X1 U1000 ( .A1(G142), .A2(n904), .ZN(n899) );
  NAND2_X1 U1001 ( .A1(G106), .A2(n705), .ZN(n898) );
  NAND2_X1 U1002 ( .A1(n899), .A2(n898), .ZN(n900) );
  XOR2_X1 U1003 ( .A(KEYINPUT45), .B(n900), .Z(n901) );
  NOR2_X1 U1004 ( .A1(n902), .A2(n901), .ZN(n903) );
  XNOR2_X1 U1005 ( .A(G164), .B(n903), .ZN(n925) );
  XOR2_X1 U1006 ( .A(KEYINPUT109), .B(KEYINPUT48), .Z(n916) );
  NAND2_X1 U1007 ( .A1(G139), .A2(n904), .ZN(n906) );
  NAND2_X1 U1008 ( .A1(G103), .A2(n705), .ZN(n905) );
  NAND2_X1 U1009 ( .A1(n906), .A2(n905), .ZN(n907) );
  XNOR2_X1 U1010 ( .A(KEYINPUT108), .B(n907), .ZN(n914) );
  NAND2_X1 U1011 ( .A1(G115), .A2(n908), .ZN(n911) );
  NAND2_X1 U1012 ( .A1(G127), .A2(n909), .ZN(n910) );
  NAND2_X1 U1013 ( .A1(n911), .A2(n910), .ZN(n912) );
  XOR2_X1 U1014 ( .A(KEYINPUT47), .B(n912), .Z(n913) );
  NOR2_X1 U1015 ( .A1(n914), .A2(n913), .ZN(n992) );
  XNOR2_X1 U1016 ( .A(n992), .B(KEYINPUT46), .ZN(n915) );
  XNOR2_X1 U1017 ( .A(n916), .B(n915), .ZN(n917) );
  XOR2_X1 U1018 ( .A(n918), .B(n917), .Z(n923) );
  XNOR2_X1 U1019 ( .A(n998), .B(G162), .ZN(n921) );
  XOR2_X1 U1020 ( .A(G160), .B(n919), .Z(n920) );
  XNOR2_X1 U1021 ( .A(n921), .B(n920), .ZN(n922) );
  XNOR2_X1 U1022 ( .A(n923), .B(n922), .ZN(n924) );
  XNOR2_X1 U1023 ( .A(n925), .B(n924), .ZN(n927) );
  XOR2_X1 U1024 ( .A(n927), .B(n926), .Z(n928) );
  NOR2_X1 U1025 ( .A1(G37), .A2(n928), .ZN(G395) );
  NAND2_X1 U1026 ( .A1(G319), .A2(n929), .ZN(n930) );
  NOR2_X1 U1027 ( .A1(G397), .A2(n930), .ZN(n933) );
  NOR2_X1 U1028 ( .A1(G227), .A2(G229), .ZN(n931) );
  XOR2_X1 U1029 ( .A(KEYINPUT49), .B(n931), .Z(n932) );
  NAND2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1031 ( .A1(n934), .A2(G395), .ZN(n935) );
  XNOR2_X1 U1032 ( .A(n935), .B(KEYINPUT111), .ZN(G225) );
  INV_X1 U1033 ( .A(G225), .ZN(G308) );
  INV_X1 U1034 ( .A(G57), .ZN(G237) );
  XOR2_X1 U1035 ( .A(KEYINPUT120), .B(G16), .Z(n963) );
  XNOR2_X1 U1036 ( .A(G1986), .B(G24), .ZN(n937) );
  XNOR2_X1 U1037 ( .A(G1971), .B(G22), .ZN(n936) );
  NOR2_X1 U1038 ( .A1(n937), .A2(n936), .ZN(n939) );
  XOR2_X1 U1039 ( .A(G1976), .B(G23), .Z(n938) );
  NAND2_X1 U1040 ( .A1(n939), .A2(n938), .ZN(n941) );
  XOR2_X1 U1041 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n940) );
  XNOR2_X1 U1042 ( .A(n941), .B(n940), .ZN(n958) );
  XNOR2_X1 U1043 ( .A(G1966), .B(G21), .ZN(n955) );
  XOR2_X1 U1044 ( .A(G1981), .B(G6), .Z(n944) );
  XNOR2_X1 U1045 ( .A(G20), .B(KEYINPUT121), .ZN(n942) );
  XNOR2_X1 U1046 ( .A(n942), .B(G1956), .ZN(n943) );
  NAND2_X1 U1047 ( .A1(n944), .A2(n943), .ZN(n946) );
  XNOR2_X1 U1048 ( .A(G19), .B(G1341), .ZN(n945) );
  NOR2_X1 U1049 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1050 ( .A(KEYINPUT122), .B(n947), .ZN(n951) );
  XOR2_X1 U1051 ( .A(KEYINPUT123), .B(G4), .Z(n949) );
  XNOR2_X1 U1052 ( .A(G1348), .B(KEYINPUT59), .ZN(n948) );
  XNOR2_X1 U1053 ( .A(n949), .B(n948), .ZN(n950) );
  NAND2_X1 U1054 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1055 ( .A(n952), .B(KEYINPUT60), .ZN(n953) );
  XNOR2_X1 U1056 ( .A(n953), .B(KEYINPUT124), .ZN(n954) );
  NOR2_X1 U1057 ( .A1(n955), .A2(n954), .ZN(n956) );
  XOR2_X1 U1058 ( .A(KEYINPUT125), .B(n956), .Z(n957) );
  NAND2_X1 U1059 ( .A1(n958), .A2(n957), .ZN(n960) );
  XNOR2_X1 U1060 ( .A(G5), .B(G1961), .ZN(n959) );
  NOR2_X1 U1061 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1062 ( .A(KEYINPUT61), .B(n961), .ZN(n962) );
  NAND2_X1 U1063 ( .A1(n963), .A2(n962), .ZN(n1043) );
  XOR2_X1 U1064 ( .A(G25), .B(G1991), .Z(n964) );
  NAND2_X1 U1065 ( .A1(n964), .A2(G28), .ZN(n965) );
  XNOR2_X1 U1066 ( .A(KEYINPUT115), .B(n965), .ZN(n977) );
  XNOR2_X1 U1067 ( .A(G32), .B(n966), .ZN(n971) );
  XNOR2_X1 U1068 ( .A(G2067), .B(G26), .ZN(n969) );
  XNOR2_X1 U1069 ( .A(G27), .B(n967), .ZN(n968) );
  NOR2_X1 U1070 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1071 ( .A1(n971), .A2(n970), .ZN(n974) );
  XNOR2_X1 U1072 ( .A(KEYINPUT116), .B(G2072), .ZN(n972) );
  XNOR2_X1 U1073 ( .A(G33), .B(n972), .ZN(n973) );
  NOR2_X1 U1074 ( .A1(n974), .A2(n973), .ZN(n975) );
  XOR2_X1 U1075 ( .A(KEYINPUT117), .B(n975), .Z(n976) );
  NAND2_X1 U1076 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1077 ( .A(KEYINPUT53), .B(n978), .ZN(n982) );
  XOR2_X1 U1078 ( .A(G34), .B(KEYINPUT118), .Z(n980) );
  XNOR2_X1 U1079 ( .A(G2084), .B(KEYINPUT54), .ZN(n979) );
  XNOR2_X1 U1080 ( .A(n980), .B(n979), .ZN(n981) );
  NAND2_X1 U1081 ( .A1(n982), .A2(n981), .ZN(n985) );
  XNOR2_X1 U1082 ( .A(KEYINPUT114), .B(G2090), .ZN(n983) );
  XNOR2_X1 U1083 ( .A(G35), .B(n983), .ZN(n984) );
  NOR2_X1 U1084 ( .A1(n985), .A2(n984), .ZN(n986) );
  XOR2_X1 U1085 ( .A(KEYINPUT119), .B(n986), .Z(n987) );
  NOR2_X1 U1086 ( .A1(G29), .A2(n987), .ZN(n988) );
  XNOR2_X1 U1087 ( .A(KEYINPUT55), .B(n988), .ZN(n989) );
  NAND2_X1 U1088 ( .A1(n989), .A2(G11), .ZN(n1041) );
  NAND2_X1 U1089 ( .A1(n991), .A2(n990), .ZN(n997) );
  XOR2_X1 U1090 ( .A(G2072), .B(n992), .Z(n994) );
  XOR2_X1 U1091 ( .A(G164), .B(G2078), .Z(n993) );
  NOR2_X1 U1092 ( .A1(n994), .A2(n993), .ZN(n995) );
  XOR2_X1 U1093 ( .A(KEYINPUT50), .B(n995), .Z(n996) );
  NOR2_X1 U1094 ( .A1(n997), .A2(n996), .ZN(n1012) );
  XNOR2_X1 U1095 ( .A(G160), .B(G2084), .ZN(n999) );
  NAND2_X1 U1096 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NOR2_X1 U1097 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XOR2_X1 U1098 ( .A(KEYINPUT112), .B(n1002), .Z(n1003) );
  NOR2_X1 U1099 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1100 ( .A(KEYINPUT113), .B(n1005), .ZN(n1010) );
  XOR2_X1 U1101 ( .A(G2090), .B(G162), .Z(n1006) );
  NOR2_X1 U1102 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1103 ( .A(KEYINPUT51), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1104 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1105 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1106 ( .A(n1013), .B(KEYINPUT52), .ZN(n1014) );
  NAND2_X1 U1107 ( .A1(n1014), .A2(G29), .ZN(n1039) );
  XNOR2_X1 U1108 ( .A(KEYINPUT56), .B(G16), .ZN(n1037) );
  XNOR2_X1 U1109 ( .A(G1966), .B(G168), .ZN(n1016) );
  NAND2_X1 U1110 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1111 ( .A(n1017), .B(KEYINPUT57), .ZN(n1035) );
  XNOR2_X1 U1112 ( .A(G1341), .B(n1018), .ZN(n1019) );
  NOR2_X1 U1113 ( .A1(n1020), .A2(n1019), .ZN(n1030) );
  NAND2_X1 U1114 ( .A1(G1971), .A2(G303), .ZN(n1021) );
  NAND2_X1 U1115 ( .A1(n1022), .A2(n1021), .ZN(n1028) );
  XNOR2_X1 U1116 ( .A(G299), .B(G1956), .ZN(n1024) );
  XNOR2_X1 U1117 ( .A(G301), .B(G1961), .ZN(n1023) );
  NOR2_X1 U1118 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1119 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1120 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1121 ( .A1(n1030), .A2(n1029), .ZN(n1033) );
  XNOR2_X1 U1122 ( .A(G1348), .B(n1031), .ZN(n1032) );
  NOR2_X1 U1123 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NAND2_X1 U1124 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NAND2_X1 U1125 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  NAND2_X1 U1126 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  NOR2_X1 U1127 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  NAND2_X1 U1128 ( .A1(n1043), .A2(n1042), .ZN(n1044) );
  XOR2_X1 U1129 ( .A(KEYINPUT62), .B(n1044), .Z(G311) );
  INV_X1 U1130 ( .A(G311), .ZN(G150) );
endmodule

