//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 0 0 0 0 0 0 0 1 0 1 0 0 1 0 1 0 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 1 0 0 0 0 0 0 0 1 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:45 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n209, new_n210, new_n211, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n247, new_n248, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n258, new_n259, new_n260,
    new_n261, new_n262, new_n263, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1188,
    new_n1189, new_n1191, new_n1192, new_n1193, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1252, new_n1253, new_n1254;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NOR3_X1   g0007(.A1(new_n207), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0008(.A(G97), .ZN(new_n209));
  INV_X1    g0009(.A(G107), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(G87), .ZN(G355));
  INV_X1    g0012(.A(G50), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n206), .A2(new_n213), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT67), .Z(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(KEYINPUT66), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT66), .ZN(new_n218));
  NAND3_X1  g0018(.A1(new_n218), .A2(G1), .A3(G13), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n215), .A2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(KEYINPUT1), .ZN(new_n225));
  INV_X1    g0025(.A(G1), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n226), .A2(new_n222), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT68), .Z(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  INV_X1    g0030(.A(G238), .ZN(new_n231));
  OAI22_X1  g0031(.A1(new_n201), .A2(new_n230), .B1(new_n202), .B2(new_n231), .ZN(new_n232));
  INV_X1    g0032(.A(G77), .ZN(new_n233));
  INV_X1    g0033(.A(G244), .ZN(new_n234));
  INV_X1    g0034(.A(G87), .ZN(new_n235));
  INV_X1    g0035(.A(G250), .ZN(new_n236));
  OAI22_X1  g0036(.A1(new_n233), .A2(new_n234), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g0037(.A(G257), .ZN(new_n238));
  INV_X1    g0038(.A(G264), .ZN(new_n239));
  OAI22_X1  g0039(.A1(new_n209), .A2(new_n238), .B1(new_n210), .B2(new_n239), .ZN(new_n240));
  NOR3_X1   g0040(.A1(new_n232), .A2(new_n237), .A3(new_n240), .ZN(new_n241));
  AOI21_X1  g0041(.A(new_n227), .B1(new_n229), .B2(new_n241), .ZN(new_n242));
  OAI21_X1  g0042(.A(new_n224), .B1(new_n225), .B2(new_n242), .ZN(new_n243));
  INV_X1    g0043(.A(G13), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n227), .A2(new_n244), .ZN(new_n245));
  AOI211_X1 g0045(.A(new_n236), .B(new_n245), .C1(new_n238), .C2(new_n239), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT65), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT0), .ZN(new_n248));
  AOI211_X1 g0048(.A(new_n243), .B(new_n248), .C1(new_n225), .C2(new_n242), .ZN(G361));
  XNOR2_X1  g0049(.A(G238), .B(G244), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(new_n230), .ZN(new_n251));
  XOR2_X1   g0051(.A(KEYINPUT2), .B(G226), .Z(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(G250), .B(G257), .ZN(new_n254));
  XNOR2_X1  g0054(.A(G264), .B(G270), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XOR2_X1   g0056(.A(new_n253), .B(new_n256), .Z(G358));
  XNOR2_X1  g0057(.A(G50), .B(G68), .ZN(new_n258));
  XNOR2_X1  g0058(.A(G58), .B(G77), .ZN(new_n259));
  XOR2_X1   g0059(.A(new_n258), .B(new_n259), .Z(new_n260));
  XOR2_X1   g0060(.A(G87), .B(G97), .Z(new_n261));
  XOR2_X1   g0061(.A(G107), .B(G116), .Z(new_n262));
  XNOR2_X1  g0062(.A(new_n261), .B(new_n262), .ZN(new_n263));
  XOR2_X1   g0063(.A(new_n260), .B(new_n263), .Z(G351));
  INV_X1    g0064(.A(KEYINPUT69), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n226), .B1(G41), .B2(G45), .ZN(new_n266));
  INV_X1    g0066(.A(G274), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G41), .ZN(new_n269));
  INV_X1    g0069(.A(G45), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND4_X1  g0071(.A1(new_n271), .A2(KEYINPUT69), .A3(new_n226), .A4(G274), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G33), .A2(G41), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n275), .A2(G1), .A3(G13), .ZN(new_n276));
  AND2_X1   g0076(.A1(new_n276), .A2(new_n266), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n274), .B1(G226), .B2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT3), .ZN(new_n279));
  INV_X1    g0079(.A(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G1698), .ZN(new_n284));
  INV_X1    g0084(.A(G223), .ZN(new_n285));
  OAI22_X1  g0085(.A1(new_n284), .A2(new_n285), .B1(new_n233), .B2(new_n283), .ZN(new_n286));
  AND2_X1   g0086(.A1(KEYINPUT3), .A2(G33), .ZN(new_n287));
  NOR2_X1   g0087(.A1(KEYINPUT3), .A2(G33), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n289), .A2(G1698), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n286), .B1(G222), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n220), .A2(new_n275), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n278), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G169), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n226), .A2(G20), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n217), .A2(new_n219), .A3(new_n296), .A4(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G50), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n244), .A2(G1), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G20), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n299), .B1(G50), .B2(new_n302), .ZN(new_n303));
  XOR2_X1   g0103(.A(new_n303), .B(KEYINPUT70), .Z(new_n304));
  NAND3_X1  g0104(.A1(new_n217), .A2(new_n219), .A3(new_n296), .ZN(new_n305));
  XOR2_X1   g0105(.A(KEYINPUT8), .B(G58), .Z(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n280), .A2(G20), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G150), .ZN(new_n310));
  NOR2_X1   g0110(.A1(G20), .A2(G33), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  OAI22_X1  g0112(.A1(new_n307), .A2(new_n309), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n222), .B1(new_n206), .B2(new_n213), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n305), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n304), .A2(new_n315), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n295), .B(new_n316), .C1(G179), .C2(new_n293), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G190), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n293), .A2(new_n319), .ZN(new_n320));
  AOI211_X1 g0120(.A(KEYINPUT72), .B(new_n320), .C1(G200), .C2(new_n293), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT9), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n316), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n304), .A2(KEYINPUT9), .A3(new_n315), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n321), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  OR2_X1    g0125(.A1(new_n325), .A2(KEYINPUT10), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(KEYINPUT10), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n318), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n307), .A2(new_n301), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n298), .A2(new_n306), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n332), .A2(KEYINPUT77), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT77), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n334), .B1(new_n330), .B2(new_n331), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT76), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT7), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n281), .A2(new_n338), .A3(new_n222), .A4(new_n282), .ZN(new_n339));
  NOR3_X1   g0139(.A1(new_n287), .A2(new_n288), .A3(G20), .ZN(new_n340));
  XNOR2_X1  g0140(.A(KEYINPUT75), .B(KEYINPUT7), .ZN(new_n341));
  OAI211_X1 g0141(.A(G68), .B(new_n339), .C1(new_n340), .C2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(G58), .A2(G68), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n203), .A2(new_n205), .A3(new_n343), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n344), .A2(G20), .B1(G159), .B2(new_n311), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT16), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n337), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  AOI211_X1 g0148(.A(KEYINPUT76), .B(KEYINPUT16), .C1(new_n342), .C2(new_n345), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AND2_X1   g0150(.A1(new_n340), .A2(new_n341), .ZN(new_n351));
  OAI21_X1  g0151(.A(G68), .B1(new_n340), .B2(new_n338), .ZN(new_n352));
  OAI211_X1 g0152(.A(KEYINPUT16), .B(new_n345), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  AND2_X1   g0153(.A1(new_n353), .A2(new_n305), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n336), .B1(new_n350), .B2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT79), .ZN(new_n356));
  AND3_X1   g0156(.A1(new_n276), .A2(G232), .A3(new_n266), .ZN(new_n357));
  INV_X1    g0157(.A(G1698), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n285), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G226), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(G1698), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n359), .B(new_n361), .C1(new_n287), .C2(new_n288), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n280), .A2(new_n235), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n217), .A2(new_n219), .B1(G33), .B2(G41), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n357), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT78), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n367), .A2(new_n368), .A3(new_n319), .A4(new_n273), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n276), .A2(G232), .A3(new_n266), .ZN(new_n370));
  NOR2_X1   g0170(.A1(G223), .A2(G1698), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n371), .B1(new_n360), .B2(G1698), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n363), .B1(new_n372), .B2(new_n283), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n273), .B(new_n370), .C1(new_n373), .C2(new_n292), .ZN(new_n374));
  INV_X1    g0174(.A(G200), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AND2_X1   g0176(.A1(new_n369), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT78), .B1(new_n374), .B2(G190), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n356), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n378), .A2(new_n356), .A3(new_n369), .A4(new_n376), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n355), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT17), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n346), .A2(new_n347), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(KEYINPUT76), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n346), .A2(new_n337), .A3(new_n347), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n354), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n336), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n374), .A2(G169), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n367), .A2(G179), .A3(new_n273), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(KEYINPUT18), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT18), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n390), .A2(new_n396), .A3(new_n393), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n378), .A2(new_n369), .A3(new_n376), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(KEYINPUT79), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n380), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n400), .A2(KEYINPUT17), .A3(new_n355), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n384), .A2(new_n395), .A3(new_n397), .A4(new_n401), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n311), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(new_n309), .B2(new_n233), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n305), .ZN(new_n405));
  XOR2_X1   g0205(.A(new_n405), .B(KEYINPUT11), .Z(new_n406));
  NOR2_X1   g0206(.A1(new_n222), .A2(G68), .ZN(new_n407));
  AOI21_X1  g0207(.A(KEYINPUT74), .B1(new_n300), .B2(new_n407), .ZN(new_n408));
  XNOR2_X1  g0208(.A(new_n408), .B(KEYINPUT12), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n409), .B1(new_n202), .B2(new_n298), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n406), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n283), .A2(G232), .A3(G1698), .ZN(new_n413));
  NAND2_X1  g0213(.A1(G33), .A2(G97), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n283), .A2(new_n358), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n413), .B(new_n414), .C1(new_n415), .C2(new_n360), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n366), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n231), .B1(new_n277), .B2(KEYINPUT73), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(KEYINPUT73), .B2(new_n277), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n417), .A2(new_n419), .A3(new_n273), .ZN(new_n420));
  OR2_X1    g0220(.A1(new_n420), .A2(KEYINPUT13), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(KEYINPUT13), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n294), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT14), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n421), .A2(new_n422), .ZN(new_n425));
  INV_X1    g0225(.A(G179), .ZN(new_n426));
  OAI22_X1  g0226(.A1(new_n423), .A2(new_n424), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n423), .A2(new_n424), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n412), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n425), .A2(G200), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n430), .B(new_n411), .C1(new_n319), .C2(new_n425), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  XNOR2_X1  g0233(.A(KEYINPUT15), .B(G87), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n435), .A2(new_n308), .B1(G20), .B2(G77), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n436), .B1(new_n307), .B2(new_n312), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n437), .A2(new_n305), .B1(new_n233), .B2(new_n302), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n298), .A2(new_n233), .ZN(new_n439));
  XNOR2_X1  g0239(.A(new_n439), .B(KEYINPUT71), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n283), .A2(G232), .A3(new_n358), .ZN(new_n442));
  OAI221_X1 g0242(.A(new_n442), .B1(new_n210), .B2(new_n283), .C1(new_n284), .C2(new_n231), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(new_n366), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n274), .B1(G244), .B2(new_n277), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n441), .B1(G200), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n447), .B1(new_n319), .B2(new_n446), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n446), .A2(new_n294), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n444), .A2(new_n426), .A3(new_n445), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n449), .A2(new_n441), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  NOR4_X1   g0252(.A1(new_n329), .A2(new_n402), .A3(new_n433), .A4(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT83), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT19), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n222), .B1(new_n414), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n456), .B1(G87), .B2(new_n211), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n283), .A2(new_n222), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n457), .B1(new_n458), .B2(new_n202), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n222), .A2(G33), .A3(G97), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT82), .ZN(new_n461));
  AND3_X1   g0261(.A1(new_n460), .A2(new_n461), .A3(new_n455), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n461), .B1(new_n460), .B2(new_n455), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n305), .B1(new_n459), .B2(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n435), .A2(new_n301), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n305), .ZN(new_n468));
  AOI22_X1  g0268(.A1(new_n300), .A2(G20), .B1(new_n226), .B2(G33), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n465), .B(new_n467), .C1(new_n235), .C2(new_n470), .ZN(new_n471));
  OAI211_X1 g0271(.A(G244), .B(G1698), .C1(new_n287), .C2(new_n288), .ZN(new_n472));
  OAI211_X1 g0272(.A(G238), .B(new_n358), .C1(new_n287), .C2(new_n288), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G33), .A2(G116), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n366), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n226), .A2(G45), .A3(G274), .ZN(new_n477));
  INV_X1    g0277(.A(new_n276), .ZN(new_n478));
  OAI21_X1  g0278(.A(G250), .B1(new_n270), .B2(G1), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n476), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n482), .A2(new_n319), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n480), .B1(new_n475), .B2(new_n366), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n484), .A2(new_n375), .ZN(new_n485));
  NOR3_X1   g0285(.A1(new_n471), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n470), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n435), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n488), .A2(new_n465), .A3(new_n467), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n476), .A2(new_n426), .A3(new_n481), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(KEYINPUT80), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT80), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n484), .A2(new_n493), .A3(new_n426), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n482), .A2(new_n294), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n492), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT81), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n490), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n492), .A2(new_n495), .A3(KEYINPUT81), .A4(new_n494), .ZN(new_n499));
  AOI211_X1 g0299(.A(new_n454), .B(new_n486), .C1(new_n498), .C2(new_n499), .ZN(new_n500));
  OAI22_X1  g0300(.A1(new_n491), .A2(KEYINPUT80), .B1(G169), .B2(new_n484), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n493), .B1(new_n484), .B2(new_n426), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n497), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n503), .A2(new_n499), .A3(new_n489), .ZN(new_n504));
  OR3_X1    g0304(.A1(new_n471), .A2(new_n483), .A3(new_n485), .ZN(new_n505));
  AOI21_X1  g0305(.A(KEYINPUT83), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n500), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g0307(.A(KEYINPUT5), .B(G41), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n270), .A2(G1), .ZN(new_n509));
  INV_X1    g0309(.A(new_n216), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n508), .A2(new_n509), .B1(new_n510), .B2(new_n275), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n477), .B1(new_n510), .B2(new_n275), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n511), .A2(G270), .B1(new_n508), .B2(new_n512), .ZN(new_n513));
  OAI211_X1 g0313(.A(G264), .B(G1698), .C1(new_n287), .C2(new_n288), .ZN(new_n514));
  OAI211_X1 g0314(.A(G257), .B(new_n358), .C1(new_n287), .C2(new_n288), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n281), .A2(G303), .A3(new_n282), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n366), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n294), .B1(new_n513), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n468), .A2(G116), .A3(new_n469), .ZN(new_n520));
  INV_X1    g0320(.A(G116), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n300), .A2(G20), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(G20), .B1(G33), .B2(G283), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n280), .A2(G97), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n523), .A2(new_n524), .B1(G20), .B2(new_n521), .ZN(new_n525));
  AND3_X1   g0325(.A1(new_n525), .A2(new_n305), .A3(KEYINPUT20), .ZN(new_n526));
  AOI21_X1  g0326(.A(KEYINPUT20), .B1(new_n525), .B2(new_n305), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n520), .B(new_n522), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  AND3_X1   g0328(.A1(new_n519), .A2(KEYINPUT21), .A3(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n528), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n513), .A2(new_n518), .A3(G179), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(KEYINPUT21), .B1(new_n519), .B2(new_n528), .ZN(new_n533));
  NOR3_X1   g0333(.A1(new_n529), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  OAI211_X1 g0334(.A(G107), .B(new_n339), .C1(new_n340), .C2(new_n341), .ZN(new_n535));
  NAND2_X1  g0335(.A1(G97), .A2(G107), .ZN(new_n536));
  AOI21_X1  g0336(.A(KEYINPUT6), .B1(new_n211), .B2(new_n536), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n210), .A2(KEYINPUT6), .A3(G97), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OAI221_X1 g0339(.A(new_n535), .B1(new_n233), .B2(new_n312), .C1(new_n222), .C2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n305), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n301), .A2(G97), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n543), .B1(new_n470), .B2(new_n209), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n541), .A2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT4), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n547), .B1(new_n415), .B2(new_n234), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n290), .A2(KEYINPUT4), .A3(G244), .ZN(new_n549));
  NAND2_X1  g0349(.A1(G33), .A2(G283), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n283), .A2(G250), .A3(G1698), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n548), .A2(new_n549), .A3(new_n550), .A4(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n366), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n511), .A2(G257), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n512), .A2(new_n508), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n553), .A2(new_n426), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n556), .B1(new_n552), .B2(new_n366), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n546), .B(new_n558), .C1(G169), .C2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n553), .A2(G190), .A3(new_n557), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n544), .B1(new_n540), .B2(new_n305), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n561), .B(new_n562), .C1(new_n375), .C2(new_n559), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n513), .A2(new_n518), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n528), .B1(new_n564), .B2(G200), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n319), .B2(new_n564), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n534), .A2(new_n560), .A3(new_n563), .A4(new_n566), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n222), .B(G87), .C1(new_n287), .C2(new_n288), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(KEYINPUT22), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT22), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n283), .A2(new_n570), .A3(new_n222), .A4(G87), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT24), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n474), .A2(G20), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT23), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n222), .B2(G107), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n210), .A2(KEYINPUT23), .A3(G20), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n574), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n572), .A2(new_n573), .A3(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n573), .B1(new_n572), .B2(new_n578), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n305), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n283), .A2(G250), .A3(new_n358), .ZN(new_n583));
  OAI211_X1 g0383(.A(G257), .B(G1698), .C1(new_n287), .C2(new_n288), .ZN(new_n584));
  NAND2_X1  g0384(.A1(G33), .A2(G294), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n366), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n511), .A2(G264), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n587), .A2(new_n588), .A3(new_n555), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(G200), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT25), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n591), .B1(new_n301), .B2(G107), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n302), .A2(KEYINPUT25), .A3(new_n210), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n487), .A2(G107), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n586), .A2(new_n366), .B1(G264), .B2(new_n511), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n595), .A2(G190), .A3(new_n555), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n582), .A2(new_n590), .A3(new_n594), .A4(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT84), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n595), .A2(new_n598), .A3(G179), .A4(new_n555), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n572), .A2(new_n578), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(KEYINPUT24), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n468), .B1(new_n601), .B2(new_n579), .ZN(new_n602));
  INV_X1    g0402(.A(new_n594), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n599), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(KEYINPUT84), .B1(new_n589), .B2(new_n426), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n294), .B1(new_n595), .B2(new_n555), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n597), .B1(new_n604), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(KEYINPUT85), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n582), .A2(new_n594), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n610), .B(new_n599), .C1(new_n606), .C2(new_n605), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT85), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n611), .A2(new_n612), .A3(new_n597), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n567), .B1(new_n609), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n453), .A2(new_n507), .A3(new_n614), .ZN(new_n615));
  XOR2_X1   g0415(.A(new_n615), .B(KEYINPUT86), .Z(G372));
  AND2_X1   g0416(.A1(new_n429), .A2(new_n451), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n431), .A2(new_n384), .A3(new_n401), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n395), .B(new_n397), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n326), .A2(new_n327), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n318), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n453), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT26), .ZN(new_n623));
  INV_X1    g0423(.A(new_n560), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n623), .B1(new_n507), .B2(new_n624), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n495), .A2(new_n491), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n489), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n505), .A2(new_n627), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n629), .A2(new_n560), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n628), .B1(new_n630), .B2(new_n623), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n611), .A2(new_n534), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n560), .A2(new_n563), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n505), .A2(new_n627), .A3(new_n597), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n631), .B1(new_n633), .B2(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n625), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n621), .B1(new_n622), .B2(new_n638), .ZN(G369));
  INV_X1    g0439(.A(new_n300), .ZN(new_n640));
  OR3_X1    g0440(.A1(new_n640), .A2(KEYINPUT27), .A3(G20), .ZN(new_n641));
  OAI21_X1  g0441(.A(KEYINPUT27), .B1(new_n640), .B2(G20), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n641), .A2(G213), .A3(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(G343), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n611), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n609), .A2(new_n613), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n534), .A2(new_n645), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n645), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n611), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n610), .A2(new_n645), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n651), .B1(new_n647), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n645), .A2(new_n528), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n534), .A2(new_n566), .A3(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n655), .B1(new_n534), .B2(new_n654), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(G330), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n649), .B1(new_n653), .B2(new_n657), .ZN(new_n658));
  XNOR2_X1  g0458(.A(new_n658), .B(KEYINPUT87), .ZN(G399));
  NOR2_X1   g0459(.A1(new_n245), .A2(G41), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NOR3_X1   g0461(.A1(new_n211), .A2(G87), .A3(G116), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(G1), .A3(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n214), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n663), .B1(new_n664), .B2(new_n661), .ZN(new_n665));
  XNOR2_X1  g0465(.A(new_n665), .B(KEYINPUT28), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT31), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n614), .A2(new_n507), .A3(new_n650), .ZN(new_n668));
  INV_X1    g0468(.A(new_n559), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n484), .A2(G179), .ZN(new_n670));
  AND4_X1   g0470(.A1(new_n589), .A2(new_n669), .A3(new_n564), .A4(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n531), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n672), .A2(new_n484), .A3(new_n595), .ZN(new_n673));
  OAI21_X1  g0473(.A(KEYINPUT88), .B1(new_n673), .B2(new_n669), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n671), .B1(KEYINPUT30), .B2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n675), .B1(KEYINPUT30), .B2(new_n674), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n645), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n667), .B1(new_n668), .B2(new_n677), .ZN(new_n678));
  AOI21_X1  g0478(.A(KEYINPUT31), .B1(new_n676), .B2(new_n645), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(G330), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT90), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n636), .B2(new_n633), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n632), .A2(new_n634), .A3(new_n635), .A4(KEYINPUT90), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n628), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n504), .A2(new_n505), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n454), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n504), .A2(KEYINPUT83), .A3(new_n505), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n688), .A2(new_n689), .A3(new_n624), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n690), .A2(KEYINPUT89), .A3(new_n623), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n630), .A2(KEYINPUT26), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(KEYINPUT89), .B1(new_n690), .B2(new_n623), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n686), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n695), .A2(KEYINPUT29), .A3(new_n650), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n638), .A2(new_n645), .ZN(new_n697));
  OR2_X1    g0497(.A1(new_n697), .A2(KEYINPUT29), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n682), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n666), .B1(new_n699), .B2(G1), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT91), .ZN(G364));
  NOR2_X1   g0501(.A1(new_n244), .A2(G20), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n226), .B1(new_n702), .B2(G45), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n660), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n245), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(G116), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n245), .A2(new_n283), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(new_n260), .B2(new_n270), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n709), .B1(new_n270), .B2(new_n215), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n245), .A2(new_n289), .ZN(new_n711));
  AOI211_X1 g0511(.A(new_n707), .B(new_n710), .C1(G355), .C2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(G13), .A2(G33), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(G20), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n715), .B(KEYINPUT92), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n221), .B1(G20), .B2(new_n294), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n705), .B1(new_n712), .B2(new_n720), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n721), .A2(KEYINPUT93), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n222), .A2(new_n319), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n723), .A2(new_n426), .A3(G200), .ZN(new_n724));
  INV_X1    g0524(.A(G303), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n426), .A2(new_n375), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(new_n723), .ZN(new_n727));
  INV_X1    g0527(.A(G326), .ZN(new_n728));
  OAI22_X1  g0528(.A1(new_n724), .A2(new_n725), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(G179), .A2(G200), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n222), .B1(new_n730), .B2(G190), .ZN(new_n731));
  INV_X1    g0531(.A(G294), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n222), .A2(G190), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n734), .A2(G179), .A3(new_n375), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(G283), .ZN(new_n737));
  OAI221_X1 g0537(.A(new_n289), .B1(new_n731), .B2(new_n732), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n733), .A2(new_n730), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  AOI211_X1 g0540(.A(new_n729), .B(new_n738), .C1(G329), .C2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(G311), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n426), .A2(G200), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT94), .ZN(new_n744));
  AND3_X1   g0544(.A1(new_n733), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n744), .B1(new_n733), .B2(new_n743), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n741), .B1(new_n742), .B2(new_n747), .ZN(new_n748));
  XOR2_X1   g0548(.A(KEYINPUT33), .B(G317), .Z(new_n749));
  NAND2_X1  g0549(.A1(new_n726), .A2(new_n733), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n723), .A2(new_n743), .ZN(new_n751));
  INV_X1    g0551(.A(G322), .ZN(new_n752));
  OAI22_X1  g0552(.A1(new_n749), .A2(new_n750), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT96), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n736), .A2(new_n210), .ZN(new_n755));
  INV_X1    g0555(.A(new_n751), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n755), .B1(G58), .B2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n731), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G97), .ZN(new_n759));
  INV_X1    g0559(.A(new_n727), .ZN(new_n760));
  INV_X1    g0560(.A(new_n750), .ZN(new_n761));
  AOI22_X1  g0561(.A1(G50), .A2(new_n760), .B1(new_n761), .B2(G68), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n757), .A2(new_n759), .A3(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT32), .ZN(new_n764));
  INV_X1    g0564(.A(G159), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n764), .B1(new_n739), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n740), .A2(KEYINPUT32), .A3(G159), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n283), .B1(new_n724), .B2(new_n235), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n766), .A2(new_n767), .B1(new_n768), .B2(KEYINPUT95), .ZN(new_n769));
  INV_X1    g0569(.A(new_n747), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G77), .ZN(new_n771));
  OR2_X1    g0571(.A1(new_n768), .A2(KEYINPUT95), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n769), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  OAI22_X1  g0573(.A1(new_n748), .A2(new_n754), .B1(new_n763), .B2(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n722), .B1(new_n718), .B2(new_n774), .ZN(new_n775));
  OAI221_X1 g0575(.A(new_n775), .B1(KEYINPUT93), .B2(new_n721), .C1(new_n656), .C2(new_n716), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n705), .B1(new_n656), .B2(G330), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(G330), .B2(new_n656), .ZN(new_n778));
  AND2_X1   g0578(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(G396));
  NOR2_X1   g0580(.A1(new_n451), .A2(new_n645), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n441), .A2(new_n645), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n448), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n781), .B1(new_n783), .B2(new_n451), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n697), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(KEYINPUT100), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n697), .A2(new_n784), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(new_n682), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n705), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n791), .B1(new_n788), .B2(new_n682), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n784), .A2(new_n714), .ZN(new_n793));
  INV_X1    g0593(.A(new_n718), .ZN(new_n794));
  AOI22_X1  g0594(.A1(G137), .A2(new_n760), .B1(new_n756), .B2(G143), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n795), .B1(new_n310), .B2(new_n750), .C1(new_n747), .C2(new_n765), .ZN(new_n796));
  INV_X1    g0596(.A(KEYINPUT34), .ZN(new_n797));
  AND2_X1   g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n736), .A2(new_n202), .ZN(new_n799));
  INV_X1    g0599(.A(new_n724), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n799), .B1(G50), .B2(new_n800), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n801), .B1(new_n201), .B2(new_n731), .ZN(new_n802));
  INV_X1    g0602(.A(G132), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n283), .B1(new_n739), .B2(new_n803), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT98), .ZN(new_n805));
  NOR3_X1   g0605(.A1(new_n798), .A2(new_n802), .A3(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n806), .B1(new_n797), .B2(new_n796), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n751), .A2(new_n732), .B1(new_n750), .B2(new_n737), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n759), .B1(new_n725), .B2(new_n727), .C1(new_n742), .C2(new_n739), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n808), .B(new_n809), .C1(G87), .C2(new_n735), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n289), .B1(new_n724), .B2(new_n210), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT97), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n810), .B(new_n812), .C1(new_n521), .C2(new_n747), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n794), .B1(new_n807), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n718), .A2(new_n713), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n791), .B(new_n814), .C1(new_n233), .C2(new_n815), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT99), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n790), .A2(new_n792), .B1(new_n793), .B2(new_n817), .ZN(G384));
  INV_X1    g0618(.A(new_n539), .ZN(new_n819));
  OR2_X1    g0619(.A1(new_n819), .A2(KEYINPUT35), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(KEYINPUT35), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n820), .A2(G116), .A3(new_n223), .A4(new_n821), .ZN(new_n822));
  XOR2_X1   g0622(.A(new_n822), .B(KEYINPUT36), .Z(new_n823));
  NAND3_X1  g0623(.A1(new_n214), .A2(G77), .A3(new_n343), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n213), .A2(G68), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n226), .B(G13), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n382), .ZN(new_n828));
  INV_X1    g0628(.A(new_n354), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n345), .B1(new_n351), .B2(new_n352), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n830), .A2(new_n347), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n332), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n391), .A2(new_n392), .A3(new_n643), .ZN(new_n833));
  AND2_X1   g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(KEYINPUT37), .B1(new_n828), .B2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n833), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(new_n388), .B2(new_n389), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n837), .B1(new_n355), .B2(new_n400), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT37), .ZN(new_n839));
  AOI21_X1  g0639(.A(KEYINPUT101), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n390), .A2(new_n833), .ZN(new_n841));
  AND4_X1   g0641(.A1(KEYINPUT101), .A2(new_n382), .A3(new_n839), .A4(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n835), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n643), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n402), .A2(new_n844), .A3(new_n832), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n843), .A2(new_n845), .A3(KEYINPUT38), .ZN(new_n846));
  AOI21_X1  g0646(.A(KEYINPUT38), .B1(new_n843), .B2(new_n845), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n846), .B1(new_n847), .B2(KEYINPUT102), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT102), .ZN(new_n849));
  AOI211_X1 g0649(.A(new_n849), .B(KEYINPUT38), .C1(new_n843), .C2(new_n845), .ZN(new_n850));
  OAI21_X1  g0650(.A(KEYINPUT39), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n402), .A2(new_n390), .A3(new_n844), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT103), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n402), .A2(KEYINPUT103), .A3(new_n390), .A4(new_n844), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT101), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n382), .A2(new_n841), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n856), .B1(new_n857), .B2(KEYINPUT37), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n838), .A2(KEYINPUT101), .A3(new_n839), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n857), .A2(KEYINPUT37), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n854), .A2(new_n855), .A3(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT38), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT39), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n865), .A2(new_n866), .A3(new_n846), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n851), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(KEYINPUT104), .ZN(new_n869));
  INV_X1    g0669(.A(new_n429), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n650), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT104), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n851), .A2(new_n867), .A3(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n869), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n848), .A2(new_n850), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n781), .B1(new_n697), .B2(new_n784), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n411), .A2(new_n650), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n429), .A2(new_n431), .A3(new_n879), .ZN(new_n880));
  OR2_X1    g0680(.A1(new_n427), .A2(new_n428), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n880), .B1(new_n882), .B2(new_n879), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NOR3_X1   g0684(.A1(new_n876), .A2(new_n877), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n844), .B1(new_n395), .B2(new_n397), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n875), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n453), .A2(new_n698), .A3(new_n696), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n621), .ZN(new_n890));
  XOR2_X1   g0690(.A(new_n888), .B(new_n890), .Z(new_n891));
  INV_X1    g0691(.A(KEYINPUT40), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n784), .B(new_n883), .C1(new_n678), .C2(new_n679), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n892), .B1(new_n876), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT105), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n892), .B1(new_n865), .B2(new_n846), .ZN(new_n896));
  INV_X1    g0696(.A(new_n893), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n843), .A2(KEYINPUT38), .A3(new_n845), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n899), .B1(new_n863), .B2(new_n864), .ZN(new_n900));
  NOR4_X1   g0700(.A1(new_n900), .A2(new_n893), .A3(KEYINPUT105), .A4(new_n892), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n894), .B1(new_n898), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n453), .A2(new_n680), .ZN(new_n903));
  OAI21_X1  g0703(.A(G330), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(new_n903), .B2(new_n902), .ZN(new_n905));
  OAI22_X1  g0705(.A1(new_n891), .A2(new_n905), .B1(new_n226), .B2(new_n702), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n891), .A2(new_n905), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n827), .B1(new_n906), .B2(new_n907), .ZN(G367));
  NOR2_X1   g0708(.A1(new_n653), .A2(new_n657), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n634), .B1(new_n562), .B2(new_n650), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n624), .A2(new_n645), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n471), .A2(new_n645), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n505), .A2(new_n627), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n627), .B2(new_n914), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n916), .A2(KEYINPUT43), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n917), .B(KEYINPUT106), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n913), .B(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n916), .A2(KEYINPUT43), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n912), .A2(new_n647), .A3(new_n648), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(KEYINPUT42), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n560), .B1(new_n910), .B2(new_n611), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n650), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n921), .A2(KEYINPUT42), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n920), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n919), .B(new_n927), .ZN(new_n928));
  XOR2_X1   g0728(.A(new_n660), .B(KEYINPUT41), .Z(new_n929));
  MUX2_X1   g0729(.A(new_n653), .B(new_n647), .S(new_n648), .Z(new_n930));
  XOR2_X1   g0730(.A(new_n930), .B(new_n657), .Z(new_n931));
  NAND2_X1  g0731(.A1(new_n699), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n649), .A2(new_n912), .ZN(new_n933));
  XOR2_X1   g0733(.A(new_n933), .B(KEYINPUT45), .Z(new_n934));
  NOR2_X1   g0734(.A1(new_n649), .A2(new_n912), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT44), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(new_n909), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n932), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n929), .B1(new_n939), .B2(new_n699), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT107), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n928), .B1(new_n941), .B2(new_n704), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n720), .B1(new_n245), .B2(new_n435), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n256), .A2(new_n708), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n791), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n724), .A2(new_n521), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n946), .A2(KEYINPUT46), .ZN(new_n947));
  AOI211_X1 g0747(.A(new_n283), .B(new_n947), .C1(G311), .C2(new_n760), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n946), .A2(KEYINPUT46), .B1(G107), .B2(new_n758), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n770), .A2(G283), .ZN(new_n950));
  OAI22_X1  g0750(.A1(new_n736), .A2(new_n209), .B1(new_n732), .B2(new_n750), .ZN(new_n951));
  XOR2_X1   g0751(.A(KEYINPUT108), .B(G317), .Z(new_n952));
  OAI22_X1  g0752(.A1(new_n952), .A2(new_n739), .B1(new_n751), .B2(new_n725), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NAND4_X1  g0754(.A1(new_n948), .A2(new_n949), .A3(new_n950), .A4(new_n954), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n736), .A2(new_n233), .B1(new_n765), .B2(new_n750), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n956), .B1(G137), .B2(new_n740), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n758), .A2(G68), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n751), .A2(new_n310), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n283), .B1(new_n724), .B2(new_n201), .ZN(new_n960));
  AOI211_X1 g0760(.A(new_n959), .B(new_n960), .C1(G143), .C2(new_n760), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n770), .A2(G50), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n957), .A2(new_n958), .A3(new_n961), .A4(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n955), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT110), .ZN(new_n965));
  XNOR2_X1  g0765(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n965), .B(new_n966), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n945), .B1(new_n716), .B2(new_n916), .C1(new_n967), .C2(new_n794), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n942), .A2(new_n968), .ZN(G387));
  INV_X1    g0769(.A(new_n662), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n711), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(G107), .B2(new_n706), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n306), .A2(new_n213), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n973), .B(KEYINPUT50), .Z(new_n974));
  AOI211_X1 g0774(.A(G45), .B(new_n970), .C1(G68), .C2(G77), .ZN(new_n975));
  AOI211_X1 g0775(.A(new_n245), .B(new_n283), .C1(new_n974), .C2(new_n975), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n253), .A2(new_n270), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n972), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n800), .A2(G77), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n979), .B1(new_n750), .B2(new_n307), .C1(new_n765), .C2(new_n727), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n751), .A2(new_n213), .B1(new_n739), .B2(new_n310), .ZN(new_n981));
  AOI211_X1 g0781(.A(new_n289), .B(new_n981), .C1(G97), .C2(new_n735), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n758), .A2(new_n435), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n980), .B(new_n984), .C1(G68), .C2(new_n770), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n289), .B1(new_n739), .B2(new_n728), .ZN(new_n986));
  AOI22_X1  g0786(.A1(G322), .A2(new_n760), .B1(new_n761), .B2(G311), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n751), .B2(new_n952), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n988), .B1(G303), .B2(new_n770), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n989), .A2(KEYINPUT48), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(KEYINPUT48), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n800), .A2(G294), .B1(new_n758), .B2(G283), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n990), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT49), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n986), .B(new_n995), .C1(G116), .C2(new_n735), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n993), .A2(new_n994), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n985), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n705), .B1(new_n720), .B2(new_n978), .C1(new_n998), .C2(new_n794), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(new_n653), .B2(new_n717), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(new_n931), .B2(new_n704), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n932), .A2(new_n660), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n699), .A2(new_n931), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1001), .B1(new_n1002), .B2(new_n1003), .ZN(G393));
  NAND2_X1  g0804(.A1(new_n932), .A2(new_n938), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n939), .A2(new_n660), .A3(new_n1005), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT111), .Z(new_n1007));
  OAI21_X1  g0807(.A(new_n719), .B1(new_n209), .B2(new_n706), .ZN(new_n1008));
  AND2_X1   g0808(.A1(new_n263), .A2(new_n708), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n705), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n283), .B(new_n755), .C1(G116), .C2(new_n758), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n724), .A2(new_n737), .B1(new_n739), .B2(new_n752), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(G303), .B2(new_n761), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1011), .B(new_n1013), .C1(new_n732), .C2(new_n747), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(G317), .A2(new_n760), .B1(new_n756), .B2(G311), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT52), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n731), .A2(new_n233), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n289), .B(new_n1017), .C1(G87), .C2(new_n735), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(G50), .A2(new_n761), .B1(new_n740), .B2(G143), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1018), .B(new_n1019), .C1(new_n202), .C2(new_n724), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n727), .A2(new_n310), .B1(new_n751), .B2(new_n765), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT51), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n307), .B2(new_n747), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n1014), .A2(new_n1016), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1010), .B1(new_n1024), .B2(new_n718), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n912), .B2(new_n716), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n938), .B2(new_n703), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n1007), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(G390));
  OAI211_X1 g0829(.A(G330), .B(new_n784), .C1(new_n678), .C2(new_n679), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1030), .A2(new_n884), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n900), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n871), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n783), .A2(new_n451), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n695), .A2(new_n650), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT112), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n781), .ZN(new_n1037));
  AND3_X1   g0837(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1036), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1033), .B1(new_n1040), .B2(new_n883), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n877), .A2(new_n884), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1042), .A2(new_n872), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(new_n869), .B2(new_n874), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1031), .B1(new_n1041), .B2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n900), .A2(new_n872), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(KEYINPUT112), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1046), .B1(new_n1050), .B2(new_n884), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n874), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n873), .B1(new_n851), .B2(new_n867), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n1052), .A2(new_n1053), .B1(new_n872), .B2(new_n1042), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1031), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1051), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1045), .A2(new_n1056), .A3(new_n704), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n713), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n1017), .B(new_n799), .C1(G283), .C2(new_n760), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n751), .A2(new_n521), .B1(new_n750), .B2(new_n210), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(G294), .B2(new_n740), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1059), .B(new_n1061), .C1(new_n209), .C2(new_n747), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n289), .B1(new_n724), .B2(new_n235), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT115), .Z(new_n1064));
  AOI21_X1  g0864(.A(new_n289), .B1(new_n735), .B2(G50), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT114), .Z(new_n1066));
  NOR2_X1   g0866(.A1(new_n724), .A2(new_n310), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT53), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(KEYINPUT54), .B(G143), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1066), .B(new_n1068), .C1(new_n747), .C2(new_n1069), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G128), .A2(new_n760), .B1(new_n761), .B2(G137), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(G132), .A2(new_n756), .B1(new_n740), .B2(G125), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1071), .B(new_n1072), .C1(new_n765), .C2(new_n731), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n1062), .A2(new_n1064), .B1(new_n1070), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n718), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n791), .B1(new_n815), .B2(new_n307), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1058), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1057), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(KEYINPUT116), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT116), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1057), .A2(new_n1080), .A3(new_n1077), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n889), .B(new_n621), .C1(new_n622), .C2(new_n681), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1030), .B(new_n883), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1050), .A2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1084), .A2(new_n877), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1083), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1045), .A2(new_n1056), .A3(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(KEYINPUT113), .B1(new_n1089), .B2(new_n660), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1089), .A2(KEYINPUT113), .A3(new_n660), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1088), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1045), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1056), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1092), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1091), .A2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1082), .B1(new_n1090), .B2(new_n1096), .ZN(G378));
  NAND2_X1  g0897(.A1(new_n316), .A2(new_n844), .ZN(new_n1098));
  XOR2_X1   g0898(.A(new_n1098), .B(KEYINPUT55), .Z(new_n1099));
  XNOR2_X1  g0899(.A(new_n328), .B(new_n1099), .ZN(new_n1100));
  XOR2_X1   g0900(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n1101));
  XNOR2_X1  g0901(.A(new_n1100), .B(new_n1101), .ZN(new_n1102));
  OAI211_X1 g0902(.A(G330), .B(new_n894), .C1(new_n898), .C2(new_n901), .ZN(new_n1103));
  AND3_X1   g0903(.A1(new_n1103), .A2(new_n875), .A3(new_n887), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1103), .B1(new_n875), .B2(new_n887), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1102), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1103), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n888), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1103), .A2(new_n875), .A3(new_n887), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1102), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1108), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1106), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1083), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1089), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT57), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n661), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1112), .A2(new_n1114), .A3(KEYINPUT57), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(KEYINPUT120), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT120), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1112), .A2(new_n1114), .A3(new_n1120), .A4(KEYINPUT57), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1117), .A2(new_n1119), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT119), .ZN(new_n1123));
  NOR3_X1   g0923(.A1(new_n1104), .A2(new_n1105), .A3(new_n1102), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1110), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n704), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1110), .A2(new_n713), .ZN(new_n1127));
  NOR3_X1   g0927(.A1(new_n718), .A2(G50), .A3(new_n713), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n736), .A2(new_n201), .B1(new_n739), .B2(new_n737), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n979), .A2(new_n269), .A3(new_n289), .A4(new_n958), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n727), .A2(new_n521), .B1(new_n751), .B2(new_n210), .ZN(new_n1131));
  NOR3_X1   g0931(.A1(new_n1129), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n770), .A2(new_n435), .B1(G97), .B2(new_n761), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT117), .ZN(new_n1134));
  AND2_X1   g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1132), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT58), .ZN(new_n1138));
  OR2_X1    g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n213), .B1(new_n287), .B2(G41), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n770), .A2(G137), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n758), .A2(G150), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(G128), .A2(new_n756), .B1(new_n761), .B2(G132), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1069), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n800), .A2(new_n1145), .B1(new_n760), .B2(G125), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1142), .A2(new_n1143), .A3(new_n1144), .A4(new_n1146), .ZN(new_n1147));
  OR2_X1    g0947(.A1(new_n1147), .A2(KEYINPUT59), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(KEYINPUT59), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n735), .A2(G159), .ZN(new_n1150));
  AOI211_X1 g0950(.A(G33), .B(G41), .C1(new_n740), .C2(G124), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .A4(new_n1151), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1139), .A2(new_n1140), .A3(new_n1141), .A4(new_n1152), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n791), .B(new_n1128), .C1(new_n1153), .C2(new_n718), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1127), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1123), .B1(new_n1126), .B2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n703), .B1(new_n1106), .B2(new_n1111), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1155), .ZN(new_n1158));
  NOR3_X1   g0958(.A1(new_n1157), .A2(KEYINPUT119), .A3(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1156), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1122), .A2(new_n1160), .ZN(G375));
  AOI21_X1  g0961(.A(new_n1086), .B1(new_n1050), .B2(new_n1084), .ZN(new_n1162));
  OR3_X1    g0962(.A1(new_n1162), .A2(KEYINPUT121), .A3(new_n703), .ZN(new_n1163));
  OAI21_X1  g0963(.A(KEYINPUT121), .B1(new_n1162), .B2(new_n703), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n884), .A2(new_n713), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n800), .A2(G159), .B1(new_n761), .B2(new_n1145), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1166), .B1(new_n803), .B2(new_n727), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(new_n770), .B2(G150), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n758), .A2(G50), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n289), .B1(new_n735), .B2(G58), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(G137), .A2(new_n756), .B1(new_n740), .B2(G128), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .A4(new_n1171), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n751), .A2(new_n737), .B1(new_n739), .B2(new_n725), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n283), .B(new_n1173), .C1(G77), .C2(new_n735), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n770), .A2(G107), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n724), .A2(new_n209), .B1(new_n727), .B2(new_n732), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(G116), .B2(new_n761), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1174), .A2(new_n983), .A3(new_n1175), .A4(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n794), .B1(new_n1172), .B2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n791), .B1(new_n815), .B2(new_n202), .ZN(new_n1180));
  XOR2_X1   g0980(.A(new_n1180), .B(KEYINPUT122), .Z(new_n1181));
  NOR2_X1   g0981(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n1163), .A2(new_n1164), .B1(new_n1165), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n929), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1162), .A2(new_n1083), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1092), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1183), .A2(new_n1186), .ZN(G381));
  OR4_X1    g0987(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1188));
  OR2_X1    g0988(.A1(G375), .A2(G378), .ZN(new_n1189));
  OR4_X1    g0989(.A1(G387), .A2(new_n1188), .A3(new_n1189), .A4(G381), .ZN(G407));
  NAND2_X1  g0990(.A1(new_n644), .A2(G213), .ZN(new_n1191));
  XOR2_X1   g0991(.A(new_n1191), .B(KEYINPUT123), .Z(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  OAI211_X1 g0993(.A(G407), .B(G213), .C1(new_n1189), .C2(new_n1193), .ZN(G409));
  INV_X1    g0994(.A(KEYINPUT63), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1122), .A2(new_n1160), .A3(G378), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1126), .B(new_n1155), .C1(new_n1115), .C2(new_n929), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1197), .B(new_n1082), .C1(new_n1090), .C2(new_n1096), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1196), .A2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT60), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1185), .B1(new_n1088), .B2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1162), .A2(KEYINPUT60), .A3(new_n1083), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1201), .A2(new_n660), .A3(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1183), .A2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(G384), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1183), .A2(G384), .A3(new_n1203), .ZN(new_n1207));
  AND2_X1   g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1199), .A2(new_n1191), .A3(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT124), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n1196), .A2(new_n1198), .B1(G213), .B2(new_n644), .ZN(new_n1212));
  AOI21_X1  g1012(.A(KEYINPUT124), .B1(new_n1212), .B2(new_n1208), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1195), .B1(new_n1211), .B2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT125), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(G387), .B(G390), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(G393), .B(new_n779), .ZN(new_n1218));
  OR2_X1    g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT61), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1219), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1208), .B1(G2897), .B2(new_n1192), .ZN(new_n1223));
  INV_X1    g1023(.A(G2897), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1191), .A2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1223), .B1(new_n1208), .B2(new_n1225), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1226), .A2(new_n1212), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1192), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n1228), .A2(KEYINPUT63), .A3(new_n1208), .ZN(new_n1229));
  NOR3_X1   g1029(.A1(new_n1222), .A2(new_n1227), .A3(new_n1229), .ZN(new_n1230));
  OAI211_X1 g1030(.A(KEYINPUT125), .B(new_n1195), .C1(new_n1211), .C2(new_n1213), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1216), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1220), .B1(new_n1226), .B2(new_n1228), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1208), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT62), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1199), .A2(new_n1236), .A3(new_n1193), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT127), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1228), .A2(KEYINPUT127), .A3(new_n1236), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1212), .A2(KEYINPUT124), .A3(new_n1208), .ZN(new_n1243));
  AOI21_X1  g1043(.A(KEYINPUT62), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1241), .B1(new_n1244), .B2(KEYINPUT126), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1235), .B1(new_n1211), .B2(new_n1213), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT126), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1233), .B1(new_n1245), .B2(new_n1248), .ZN(new_n1249));
  AND2_X1   g1049(.A1(new_n1219), .A2(new_n1221), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1232), .B1(new_n1249), .B2(new_n1250), .ZN(G405));
  NAND2_X1  g1051(.A1(G375), .A2(G378), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1189), .A2(new_n1252), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(new_n1253), .B(new_n1208), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(new_n1254), .B(new_n1250), .ZN(G402));
endmodule


