//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 0 1 0 0 1 0 0 1 1 0 0 1 0 0 1 1 1 0 1 0 0 1 0 1 1 1 0 0 0 0 0 0 0 1 1 1 1 1 1 1 1 0 0 1 0 1 0 1 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n797, new_n798, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n857, new_n858, new_n859, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n878, new_n879, new_n880, new_n881, new_n883, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT28), .ZN(new_n203));
  NOR2_X1   g002(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT66), .B(G183gat), .ZN(new_n205));
  AOI21_X1  g004(.A(new_n204), .B1(new_n205), .B2(KEYINPUT27), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n203), .B1(new_n206), .B2(G190gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(KEYINPUT27), .B(G183gat), .ZN(new_n208));
  INV_X1    g007(.A(G190gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n208), .A2(KEYINPUT28), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  OR2_X1    g012(.A1(new_n213), .A2(KEYINPUT26), .ZN(new_n214));
  NAND2_X1  g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n216), .B1(new_n213), .B2(KEYINPUT26), .ZN(new_n217));
  AOI22_X1  g016(.A1(new_n214), .A2(new_n217), .B1(G183gat), .B2(G190gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n211), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n212), .A2(KEYINPUT23), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n212), .B1(KEYINPUT23), .B2(new_n215), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  NAND3_X1  g021(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n223), .B1(new_n205), .B2(G190gat), .ZN(new_n224));
  AND3_X1   g023(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n225));
  AOI21_X1  g024(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n226));
  NOR3_X1   g025(.A1(new_n225), .A2(new_n226), .A3(KEYINPUT24), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n220), .B(new_n222), .C1(new_n224), .C2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT25), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT64), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n229), .B1(new_n220), .B2(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(KEYINPUT64), .B1(new_n212), .B2(KEYINPUT23), .ZN(new_n232));
  NOR3_X1   g031(.A1(new_n231), .A2(new_n221), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G183gat), .A2(G190gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT24), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n236), .B(new_n223), .C1(G183gat), .C2(G190gat), .ZN(new_n237));
  AOI22_X1  g036(.A1(new_n228), .A2(KEYINPUT25), .B1(new_n233), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n219), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT67), .ZN(new_n240));
  NAND2_X1  g039(.A1(G113gat), .A2(G120gat), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NOR2_X1   g041(.A1(G113gat), .A2(G120gat), .ZN(new_n243));
  NOR3_X1   g042(.A1(new_n242), .A2(new_n243), .A3(KEYINPUT1), .ZN(new_n244));
  XNOR2_X1  g043(.A(G127gat), .B(G134gat), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n240), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n243), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n247), .A2(KEYINPUT68), .A3(new_n241), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n249), .B1(new_n242), .B2(new_n243), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT1), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n248), .A2(new_n250), .A3(new_n251), .A4(new_n245), .ZN(new_n252));
  INV_X1    g051(.A(new_n245), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n247), .A2(new_n251), .A3(new_n241), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n253), .A2(new_n254), .A3(KEYINPUT67), .ZN(new_n255));
  AND3_X1   g054(.A1(new_n246), .A2(new_n252), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(G227gat), .ZN(new_n258));
  INV_X1    g057(.A(G233gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n246), .A2(new_n252), .A3(new_n255), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n219), .A2(new_n238), .A3(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n257), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n263), .A2(KEYINPUT32), .ZN(new_n264));
  XNOR2_X1  g063(.A(G15gat), .B(G43gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(G71gat), .B(G99gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  OR2_X1    g066(.A1(new_n267), .A2(KEYINPUT69), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(KEYINPUT69), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n268), .A2(KEYINPUT33), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n264), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n267), .B1(new_n263), .B2(KEYINPUT32), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT33), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n263), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n271), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT34), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n257), .A2(new_n262), .ZN(new_n278));
  INV_X1    g077(.A(new_n260), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AOI211_X1 g079(.A(KEYINPUT34), .B(new_n260), .C1(new_n257), .C2(new_n262), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n276), .A2(new_n283), .ZN(new_n284));
  AOI22_X1  g083(.A1(new_n264), .A2(new_n270), .B1(new_n272), .B2(new_n274), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(new_n282), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT29), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n239), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(G226gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n290), .A2(new_n259), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n239), .A2(new_n291), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT72), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT22), .ZN(new_n297));
  XOR2_X1   g096(.A(KEYINPUT71), .B(G211gat), .Z(new_n298));
  INV_X1    g097(.A(G218gat), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(G197gat), .B(G204gat), .ZN(new_n301));
  XNOR2_X1  g100(.A(G211gat), .B(G218gat), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n302), .B1(new_n300), .B2(new_n301), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n296), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n300), .A2(new_n301), .ZN(new_n307));
  INV_X1    g106(.A(new_n302), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n309), .A2(KEYINPUT72), .A3(new_n303), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n306), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n295), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n293), .A2(new_n311), .A3(new_n294), .ZN(new_n314));
  XNOR2_X1  g113(.A(G8gat), .B(G36gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(G64gat), .B(G92gat), .ZN(new_n316));
  XOR2_X1   g115(.A(new_n315), .B(new_n316), .Z(new_n317));
  NAND3_X1  g116(.A1(new_n313), .A2(new_n314), .A3(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT30), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n313), .A2(KEYINPUT30), .A3(new_n314), .A4(new_n317), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n313), .A2(new_n314), .ZN(new_n322));
  XOR2_X1   g121(.A(new_n317), .B(KEYINPUT73), .Z(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n320), .A2(new_n321), .A3(new_n324), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n287), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(G155gat), .A2(G162gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT2), .ZN(new_n328));
  INV_X1    g127(.A(G148gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n329), .A2(G141gat), .ZN(new_n330));
  INV_X1    g129(.A(G141gat), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n331), .A2(G148gat), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n328), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(G155gat), .ZN(new_n334));
  INV_X1    g133(.A(G162gat), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n334), .A2(new_n335), .A3(KEYINPUT74), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT74), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n337), .B1(G155gat), .B2(G162gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n333), .A2(new_n339), .A3(new_n327), .ZN(new_n340));
  INV_X1    g139(.A(new_n333), .ZN(new_n341));
  XNOR2_X1  g140(.A(G155gat), .B(G162gat), .ZN(new_n342));
  AOI22_X1  g141(.A1(new_n340), .A2(KEYINPUT75), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT3), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT75), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n333), .A2(new_n345), .A3(new_n339), .A4(new_n327), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n343), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(new_n288), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n348), .A2(new_n306), .A3(new_n310), .ZN(new_n349));
  XNOR2_X1  g148(.A(G141gat), .B(G148gat), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n327), .B1(new_n350), .B2(KEYINPUT2), .ZN(new_n351));
  INV_X1    g150(.A(new_n339), .ZN(new_n352));
  OAI21_X1  g151(.A(KEYINPUT75), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n341), .A2(new_n342), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n353), .A2(new_n346), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT29), .B1(new_n309), .B2(new_n303), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n355), .B1(new_n356), .B2(KEYINPUT3), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n349), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(G228gat), .A2(G233gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(G22gat), .ZN(new_n361));
  INV_X1    g160(.A(new_n359), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n349), .A2(new_n362), .A3(new_n357), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n360), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT82), .ZN(new_n365));
  XOR2_X1   g164(.A(KEYINPUT31), .B(G50gat), .Z(new_n366));
  XNOR2_X1  g165(.A(new_n366), .B(KEYINPUT81), .ZN(new_n367));
  XOR2_X1   g166(.A(G78gat), .B(G106gat), .Z(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n363), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n362), .B1(new_n349), .B2(new_n357), .ZN(new_n371));
  OAI21_X1  g170(.A(G22gat), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  AOI22_X1  g171(.A1(new_n365), .A2(new_n369), .B1(new_n372), .B2(new_n364), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT82), .ZN(new_n374));
  AND4_X1   g173(.A1(new_n374), .A2(new_n372), .A3(new_n364), .A4(new_n369), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n355), .A2(KEYINPUT3), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n377), .A2(new_n347), .A3(new_n261), .ZN(new_n378));
  NAND2_X1  g177(.A1(G225gat), .A2(G233gat), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT4), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n380), .B1(new_n355), .B2(new_n261), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n256), .A2(new_n343), .A3(KEYINPUT4), .A4(new_n346), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n378), .A2(new_n379), .A3(new_n381), .A4(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(KEYINPUT76), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n381), .A2(new_n382), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT76), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n385), .A2(new_n386), .A3(new_n379), .A4(new_n378), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n355), .B(new_n256), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT5), .B1(new_n389), .B2(new_n379), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT78), .ZN(new_n393));
  XNOR2_X1  g192(.A(G1gat), .B(G29gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(G57gat), .B(G85gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n396), .B(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n398), .B1(new_n383), .B2(KEYINPUT5), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n392), .A2(new_n393), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n398), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n390), .B1(new_n384), .B2(new_n387), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n383), .A2(KEYINPUT5), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n402), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(KEYINPUT78), .B1(new_n403), .B2(new_n399), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT6), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n401), .A2(new_n405), .A3(new_n406), .A4(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n404), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n392), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n410), .A2(KEYINPUT6), .A3(new_n402), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  AND4_X1   g211(.A1(new_n202), .A2(new_n326), .A3(new_n376), .A4(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n325), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT79), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n411), .B1(new_n408), .B2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n393), .B1(new_n392), .B2(new_n400), .ZN(new_n417));
  NOR3_X1   g216(.A1(new_n403), .A2(KEYINPUT78), .A3(new_n399), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(KEYINPUT6), .B1(new_n410), .B2(new_n402), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT79), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n414), .B1(new_n416), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT80), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT80), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n424), .B(new_n414), .C1(new_n416), .C2(new_n421), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n283), .B1(new_n285), .B2(KEYINPUT70), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT70), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n276), .A2(new_n282), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT87), .ZN(new_n430));
  AND3_X1   g229(.A1(new_n376), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n430), .B1(new_n376), .B2(new_n429), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n423), .A2(new_n425), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n413), .B1(new_n434), .B2(KEYINPUT35), .ZN(new_n435));
  OR2_X1    g234(.A1(new_n287), .A2(KEYINPUT36), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n426), .A2(new_n428), .A3(KEYINPUT36), .ZN(new_n437));
  AND2_X1   g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT86), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n313), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n295), .A2(KEYINPUT86), .A3(new_n312), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n314), .A2(KEYINPUT85), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT85), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n293), .A2(new_n443), .A3(new_n311), .A4(new_n294), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n440), .A2(new_n441), .A3(new_n442), .A4(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT37), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT37), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n313), .A2(new_n447), .A3(new_n314), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT38), .ZN(new_n449));
  AND3_X1   g248(.A1(new_n448), .A2(new_n449), .A3(new_n323), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n446), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(new_n318), .ZN(new_n452));
  INV_X1    g251(.A(new_n317), .ZN(new_n453));
  AND2_X1   g252(.A1(new_n448), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n322), .A2(KEYINPUT37), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n449), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NOR3_X1   g255(.A1(new_n452), .A2(new_n412), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n379), .B1(new_n385), .B2(new_n378), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT39), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n389), .A2(new_n379), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT39), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n460), .B(new_n398), .C1(new_n458), .C2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT83), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT40), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n464), .B1(new_n463), .B2(new_n465), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n325), .B(new_n405), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  OR2_X1    g267(.A1(new_n462), .A2(new_n458), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n469), .A2(KEYINPUT40), .A3(new_n398), .A4(new_n460), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n470), .B(KEYINPUT84), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n376), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n438), .B1(new_n457), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n423), .A2(new_n425), .ZN(new_n474));
  INV_X1    g273(.A(new_n376), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n435), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(G113gat), .B(G141gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n478), .B(G197gat), .ZN(new_n479));
  XOR2_X1   g278(.A(KEYINPUT11), .B(G169gat), .Z(new_n480));
  XNOR2_X1  g279(.A(new_n479), .B(new_n480), .ZN(new_n481));
  XOR2_X1   g280(.A(new_n481), .B(KEYINPUT12), .Z(new_n482));
  XNOR2_X1  g281(.A(G15gat), .B(G22gat), .ZN(new_n483));
  INV_X1    g282(.A(G1gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT16), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n483), .A2(G1gat), .ZN(new_n487));
  OAI21_X1  g286(.A(G8gat), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n483), .A2(new_n485), .ZN(new_n489));
  INV_X1    g288(.A(G8gat), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n489), .B(new_n490), .C1(G1gat), .C2(new_n483), .ZN(new_n491));
  AND2_X1   g290(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g291(.A(G43gat), .B(G50gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT15), .ZN(new_n494));
  OR2_X1    g293(.A1(KEYINPUT88), .A2(G36gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(KEYINPUT88), .A2(G36gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(G29gat), .ZN(new_n498));
  OR3_X1    g297(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n494), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(G43gat), .ZN(new_n503));
  INV_X1    g302(.A(G50gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT15), .ZN(new_n506));
  NAND2_X1  g305(.A1(G43gat), .A2(G50gat), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  AND3_X1   g307(.A1(new_n498), .A2(new_n494), .A3(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT89), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n499), .A2(new_n510), .ZN(new_n511));
  OR4_X1    g310(.A1(new_n510), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(new_n500), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n502), .B1(new_n509), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT90), .B1(new_n492), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n498), .A2(new_n494), .A3(new_n508), .ZN(new_n517));
  INV_X1    g316(.A(new_n500), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n518), .B1(new_n511), .B2(new_n512), .ZN(new_n519));
  AOI22_X1  g318(.A1(new_n497), .A2(G29gat), .B1(new_n499), .B2(new_n500), .ZN(new_n520));
  OAI22_X1  g319(.A1(new_n517), .A2(new_n519), .B1(new_n520), .B2(new_n494), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n488), .A2(new_n491), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT90), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n516), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(G229gat), .A2(G233gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n515), .A2(KEYINPUT17), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT17), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n521), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n527), .A2(new_n492), .A3(new_n529), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n525), .A2(KEYINPUT18), .A3(new_n526), .A4(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n492), .A2(new_n515), .ZN(new_n532));
  AND3_X1   g331(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n523), .B1(new_n521), .B2(new_n522), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  XOR2_X1   g334(.A(new_n526), .B(KEYINPUT13), .Z(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n531), .A2(new_n537), .A3(KEYINPUT91), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n525), .A2(new_n526), .A3(new_n530), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT18), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(KEYINPUT91), .B1(new_n531), .B2(new_n537), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n482), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT92), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI211_X1 g345(.A(KEYINPUT92), .B(new_n482), .C1(new_n542), .C2(new_n543), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n481), .B(KEYINPUT12), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n541), .A2(new_n537), .A3(new_n531), .A4(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  XOR2_X1   g351(.A(G71gat), .B(G78gat), .Z(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(KEYINPUT93), .ZN(new_n554));
  XOR2_X1   g353(.A(G57gat), .B(G64gat), .Z(new_n555));
  INV_X1    g354(.A(KEYINPUT9), .ZN(new_n556));
  INV_X1    g355(.A(G71gat), .ZN(new_n557));
  INV_X1    g356(.A(G78gat), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(G71gat), .B(G78gat), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT93), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n554), .A2(new_n560), .A3(new_n563), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n553), .A2(new_n555), .A3(KEYINPUT93), .A4(new_n559), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n566), .A2(KEYINPUT21), .ZN(new_n567));
  NAND2_X1  g366(.A1(G231gat), .A2(G233gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(G127gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n522), .B1(KEYINPUT21), .B2(new_n566), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(G155gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(G183gat), .B(G211gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  OR2_X1    g376(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n573), .A2(new_n577), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g379(.A1(G85gat), .A2(G92gat), .ZN(new_n581));
  NOR2_X1   g380(.A1(KEYINPUT95), .A2(KEYINPUT7), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(G85gat), .A2(G92gat), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT7), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n584), .B1(new_n585), .B2(KEYINPUT94), .ZN(new_n586));
  AND2_X1   g385(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT94), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n588), .A2(KEYINPUT95), .A3(KEYINPUT7), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n589), .A2(new_n584), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  XOR2_X1   g390(.A(G99gat), .B(G106gat), .Z(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(G99gat), .ZN(new_n594));
  INV_X1    g393(.A(G106gat), .ZN(new_n595));
  OAI21_X1  g394(.A(KEYINPUT8), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n587), .A2(new_n591), .A3(new_n593), .A4(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n583), .A2(new_n586), .A3(new_n596), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n592), .B1(new_n598), .B2(new_n590), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n527), .A2(new_n529), .A3(new_n600), .ZN(new_n601));
  AND2_X1   g400(.A1(G232gat), .A2(G233gat), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(KEYINPUT41), .ZN(new_n603));
  OAI211_X1 g402(.A(new_n601), .B(new_n603), .C1(new_n515), .C2(new_n600), .ZN(new_n604));
  XOR2_X1   g403(.A(G190gat), .B(G218gat), .Z(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n602), .A2(KEYINPUT41), .ZN(new_n607));
  XNOR2_X1  g406(.A(G134gat), .B(G162gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  OR2_X1    g409(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n606), .A2(new_n610), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(G230gat), .A2(G233gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(KEYINPUT97), .B(KEYINPUT10), .ZN(new_n615));
  AND2_X1   g414(.A1(new_n564), .A2(new_n565), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(new_n600), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n566), .A2(new_n597), .A3(new_n599), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n617), .A2(KEYINPUT96), .A3(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT96), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n616), .A2(new_n600), .A3(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n615), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT10), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n618), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n614), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n619), .A2(G230gat), .A3(G233gat), .A4(new_n621), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(G120gat), .B(G148gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(G176gat), .B(G204gat), .ZN(new_n629));
  XOR2_X1   g428(.A(new_n628), .B(new_n629), .Z(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n625), .A2(new_n626), .A3(new_n630), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n580), .A2(new_n613), .A3(new_n635), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n636), .B(KEYINPUT98), .Z(new_n637));
  NOR3_X1   g436(.A1(new_n477), .A2(new_n552), .A3(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n416), .A2(new_n421), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g440(.A1(new_n638), .A2(new_n325), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(KEYINPUT99), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(G8gat), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n643), .A2(KEYINPUT42), .A3(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT42), .ZN(new_n647));
  INV_X1    g446(.A(new_n645), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n647), .B1(new_n642), .B2(new_n648), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n646), .B(new_n649), .C1(new_n490), .C2(new_n643), .ZN(G1325gat));
  INV_X1    g449(.A(G15gat), .ZN(new_n651));
  INV_X1    g450(.A(new_n287), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n638), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n438), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n653), .B1(new_n656), .B2(new_n651), .ZN(G1326gat));
  NAND2_X1  g456(.A1(new_n638), .A2(new_n475), .ZN(new_n658));
  XNOR2_X1  g457(.A(KEYINPUT43), .B(G22gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(G1327gat));
  INV_X1    g459(.A(new_n613), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n661), .B1(new_n435), .B2(new_n476), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NOR3_X1   g462(.A1(new_n552), .A2(new_n580), .A3(new_n634), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n639), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n665), .A2(G29gat), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT100), .B(KEYINPUT45), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT44), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n662), .A2(new_n670), .ZN(new_n671));
  OAI211_X1 g470(.A(KEYINPUT44), .B(new_n661), .C1(new_n435), .C2(new_n476), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g472(.A(new_n664), .B(KEYINPUT101), .Z(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(G29gat), .B1(new_n675), .B2(new_n666), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n669), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT102), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1328gat));
  NOR3_X1   g478(.A1(new_n665), .A2(new_n414), .A3(new_n497), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT46), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n497), .B1(new_n675), .B2(new_n414), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(G1329gat));
  OAI21_X1  g482(.A(new_n503), .B1(new_n665), .B2(new_n287), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n654), .A2(G43gat), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n684), .B1(new_n675), .B2(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g486(.A(G50gat), .B1(new_n675), .B2(new_n376), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n475), .A2(new_n504), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT104), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT103), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n690), .B1(new_n665), .B2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n665), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n693), .A2(KEYINPUT103), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n688), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n695), .B(KEYINPUT48), .Z(G1331gat));
  NAND3_X1  g495(.A1(new_n580), .A2(new_n613), .A3(new_n634), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n477), .A2(new_n551), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(new_n639), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g499(.A(new_n414), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  XOR2_X1   g501(.A(new_n702), .B(KEYINPUT105), .Z(new_n703));
  NOR2_X1   g502(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n703), .B(new_n704), .ZN(G1333gat));
  AOI21_X1  g504(.A(new_n557), .B1(new_n698), .B2(new_n654), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n287), .A2(G71gat), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n706), .B1(new_n698), .B2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g508(.A1(new_n698), .A2(new_n475), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g510(.A1(new_n580), .A2(new_n551), .ZN(new_n712));
  OAI211_X1 g511(.A(new_n661), .B(new_n712), .C1(new_n435), .C2(new_n476), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT51), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n714), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  OR4_X1    g517(.A1(G85gat), .A2(new_n718), .A3(new_n666), .A4(new_n635), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n580), .A2(new_n551), .A3(new_n635), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n671), .A2(new_n672), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(KEYINPUT106), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT106), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n671), .A2(new_n723), .A3(new_n672), .A4(new_n720), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n722), .A2(new_n639), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(G85gat), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n719), .A2(new_n726), .ZN(G1336gat));
  NOR2_X1   g526(.A1(new_n414), .A2(G92gat), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n717), .A2(new_n634), .A3(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT52), .ZN(new_n730));
  OAI21_X1  g529(.A(G92gat), .B1(new_n721), .B2(new_n414), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n729), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT108), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n722), .A2(new_n325), .A3(new_n724), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(G92gat), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n715), .A2(KEYINPUT107), .A3(new_n716), .ZN(new_n736));
  OR2_X1    g535(.A1(new_n716), .A2(KEYINPUT107), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n736), .A2(new_n737), .A3(new_n634), .A4(new_n728), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n733), .B1(new_n739), .B2(KEYINPUT52), .ZN(new_n740));
  AOI211_X1 g539(.A(KEYINPUT108), .B(new_n730), .C1(new_n735), .C2(new_n738), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n732), .B1(new_n740), .B2(new_n741), .ZN(G1337gat));
  AND3_X1   g541(.A1(new_n722), .A2(new_n654), .A3(new_n724), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n652), .A2(new_n594), .A3(new_n634), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT109), .ZN(new_n745));
  OAI22_X1  g544(.A1(new_n743), .A2(new_n594), .B1(new_n718), .B2(new_n745), .ZN(G1338gat));
  AND2_X1   g545(.A1(new_n736), .A2(new_n737), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n376), .A2(G106gat), .A3(new_n635), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n722), .A2(new_n475), .A3(new_n724), .ZN(new_n749));
  AOI22_X1  g548(.A1(new_n747), .A2(new_n748), .B1(new_n749), .B2(G106gat), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT53), .ZN(new_n751));
  INV_X1    g550(.A(new_n721), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n595), .B1(new_n752), .B2(new_n475), .ZN(new_n753));
  INV_X1    g552(.A(new_n748), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n751), .B1(new_n718), .B2(new_n754), .ZN(new_n755));
  OAI22_X1  g554(.A1(new_n750), .A2(new_n751), .B1(new_n753), .B2(new_n755), .ZN(G1339gat));
  OR3_X1    g555(.A1(new_n622), .A2(new_n614), .A3(new_n624), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n757), .A2(KEYINPUT54), .A3(new_n625), .ZN(new_n758));
  XOR2_X1   g557(.A(KEYINPUT110), .B(KEYINPUT54), .Z(new_n759));
  OAI211_X1 g558(.A(new_n614), .B(new_n759), .C1(new_n622), .C2(new_n624), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n760), .A2(new_n631), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n758), .A2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n763), .A2(KEYINPUT55), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT55), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n633), .B1(new_n762), .B2(new_n765), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n525), .A2(new_n530), .ZN(new_n767));
  OAI22_X1  g566(.A1(new_n767), .A2(new_n526), .B1(new_n535), .B2(new_n536), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(new_n481), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n550), .ZN(new_n770));
  NOR4_X1   g569(.A1(new_n764), .A2(new_n766), .A3(new_n613), .A4(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n766), .B1(new_n548), .B2(new_n550), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n772), .B1(KEYINPUT55), .B2(new_n763), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n634), .A2(new_n550), .A3(new_n769), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT111), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n771), .B1(new_n776), .B2(new_n613), .ZN(new_n777));
  OAI22_X1  g576(.A1(new_n777), .A2(new_n580), .B1(new_n551), .B2(new_n636), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n778), .A2(new_n639), .A3(new_n414), .A4(new_n433), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(G113gat), .B1(new_n780), .B2(new_n551), .ZN(new_n781));
  AND3_X1   g580(.A1(new_n778), .A2(KEYINPUT112), .A3(new_n376), .ZN(new_n782));
  AOI21_X1  g581(.A(KEYINPUT112), .B1(new_n778), .B2(new_n376), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n639), .B(new_n326), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(KEYINPUT113), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n551), .A2(G113gat), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n781), .B1(new_n785), .B2(new_n786), .ZN(G1340gat));
  INV_X1    g586(.A(G120gat), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n635), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n785), .A2(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n788), .B1(new_n779), .B2(new_n635), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(KEYINPUT114), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT114), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n790), .A2(new_n794), .A3(new_n791), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n795), .ZN(G1341gat));
  NAND3_X1  g595(.A1(new_n780), .A2(new_n570), .A3(new_n580), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n785), .A2(new_n580), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n797), .B1(new_n798), .B2(new_n570), .ZN(G1342gat));
  NAND2_X1  g598(.A1(new_n785), .A2(new_n661), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(G134gat), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n779), .A2(G134gat), .A3(new_n613), .ZN(new_n802));
  XNOR2_X1  g601(.A(KEYINPUT115), .B(KEYINPUT56), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n801), .A2(new_n804), .ZN(G1343gat));
  NOR3_X1   g604(.A1(new_n654), .A2(new_n666), .A3(new_n325), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT57), .B1(new_n778), .B2(new_n475), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n475), .A2(KEYINPUT57), .ZN(new_n809));
  INV_X1    g608(.A(new_n774), .ZN(new_n810));
  AOI21_X1  g609(.A(KEYINPUT55), .B1(new_n762), .B2(KEYINPUT116), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n811), .B1(KEYINPUT116), .B2(new_n762), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n810), .B1(new_n772), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n661), .B1(new_n813), .B2(KEYINPUT117), .ZN(new_n814));
  INV_X1    g613(.A(new_n766), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n812), .A2(new_n551), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n774), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT117), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n771), .B1(new_n814), .B2(new_n819), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n820), .A2(new_n580), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n636), .A2(new_n551), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n809), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n808), .B1(new_n823), .B2(KEYINPUT118), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT118), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n825), .B(new_n809), .C1(new_n821), .C2(new_n822), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n807), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n827), .A2(G141gat), .A3(new_n551), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n778), .A2(new_n475), .A3(new_n806), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n331), .B1(new_n829), .B2(new_n552), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  XOR2_X1   g630(.A(new_n831), .B(KEYINPUT58), .Z(G1344gat));
  INV_X1    g631(.A(new_n829), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n833), .A2(new_n329), .A3(new_n634), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT59), .ZN(new_n835));
  OR2_X1    g634(.A1(new_n637), .A2(new_n551), .ZN(new_n836));
  INV_X1    g635(.A(new_n580), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n837), .B1(new_n820), .B2(KEYINPUT119), .ZN(new_n838));
  INV_X1    g637(.A(new_n771), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n816), .A2(KEYINPUT117), .A3(new_n774), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n613), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n813), .A2(KEYINPUT117), .ZN(new_n842));
  OAI211_X1 g641(.A(KEYINPUT119), .B(new_n839), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n836), .B1(new_n838), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT57), .B1(new_n845), .B2(new_n475), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n778), .A2(new_n809), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n634), .B(new_n806), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n835), .B1(new_n848), .B2(G148gat), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n835), .A2(G148gat), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n850), .B1(new_n827), .B2(new_n634), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n834), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(KEYINPUT120), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT120), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n854), .B(new_n834), .C1(new_n849), .C2(new_n851), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n853), .A2(new_n855), .ZN(G1345gat));
  AOI21_X1  g655(.A(G155gat), .B1(new_n833), .B2(new_n580), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n580), .A2(G155gat), .ZN(new_n858));
  XOR2_X1   g657(.A(new_n858), .B(KEYINPUT121), .Z(new_n859));
  AOI21_X1  g658(.A(new_n857), .B1(new_n827), .B2(new_n859), .ZN(G1346gat));
  AOI21_X1  g659(.A(G162gat), .B1(new_n833), .B2(new_n661), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n613), .A2(new_n335), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n861), .B1(new_n827), .B2(new_n862), .ZN(G1347gat));
  NAND2_X1  g662(.A1(new_n433), .A2(new_n325), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n778), .A2(new_n666), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT122), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n865), .A2(new_n866), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n864), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(G169gat), .B1(new_n870), .B2(new_n551), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n782), .A2(new_n783), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n639), .A2(new_n414), .A3(new_n287), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n551), .A2(G169gat), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n871), .B1(new_n875), .B2(new_n876), .ZN(G1348gat));
  INV_X1    g676(.A(new_n875), .ZN(new_n878));
  OAI21_X1  g677(.A(G176gat), .B1(new_n878), .B2(new_n635), .ZN(new_n879));
  INV_X1    g678(.A(G176gat), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n870), .A2(new_n880), .A3(new_n634), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n879), .A2(new_n881), .ZN(G1349gat));
  OAI21_X1  g681(.A(new_n205), .B1(new_n878), .B2(new_n837), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n580), .A2(new_n208), .ZN(new_n884));
  AOI21_X1  g683(.A(KEYINPUT123), .B1(new_n870), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n886), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g686(.A1(new_n870), .A2(new_n209), .A3(new_n661), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n888), .B(KEYINPUT124), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n661), .B(new_n873), .C1(new_n782), .C2(new_n783), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(G190gat), .ZN(new_n891));
  OR2_X1    g690(.A1(new_n891), .A2(KEYINPUT125), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(KEYINPUT125), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT61), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n892), .A2(KEYINPUT61), .A3(new_n893), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n889), .A2(new_n896), .A3(new_n897), .ZN(G1351gat));
  NAND2_X1  g697(.A1(new_n868), .A2(new_n869), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n654), .A2(new_n414), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n901), .A2(new_n376), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(G197gat), .B1(new_n903), .B2(new_n551), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n846), .A2(new_n847), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n901), .A2(new_n639), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n551), .A2(G197gat), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n904), .B1(new_n908), .B2(new_n909), .ZN(G1352gat));
  INV_X1    g709(.A(G204gat), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n903), .A2(new_n911), .A3(new_n634), .ZN(new_n912));
  OR2_X1    g711(.A1(new_n912), .A2(KEYINPUT62), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(KEYINPUT62), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n905), .A2(new_n635), .A3(new_n907), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n913), .B(new_n914), .C1(new_n911), .C2(new_n915), .ZN(G1353gat));
  NOR3_X1   g715(.A1(new_n905), .A2(new_n837), .A3(new_n907), .ZN(new_n917));
  OAI21_X1  g716(.A(G211gat), .B1(KEYINPUT126), .B2(KEYINPUT63), .ZN(new_n918));
  AND2_X1   g717(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n919));
  OR3_X1    g718(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n919), .B1(new_n917), .B2(new_n918), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n903), .A2(new_n298), .A3(new_n580), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(G1354gat));
  NOR2_X1   g722(.A1(new_n613), .A2(G218gat), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n903), .A2(new_n924), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n905), .A2(new_n613), .A3(new_n907), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n925), .B1(new_n926), .B2(new_n299), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(KEYINPUT127), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT127), .ZN(new_n929));
  OAI211_X1 g728(.A(new_n925), .B(new_n929), .C1(new_n926), .C2(new_n299), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(G1355gat));
endmodule


