//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 1 0 1 1 1 1 0 1 0 0 0 1 0 0 1 0 0 0 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 1 1 0 0 0 0 1 1 1 0 0 1 0 1 0 1 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:31 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT65), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT65), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(G125), .B(G140), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n193), .B1(new_n187), .B2(new_n192), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT81), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT81), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n193), .B(new_n196), .C1(new_n187), .C2(new_n192), .ZN(new_n197));
  INV_X1    g011(.A(G237), .ZN(new_n198));
  INV_X1    g012(.A(G953), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n198), .A2(new_n199), .A3(G214), .ZN(new_n200));
  INV_X1    g014(.A(G143), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n198), .A2(new_n199), .A3(G143), .A4(G214), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT18), .ZN(new_n205));
  INV_X1    g019(.A(G131), .ZN(new_n206));
  OAI22_X1  g020(.A1(new_n204), .A2(KEYINPUT82), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT82), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n205), .A2(new_n206), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n202), .A2(new_n208), .A3(new_n209), .A4(new_n203), .ZN(new_n210));
  AOI22_X1  g024(.A1(new_n195), .A2(new_n197), .B1(new_n207), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  XNOR2_X1  g026(.A(new_n192), .B(KEYINPUT19), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(new_n191), .ZN(new_n214));
  INV_X1    g028(.A(G140), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G125), .ZN(new_n216));
  OAI21_X1  g030(.A(KEYINPUT71), .B1(new_n216), .B2(KEYINPUT16), .ZN(new_n217));
  INV_X1    g031(.A(G125), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G140), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n216), .A2(new_n219), .A3(KEYINPUT16), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT71), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT16), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n221), .A2(new_n222), .A3(new_n215), .A4(G125), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n217), .A2(new_n220), .A3(G146), .A4(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n206), .B1(new_n202), .B2(new_n203), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n204), .A2(G131), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n214), .B(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n212), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(G113), .B(G122), .ZN(new_n229));
  INV_X1    g043(.A(G104), .ZN(new_n230));
  XNOR2_X1  g044(.A(new_n229), .B(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n228), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n217), .A2(new_n220), .A3(new_n223), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(new_n187), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n235), .A2(KEYINPUT72), .A3(new_n224), .ZN(new_n236));
  AND2_X1   g050(.A1(new_n220), .A2(new_n223), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT72), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n237), .A2(new_n238), .A3(G146), .A4(new_n217), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n236), .A2(new_n239), .ZN(new_n240));
  OR3_X1    g054(.A1(new_n226), .A2(KEYINPUT17), .A3(new_n225), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n225), .A2(KEYINPUT17), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n240), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n243), .A2(new_n212), .A3(new_n231), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT83), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n242), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n247), .B1(new_n236), .B2(new_n239), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n211), .B1(new_n248), .B2(new_n241), .ZN(new_n249));
  AOI21_X1  g063(.A(KEYINPUT83), .B1(new_n249), .B2(new_n231), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n233), .B1(new_n246), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G475), .ZN(new_n252));
  INV_X1    g066(.A(G902), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT20), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT20), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n251), .A2(new_n256), .A3(new_n252), .A4(new_n253), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  OAI22_X1  g072(.A1(new_n246), .A2(new_n250), .B1(new_n231), .B2(new_n249), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n259), .A2(KEYINPUT84), .A3(new_n253), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT84), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n249), .A2(new_n231), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n244), .A2(new_n245), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n249), .A2(KEYINPUT83), .A3(new_n231), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n262), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n261), .B1(new_n265), .B2(G902), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n260), .A2(new_n266), .A3(G475), .ZN(new_n267));
  INV_X1    g081(.A(G116), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n268), .A2(KEYINPUT14), .A3(G122), .ZN(new_n269));
  XNOR2_X1  g083(.A(G116), .B(G122), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  OAI211_X1 g085(.A(G107), .B(new_n269), .C1(new_n271), .C2(KEYINPUT14), .ZN(new_n272));
  INV_X1    g086(.A(G107), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(G128), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G143), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT85), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n276), .B(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G134), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n201), .A2(G128), .ZN(new_n280));
  AND3_X1   g094(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n279), .B1(new_n278), .B2(new_n280), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n272), .B(new_n274), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n278), .A2(new_n280), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT13), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n276), .A2(new_n277), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT85), .B1(new_n275), .B2(G143), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n284), .A2(G134), .A3(new_n288), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n270), .B(new_n273), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n278), .B(new_n280), .C1(new_n285), .C2(new_n279), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n283), .A2(new_n292), .ZN(new_n293));
  XOR2_X1   g107(.A(KEYINPUT9), .B(G234), .Z(new_n294));
  NAND3_X1  g108(.A1(new_n294), .A2(G217), .A3(new_n199), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT86), .ZN(new_n297));
  INV_X1    g111(.A(new_n295), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n283), .A2(new_n292), .A3(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n296), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n283), .A2(new_n292), .A3(KEYINPUT86), .A4(new_n298), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n300), .A2(new_n253), .A3(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G478), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n303), .A2(KEYINPUT15), .ZN(new_n304));
  OR2_X1    g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n302), .A2(new_n304), .ZN(new_n306));
  XNOR2_X1  g120(.A(KEYINPUT87), .B(G952), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n307), .A2(G953), .ZN(new_n308));
  NAND2_X1  g122(.A1(G234), .A2(G237), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n309), .A2(G902), .A3(G953), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n312), .B(KEYINPUT88), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  XOR2_X1   g128(.A(KEYINPUT21), .B(G898), .Z(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n311), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n305), .A2(new_n306), .A3(new_n318), .ZN(new_n319));
  AND3_X1   g133(.A1(new_n258), .A2(new_n267), .A3(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(G214), .B1(G237), .B2(G902), .ZN(new_n321));
  OAI21_X1  g135(.A(G210), .B1(G237), .B2(G902), .ZN(new_n322));
  OAI21_X1  g136(.A(KEYINPUT3), .B1(new_n230), .B2(G107), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT3), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n324), .A2(new_n273), .A3(G104), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n230), .A2(G107), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n323), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT75), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n323), .A2(new_n325), .A3(KEYINPUT75), .A4(new_n326), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(G101), .A3(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(G101), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n323), .A2(new_n325), .A3(new_n332), .A4(new_n326), .ZN(new_n333));
  AND2_X1   g147(.A1(new_n333), .A2(KEYINPUT4), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT76), .ZN(new_n336));
  OR2_X1    g150(.A1(new_n331), .A2(KEYINPUT4), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT76), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n331), .A2(new_n338), .A3(new_n334), .ZN(new_n339));
  XNOR2_X1  g153(.A(G116), .B(G119), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT68), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  XOR2_X1   g156(.A(KEYINPUT2), .B(G113), .Z(new_n343));
  XNOR2_X1  g157(.A(new_n342), .B(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n336), .A2(new_n337), .A3(new_n339), .A4(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n326), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n230), .A2(G107), .ZN(new_n348));
  OAI21_X1  g162(.A(G101), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n333), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n343), .A2(new_n340), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n340), .A2(KEYINPUT5), .ZN(new_n353));
  INV_X1    g167(.A(G119), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(G116), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n353), .B(G113), .C1(KEYINPUT5), .C2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n351), .A2(new_n352), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n346), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(G110), .B(G122), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n346), .A2(new_n357), .A3(new_n359), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(KEYINPUT6), .A3(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT6), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n358), .A2(new_n364), .A3(new_n360), .ZN(new_n365));
  XNOR2_X1  g179(.A(KEYINPUT65), .B(G146), .ZN(new_n366));
  OAI21_X1  g180(.A(KEYINPUT1), .B1(new_n366), .B2(new_n201), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n201), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n187), .A2(G143), .ZN(new_n369));
  AOI22_X1  g183(.A1(new_n367), .A2(G128), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n201), .B1(new_n188), .B2(new_n190), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n187), .A2(G143), .ZN(new_n372));
  NOR4_X1   g186(.A1(new_n371), .A2(KEYINPUT1), .A3(new_n275), .A4(new_n372), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n218), .ZN(new_n375));
  XNOR2_X1  g189(.A(KEYINPUT0), .B(G128), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n376), .B1(new_n368), .B2(new_n369), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n372), .B1(new_n191), .B2(G143), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n379), .A2(KEYINPUT0), .A3(G128), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G125), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n375), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G224), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n384), .A2(G953), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n383), .B(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n363), .A2(new_n365), .A3(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT79), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n363), .A2(KEYINPUT79), .A3(new_n365), .A4(new_n386), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  XOR2_X1   g205(.A(new_n359), .B(KEYINPUT8), .Z(new_n392));
  NAND2_X1  g206(.A1(new_n356), .A2(new_n352), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n350), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n392), .B1(new_n394), .B2(new_n357), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n395), .B(KEYINPUT80), .ZN(new_n396));
  OAI21_X1  g210(.A(KEYINPUT7), .B1(new_n384), .B2(G953), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n383), .A2(new_n397), .ZN(new_n398));
  OR2_X1    g212(.A1(new_n383), .A2(new_n397), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n396), .A2(new_n362), .A3(new_n398), .A4(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n253), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n322), .B1(new_n391), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n322), .ZN(new_n404));
  AOI211_X1 g218(.A(new_n404), .B(new_n401), .C1(new_n389), .C2(new_n390), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n320), .B(new_n321), .C1(new_n403), .C2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(G469), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n189), .A2(G146), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n187), .A2(KEYINPUT65), .ZN(new_n409));
  OAI21_X1  g223(.A(G143), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT1), .ZN(new_n411));
  INV_X1    g225(.A(new_n372), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n410), .A2(new_n411), .A3(G128), .A4(new_n412), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n201), .A2(G146), .ZN(new_n414));
  OAI21_X1  g228(.A(G128), .B1(new_n414), .B2(new_n411), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n415), .B(KEYINPUT77), .C1(new_n371), .C2(new_n372), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n412), .B1(new_n366), .B2(new_n201), .ZN(new_n418));
  AOI21_X1  g232(.A(KEYINPUT77), .B1(new_n418), .B2(new_n415), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n351), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT78), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  OAI211_X1 g236(.A(KEYINPUT78), .B(new_n351), .C1(new_n417), .C2(new_n419), .ZN(new_n423));
  AOI22_X1  g237(.A1(new_n422), .A2(new_n423), .B1(new_n350), .B2(new_n374), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT12), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT11), .ZN(new_n426));
  AOI22_X1  g240(.A1(KEYINPUT66), .A2(new_n426), .B1(new_n279), .B2(G137), .ZN(new_n427));
  OAI22_X1  g241(.A1(KEYINPUT66), .A2(new_n426), .B1(new_n279), .B2(G137), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT66), .ZN(new_n429));
  INV_X1    g243(.A(G137), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n429), .A2(new_n430), .A3(KEYINPUT11), .A4(G134), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n427), .A2(new_n428), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(G131), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n427), .A2(new_n428), .A3(new_n206), .A4(new_n431), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  NOR3_X1   g250(.A1(new_n424), .A2(new_n425), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n374), .A2(new_n350), .ZN(new_n438));
  INV_X1    g252(.A(new_n423), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT77), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n275), .B1(new_n369), .B2(KEYINPUT1), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n440), .B1(new_n379), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n442), .A2(new_n416), .A3(new_n413), .ZN(new_n443));
  AOI21_X1  g257(.A(KEYINPUT78), .B1(new_n443), .B2(new_n351), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n438), .B1(new_n439), .B2(new_n444), .ZN(new_n445));
  AND3_X1   g259(.A1(new_n433), .A2(KEYINPUT69), .A3(new_n434), .ZN(new_n446));
  AOI21_X1  g260(.A(KEYINPUT69), .B1(new_n433), .B2(new_n434), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(KEYINPUT12), .B1(new_n445), .B2(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n437), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT10), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n452), .B1(new_n439), .B2(new_n444), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n418), .A2(new_n275), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n377), .B1(new_n454), .B2(KEYINPUT0), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n336), .A2(new_n337), .A3(new_n339), .A4(new_n455), .ZN(new_n456));
  OAI211_X1 g270(.A(KEYINPUT10), .B(new_n351), .C1(new_n370), .C2(new_n373), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n453), .A2(new_n456), .A3(new_n457), .A4(new_n448), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n199), .A2(G227), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n459), .B(KEYINPUT74), .ZN(new_n460));
  XNOR2_X1  g274(.A(G110), .B(G140), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n460), .B(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n458), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n451), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n456), .A2(new_n457), .ZN(new_n465));
  AOI21_X1  g279(.A(KEYINPUT10), .B1(new_n422), .B2(new_n423), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n449), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n462), .B1(new_n467), .B2(new_n458), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n407), .B(new_n253), .C1(new_n464), .C2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n467), .A2(new_n458), .A3(new_n462), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n425), .B1(new_n424), .B2(new_n448), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n445), .A2(KEYINPUT12), .A3(new_n435), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n465), .A2(new_n466), .ZN(new_n473));
  AOI22_X1  g287(.A1(new_n471), .A2(new_n472), .B1(new_n473), .B2(new_n448), .ZN(new_n474));
  OAI211_X1 g288(.A(G469), .B(new_n470), .C1(new_n474), .C2(new_n462), .ZN(new_n475));
  NAND2_X1  g289(.A1(G469), .A2(G902), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n469), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(G221), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n478), .B1(new_n294), .B2(new_n253), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(KEYINPUT89), .B1(new_n406), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n321), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n391), .A2(new_n402), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n404), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n391), .A2(new_n322), .A3(new_n402), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n483), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n481), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT89), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n487), .A2(new_n488), .A3(new_n489), .A4(new_n320), .ZN(new_n490));
  XNOR2_X1  g304(.A(G134), .B(G137), .ZN(new_n491));
  OR3_X1    g305(.A1(new_n491), .A2(KEYINPUT67), .A3(new_n206), .ZN(new_n492));
  OAI21_X1  g306(.A(KEYINPUT67), .B1(new_n491), .B2(new_n206), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n434), .A2(new_n493), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n492), .B(new_n494), .C1(new_n370), .C2(new_n373), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n435), .A2(new_n378), .A3(new_n380), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  XNOR2_X1  g311(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n455), .B1(new_n446), .B2(new_n447), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n500), .A2(KEYINPUT30), .A3(new_n495), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n499), .A2(new_n501), .A3(new_n345), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n500), .A2(new_n344), .A3(new_n495), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n198), .A2(new_n199), .A3(G210), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n504), .B(new_n332), .ZN(new_n505));
  XNOR2_X1  g319(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n506));
  XOR2_X1   g320(.A(new_n505), .B(new_n506), .Z(new_n507));
  NAND3_X1  g321(.A1(new_n502), .A2(new_n503), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT31), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n503), .A2(KEYINPUT28), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT28), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n500), .A2(new_n511), .A3(new_n344), .A4(new_n495), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n497), .A2(new_n345), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n507), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT31), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n502), .A2(new_n518), .A3(new_n503), .A4(new_n507), .ZN(new_n519));
  AND2_X1   g333(.A1(new_n519), .A2(KEYINPUT70), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n519), .A2(KEYINPUT70), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n509), .B(new_n517), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(G472), .A2(G902), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT32), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n522), .A2(KEYINPUT32), .A3(new_n523), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n515), .A2(new_n516), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n507), .B1(new_n502), .B2(new_n503), .ZN(new_n529));
  NOR3_X1   g343(.A1(new_n528), .A2(new_n529), .A3(KEYINPUT29), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n500), .A2(new_n495), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n345), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n533), .B1(new_n510), .B2(new_n512), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n534), .A2(KEYINPUT29), .A3(new_n507), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n253), .ZN(new_n536));
  OAI21_X1  g350(.A(G472), .B1(new_n530), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n526), .A2(new_n527), .A3(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT23), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n539), .B1(new_n354), .B2(G128), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n354), .A2(G128), .ZN(new_n541));
  MUX2_X1   g355(.A(new_n540), .B(new_n539), .S(new_n541), .Z(new_n542));
  INV_X1    g356(.A(G110), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  XOR2_X1   g358(.A(new_n544), .B(KEYINPUT73), .Z(new_n545));
  XOR2_X1   g359(.A(G119), .B(G128), .Z(new_n546));
  XNOR2_X1  g360(.A(KEYINPUT24), .B(G110), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n193), .B(new_n224), .C1(new_n545), .C2(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n542), .A2(new_n543), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n240), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n551), .B1(new_n546), .B2(new_n547), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g367(.A(KEYINPUT22), .B(G137), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n199), .A2(G221), .A3(G234), .ZN(new_n555));
  XOR2_X1   g369(.A(new_n554), .B(new_n555), .Z(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n549), .A2(new_n552), .A3(new_n556), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(G217), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n561), .B1(G234), .B2(new_n253), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n562), .A2(G902), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n558), .A2(new_n253), .A3(new_n559), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT25), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n566), .B(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n565), .B1(new_n568), .B2(new_n562), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n538), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n482), .A2(new_n490), .A3(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n572), .B(G101), .ZN(G3));
  NAND2_X1  g387(.A1(new_n487), .A2(new_n318), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n522), .A2(new_n253), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(G472), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n524), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n566), .A2(new_n567), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n566), .A2(new_n567), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n562), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n581), .B1(new_n560), .B2(new_n564), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n578), .A2(new_n582), .A3(new_n481), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n575), .A2(new_n583), .ZN(new_n584));
  AOI22_X1  g398(.A1(new_n263), .A2(new_n264), .B1(new_n232), .B2(new_n228), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n585), .A2(G475), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n256), .B1(new_n586), .B2(new_n253), .ZN(new_n587));
  INV_X1    g401(.A(new_n257), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n267), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT33), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n300), .A2(new_n590), .A3(new_n301), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n296), .A2(KEYINPUT33), .A3(new_n299), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n591), .A2(G478), .A3(new_n253), .A4(new_n592), .ZN(new_n593));
  OR2_X1    g407(.A1(new_n593), .A2(KEYINPUT90), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n302), .A2(new_n303), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n593), .A2(KEYINPUT90), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n589), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n584), .A2(new_n598), .ZN(new_n599));
  XOR2_X1   g413(.A(KEYINPUT34), .B(G104), .Z(new_n600));
  XNOR2_X1  g414(.A(new_n599), .B(new_n600), .ZN(G6));
  NAND2_X1  g415(.A1(new_n588), .A2(KEYINPUT91), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT91), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n257), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n602), .A2(new_n255), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n305), .A2(new_n306), .ZN(new_n606));
  AND3_X1   g420(.A1(new_n605), .A2(new_n267), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n584), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(G107), .ZN(new_n609));
  XNOR2_X1  g423(.A(KEYINPUT92), .B(KEYINPUT35), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(G9));
  INV_X1    g425(.A(new_n578), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n557), .A2(KEYINPUT36), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n553), .B(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n563), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n581), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n482), .A2(new_n490), .A3(new_n612), .A4(new_n616), .ZN(new_n617));
  XOR2_X1   g431(.A(KEYINPUT37), .B(G110), .Z(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(KEYINPUT93), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n617), .B(new_n619), .ZN(G12));
  AND3_X1   g434(.A1(new_n522), .A2(KEYINPUT32), .A3(new_n523), .ZN(new_n621));
  AOI21_X1  g435(.A(KEYINPUT32), .B1(new_n522), .B2(new_n523), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n481), .B1(new_n623), .B2(new_n537), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n310), .B(KEYINPUT94), .ZN(new_n625));
  INV_X1    g439(.A(G900), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n625), .B1(new_n626), .B2(new_n314), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  AND4_X1   g442(.A1(new_n267), .A2(new_n605), .A3(new_n606), .A4(new_n628), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n624), .A2(new_n487), .A3(new_n616), .A4(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(G128), .ZN(G30));
  XNOR2_X1  g445(.A(KEYINPUT97), .B(KEYINPUT39), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n627), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n488), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(KEYINPUT40), .ZN(new_n635));
  AOI22_X1  g449(.A1(new_n568), .A2(new_n562), .B1(new_n563), .B2(new_n614), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT40), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n488), .A2(new_n637), .A3(new_n633), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n635), .A2(new_n321), .A3(new_n636), .A4(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n503), .A2(new_n516), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n253), .B1(new_n533), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n516), .B1(new_n502), .B2(new_n503), .ZN(new_n642));
  OAI21_X1  g456(.A(G472), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n623), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT96), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n485), .A2(new_n486), .A3(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n647), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n649), .B1(new_n403), .B2(new_n405), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n589), .A2(new_n606), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n639), .A2(new_n646), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(new_n201), .ZN(G45));
  NAND3_X1  g470(.A1(new_n589), .A2(new_n597), .A3(new_n628), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n624), .A2(new_n487), .A3(new_n616), .A4(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G146), .ZN(G48));
  INV_X1    g474(.A(new_n468), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n661), .B1(new_n451), .B2(new_n463), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n253), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(G469), .ZN(new_n664));
  AND3_X1   g478(.A1(new_n664), .A2(new_n480), .A3(new_n469), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n575), .A2(new_n571), .A3(new_n598), .A4(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT41), .B(G113), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G15));
  NAND4_X1  g482(.A1(new_n487), .A2(new_n607), .A3(new_n665), .A4(new_n538), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n569), .A2(new_n318), .ZN(new_n670));
  OR2_X1    g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G116), .ZN(G18));
  NAND4_X1  g486(.A1(new_n665), .A2(new_n487), .A3(new_n538), .A4(new_n616), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT98), .ZN(new_n674));
  INV_X1    g488(.A(new_n320), .ZN(new_n675));
  OR3_X1    g489(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n674), .B1(new_n673), .B2(new_n675), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G119), .ZN(G21));
  OAI221_X1 g493(.A(new_n509), .B1(new_n507), .B2(new_n534), .C1(new_n520), .C2(new_n521), .ZN(new_n680));
  XOR2_X1   g494(.A(new_n523), .B(KEYINPUT99), .Z(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n577), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n683), .A2(new_n582), .ZN(new_n684));
  AND2_X1   g498(.A1(new_n684), .A2(new_n665), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n652), .A2(KEYINPUT100), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT100), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n589), .A2(new_n687), .A3(new_n606), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n685), .A2(new_n575), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G122), .ZN(G24));
  NOR2_X1   g505(.A1(new_n683), .A2(new_n636), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n692), .A2(new_n487), .A3(new_n658), .A4(new_n665), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G125), .ZN(G27));
  INV_X1    g508(.A(KEYINPUT106), .ZN(new_n695));
  AND3_X1   g509(.A1(new_n538), .A2(KEYINPUT105), .A3(new_n569), .ZN(new_n696));
  AOI21_X1  g510(.A(KEYINPUT105), .B1(new_n538), .B2(new_n569), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n485), .A2(new_n321), .A3(new_n486), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n699), .A2(new_n657), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT101), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n475), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n458), .B1(new_n437), .B2(new_n450), .ZN(new_n703));
  INV_X1    g517(.A(new_n462), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n705), .A2(KEYINPUT101), .A3(G469), .A4(new_n470), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n702), .A2(new_n469), .A3(new_n476), .A4(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT102), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n707), .A2(new_n708), .A3(new_n480), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n708), .B1(new_n707), .B2(new_n480), .ZN(new_n711));
  OAI211_X1 g525(.A(new_n700), .B(KEYINPUT42), .C1(new_n710), .C2(new_n711), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n695), .B1(new_n698), .B2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT105), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n570), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n538), .A2(KEYINPUT105), .A3(new_n569), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT42), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n707), .A2(new_n480), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(KEYINPUT102), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n718), .B1(new_n720), .B2(new_n709), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n717), .A2(KEYINPUT106), .A3(new_n721), .A4(new_n700), .ZN(new_n722));
  AND2_X1   g536(.A1(new_n713), .A2(new_n722), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n403), .A2(new_n405), .A3(new_n483), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n724), .A2(new_n538), .A3(new_n569), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n720), .A2(new_n709), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n725), .A2(new_n726), .A3(new_n658), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT103), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n725), .A2(new_n726), .A3(KEYINPUT103), .A4(new_n658), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n729), .A2(new_n718), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(KEYINPUT104), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT104), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n729), .A2(new_n733), .A3(new_n718), .A4(new_n730), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n723), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(new_n206), .ZN(G33));
  NAND3_X1  g550(.A1(new_n725), .A2(new_n726), .A3(new_n629), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT107), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n737), .B(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G134), .ZN(G36));
  NAND2_X1  g554(.A1(new_n705), .A2(new_n470), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT45), .ZN(new_n742));
  OAI21_X1  g556(.A(KEYINPUT108), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n407), .B1(new_n741), .B2(new_n742), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT108), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n705), .A2(new_n745), .A3(KEYINPUT45), .A4(new_n470), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n743), .A2(new_n744), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n476), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT46), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n747), .A2(KEYINPUT46), .A3(new_n476), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n750), .A2(new_n469), .A3(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(new_n480), .A3(new_n633), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n597), .A2(new_n258), .A3(new_n267), .ZN(new_n755));
  NOR2_X1   g569(.A1(KEYINPUT109), .A2(KEYINPUT43), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(KEYINPUT109), .A2(KEYINPUT43), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n756), .B1(new_n755), .B2(new_n758), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n578), .B(new_n616), .C1(new_n757), .C2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT44), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n699), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n754), .B(new_n762), .C1(new_n761), .C2(new_n760), .ZN(new_n763));
  XNOR2_X1  g577(.A(KEYINPUT110), .B(G137), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n763), .B(new_n764), .ZN(G39));
  NOR2_X1   g579(.A1(new_n538), .A2(new_n569), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n752), .A2(KEYINPUT47), .A3(new_n480), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(KEYINPUT47), .B1(new_n752), .B2(new_n480), .ZN(new_n769));
  OAI211_X1 g583(.A(new_n700), .B(new_n766), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(KEYINPUT111), .ZN(new_n771));
  INV_X1    g585(.A(new_n769), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n767), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT111), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n773), .A2(new_n774), .A3(new_n700), .A4(new_n766), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n771), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G140), .ZN(G42));
  OR2_X1    g591(.A1(new_n757), .A2(new_n759), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n778), .A2(new_n625), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n724), .ZN(new_n780));
  INV_X1    g594(.A(new_n665), .ZN(new_n781));
  OR3_X1    g595(.A1(new_n780), .A2(KEYINPUT116), .A3(new_n781), .ZN(new_n782));
  OAI21_X1  g596(.A(KEYINPUT116), .B1(new_n780), .B2(new_n781), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n692), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n779), .A2(new_n685), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n321), .B1(new_n648), .B2(new_n650), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT50), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n786), .A2(KEYINPUT50), .A3(new_n787), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g606(.A1(KEYINPUT117), .A2(KEYINPUT51), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n785), .A2(new_n792), .A3(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT117), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT51), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n781), .A2(new_n582), .A3(new_n699), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n646), .A2(new_n311), .A3(new_n799), .ZN(new_n800));
  OR3_X1    g614(.A1(new_n800), .A2(new_n589), .A3(new_n597), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n664), .A2(new_n469), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n772), .B(new_n767), .C1(new_n480), .C2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(new_n780), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n803), .A2(new_n684), .A3(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n795), .A2(new_n798), .A3(new_n801), .A4(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n785), .A2(new_n801), .A3(new_n792), .A4(new_n794), .ZN(new_n807));
  INV_X1    g621(.A(new_n805), .ZN(new_n808));
  OAI22_X1  g622(.A1(new_n807), .A2(new_n808), .B1(new_n796), .B2(new_n797), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n806), .A2(new_n809), .A3(new_n308), .ZN(new_n810));
  XNOR2_X1  g624(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n732), .A2(new_n734), .ZN(new_n812));
  INV_X1    g626(.A(new_n723), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n321), .B1(new_n403), .B2(new_n405), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n815), .B1(new_n686), .B2(new_n688), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n616), .B1(new_n623), .B2(new_n643), .ZN(new_n817));
  INV_X1    g631(.A(new_n719), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n816), .A2(new_n817), .A3(new_n628), .A4(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n819), .A2(new_n630), .A3(new_n659), .A4(new_n693), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT52), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n487), .A2(new_n488), .A3(new_n538), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n823), .B(new_n616), .C1(new_n629), .C2(new_n658), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n824), .A2(KEYINPUT52), .A3(new_n693), .A4(new_n819), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT113), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n598), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n589), .A2(new_n597), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(KEYINPUT113), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n258), .A2(new_n267), .A3(new_n606), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n828), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n575), .A2(new_n832), .A3(new_n583), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n617), .A2(new_n572), .A3(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n683), .A2(new_n657), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n835), .B1(new_n710), .B2(new_n711), .ZN(new_n836));
  INV_X1    g650(.A(new_n606), .ZN(new_n837));
  AND4_X1   g651(.A1(new_n267), .A2(new_n605), .A3(new_n837), .A4(new_n628), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n838), .A2(new_n488), .A3(new_n538), .ZN(new_n839));
  AOI211_X1 g653(.A(new_n636), .B(new_n699), .C1(new_n836), .C2(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n834), .A2(new_n840), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n826), .A2(new_n739), .A3(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n678), .A2(new_n671), .A3(new_n666), .A4(new_n690), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n814), .A2(new_n842), .A3(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n826), .A2(KEYINPUT114), .A3(new_n739), .A4(new_n841), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n846), .A2(KEYINPUT53), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n826), .A2(new_n739), .A3(new_n841), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n735), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n846), .A2(KEYINPUT53), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n850), .A2(new_n851), .A3(new_n844), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n811), .B1(new_n848), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n845), .A2(KEYINPUT53), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT53), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n850), .A2(new_n855), .A3(new_n844), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n853), .B1(KEYINPUT54), .B2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n800), .ZN(new_n859));
  AOI22_X1  g673(.A1(new_n786), .A2(new_n487), .B1(new_n859), .B2(new_n598), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n784), .A2(new_n717), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n861), .B(KEYINPUT48), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n810), .A2(new_n858), .A3(new_n860), .A4(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n863), .B1(G952), .B2(G953), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n569), .A2(new_n480), .A3(new_n321), .ZN(new_n865));
  XOR2_X1   g679(.A(new_n865), .B(KEYINPUT112), .Z(new_n866));
  INV_X1    g680(.A(new_n755), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n867), .B1(KEYINPUT49), .B2(new_n802), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n868), .B1(KEYINPUT49), .B2(new_n802), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n866), .A2(new_n646), .A3(new_n651), .A4(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n864), .A2(new_n870), .ZN(G75));
  NOR2_X1   g685(.A1(new_n845), .A2(new_n847), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n851), .B1(new_n850), .B2(new_n844), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n872), .A2(new_n873), .A3(new_n253), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(G210), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT56), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n363), .A2(new_n365), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n877), .B(new_n386), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(KEYINPUT55), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n875), .A2(new_n876), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n879), .B1(new_n875), .B2(new_n876), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n199), .A2(G952), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(G51));
  XOR2_X1   g697(.A(new_n476), .B(KEYINPUT57), .Z(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(new_n811), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n886), .B1(new_n872), .B2(new_n873), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n848), .A2(new_n852), .A3(new_n811), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n885), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(new_n662), .ZN(new_n890));
  OAI21_X1  g704(.A(KEYINPUT118), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n848), .A2(new_n852), .A3(new_n811), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n884), .B1(new_n892), .B2(new_n853), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT118), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n893), .A2(new_n894), .A3(new_n662), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n747), .B(KEYINPUT119), .Z(new_n896));
  NAND2_X1  g710(.A1(new_n874), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n891), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(new_n882), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n898), .A2(new_n899), .ZN(G54));
  NAND3_X1  g714(.A1(new_n874), .A2(KEYINPUT58), .A3(G475), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT120), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n901), .A2(new_n902), .A3(new_n585), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n899), .B1(new_n901), .B2(new_n585), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n902), .B1(new_n901), .B2(new_n585), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(G60));
  AND2_X1   g721(.A1(new_n591), .A2(new_n592), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(G478), .A2(G902), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n910), .B(KEYINPUT59), .Z(new_n911));
  AOI211_X1 g725(.A(new_n909), .B(new_n911), .C1(new_n887), .C2(new_n888), .ZN(new_n912));
  OAI211_X1 g726(.A(KEYINPUT121), .B(new_n909), .C1(new_n858), .C2(new_n911), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT121), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n854), .A2(KEYINPUT54), .A3(new_n856), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n911), .B1(new_n887), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n914), .B1(new_n916), .B2(new_n908), .ZN(new_n917));
  AOI211_X1 g731(.A(new_n882), .B(new_n912), .C1(new_n913), .C2(new_n917), .ZN(G63));
  NOR2_X1   g732(.A1(new_n872), .A2(new_n873), .ZN(new_n919));
  NAND2_X1  g733(.A1(G217), .A2(G902), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT60), .Z(new_n921));
  NAND2_X1  g735(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(new_n560), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n919), .A2(new_n614), .A3(new_n921), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n923), .A2(new_n899), .A3(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT61), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n925), .B(new_n926), .ZN(G66));
  OAI21_X1  g741(.A(G953), .B1(new_n316), .B2(new_n384), .ZN(new_n928));
  OAI21_X1  g742(.A(KEYINPUT122), .B1(new_n843), .B2(new_n834), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n671), .A2(new_n666), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n930), .B1(new_n677), .B2(new_n676), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT122), .ZN(new_n932));
  INV_X1    g746(.A(new_n834), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n931), .A2(new_n932), .A3(new_n933), .A4(new_n690), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n929), .A2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n928), .B1(new_n936), .B2(G953), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n877), .B1(G898), .B2(new_n199), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n937), .B(new_n938), .ZN(G69));
  NAND2_X1  g753(.A1(new_n499), .A2(new_n501), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(new_n213), .ZN(new_n941));
  OR3_X1    g755(.A1(new_n639), .A2(new_n646), .A3(new_n654), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n824), .A2(new_n693), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n942), .A2(new_n944), .A3(KEYINPUT62), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT62), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n946), .B1(new_n655), .B2(new_n943), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n725), .A2(new_n832), .A3(new_n488), .A4(new_n633), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n776), .A2(new_n763), .A3(new_n948), .A4(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n941), .B1(new_n951), .B2(G953), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n626), .A2(new_n199), .ZN(new_n953));
  INV_X1    g767(.A(new_n941), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n763), .A2(new_n739), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n955), .B1(new_n771), .B2(new_n775), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n753), .A2(new_n698), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n943), .B1(new_n957), .B2(new_n816), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n956), .A2(new_n814), .A3(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n954), .B1(new_n959), .B2(G953), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n952), .B1(new_n953), .B2(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n199), .B1(G227), .B2(G900), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n961), .B(new_n962), .ZN(G72));
  NAND2_X1  g777(.A1(G472), .A2(G902), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT63), .Z(new_n965));
  OAI21_X1  g779(.A(new_n965), .B1(new_n950), .B2(new_n935), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n642), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(KEYINPUT123), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT123), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n966), .A2(new_n969), .A3(new_n642), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n508), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n529), .B(KEYINPUT126), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n857), .B(new_n965), .C1(new_n972), .C2(new_n973), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n502), .A2(new_n503), .A3(new_n516), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT124), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n936), .A2(new_n814), .A3(new_n958), .A4(new_n956), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n977), .B1(new_n978), .B2(new_n965), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT125), .ZN(new_n980));
  NOR3_X1   g794(.A1(new_n979), .A2(new_n980), .A3(new_n882), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n965), .B1(new_n959), .B2(new_n935), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n976), .ZN(new_n983));
  AOI21_X1  g797(.A(KEYINPUT125), .B1(new_n983), .B2(new_n899), .ZN(new_n984));
  OAI211_X1 g798(.A(new_n971), .B(new_n974), .C1(new_n981), .C2(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(KEYINPUT127), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n980), .B1(new_n979), .B2(new_n882), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n983), .A2(KEYINPUT125), .A3(new_n899), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT127), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n989), .A2(new_n990), .A3(new_n971), .A4(new_n974), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n986), .A2(new_n991), .ZN(G57));
endmodule


