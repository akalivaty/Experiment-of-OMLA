//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 0 1 0 0 1 0 1 1 0 1 1 0 0 0 0 0 0 1 1 1 1 1 0 0 0 0 0 1 0 1 1 0 1 0 0 1 1 1 0 1 0 1 1 1 0 0 0 1 0 1 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:28 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1283, new_n1284, new_n1285,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n221));
  INV_X1    g0021(.A(G77), .ZN(new_n222));
  INV_X1    g0022(.A(G244), .ZN(new_n223));
  INV_X1    g0023(.A(G107), .ZN(new_n224));
  INV_X1    g0024(.A(G264), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n211), .B1(new_n220), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n228), .A2(new_n209), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT64), .ZN(new_n230));
  INV_X1    g0030(.A(new_n201), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(G50), .ZN(new_n232));
  OAI221_X1 g0032(.A(new_n214), .B1(KEYINPUT1), .B2(new_n227), .C1(new_n230), .C2(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n202), .A2(G68), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n216), .A2(G50), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n245), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(G13), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(G1), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G20), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n254), .A2(G116), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n228), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  OAI211_X1 g0059(.A(new_n258), .B(new_n254), .C1(G1), .C2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n255), .B1(new_n261), .B2(G116), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G33), .A2(G283), .ZN(new_n263));
  INV_X1    g0063(.A(G97), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n263), .B(new_n209), .C1(G33), .C2(new_n264), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n265), .B(new_n257), .C1(new_n209), .C2(G116), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT20), .ZN(new_n267));
  XNOR2_X1  g0067(.A(new_n266), .B(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n262), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G169), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT21), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AND2_X1   g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  NOR2_X1   g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G264), .A2(G1698), .ZN(new_n276));
  OAI21_X1  g0076(.A(KEYINPUT81), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT3), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n259), .ZN(new_n279));
  NAND2_X1  g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G1698), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n281), .A2(G257), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n275), .A2(G303), .ZN(new_n284));
  INV_X1    g0084(.A(new_n276), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT81), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n285), .B(new_n286), .C1(new_n273), .C2(new_n274), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n277), .A2(new_n283), .A3(new_n284), .A4(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT82), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n288), .A2(KEYINPUT82), .A3(new_n289), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g0094(.A(KEYINPUT5), .B(G41), .ZN(new_n295));
  INV_X1    g0095(.A(G41), .ZN(new_n296));
  OAI211_X1 g0096(.A(G1), .B(G13), .C1(new_n259), .C2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n208), .A2(G45), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n295), .A2(new_n297), .A3(G274), .A4(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n289), .B1(new_n299), .B2(new_n295), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n301), .B1(G270), .B2(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(KEYINPUT83), .B1(new_n294), .B2(new_n303), .ZN(new_n304));
  AND3_X1   g0104(.A1(new_n288), .A2(KEYINPUT82), .A3(new_n289), .ZN(new_n305));
  AOI21_X1  g0105(.A(KEYINPUT82), .B1(new_n288), .B2(new_n289), .ZN(new_n306));
  OAI211_X1 g0106(.A(KEYINPUT83), .B(new_n303), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n272), .B1(new_n304), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n302), .A2(G270), .ZN(new_n310));
  AND3_X1   g0110(.A1(new_n310), .A2(G179), .A3(new_n300), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n294), .A2(new_n269), .A3(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n303), .B1(new_n305), .B2(new_n306), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT83), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n270), .B1(new_n315), .B2(new_n307), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n309), .B(new_n312), .C1(new_n316), .C2(KEYINPUT21), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  NOR3_X1   g0118(.A1(new_n252), .A2(new_n209), .A3(G1), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n202), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n257), .B1(new_n208), .B2(G20), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n320), .B1(new_n322), .B2(new_n202), .ZN(new_n323));
  NOR2_X1   g0123(.A1(KEYINPUT8), .A2(G58), .ZN(new_n324));
  INV_X1    g0124(.A(G58), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT65), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT65), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G58), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n324), .B1(new_n329), .B2(KEYINPUT8), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n330), .A2(new_n209), .A3(G33), .ZN(new_n331));
  NOR2_X1   g0131(.A1(G20), .A2(G33), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n323), .B1(new_n334), .B2(new_n257), .ZN(new_n335));
  OR2_X1    g0135(.A1(new_n335), .A2(KEYINPUT9), .ZN(new_n336));
  INV_X1    g0136(.A(G45), .ZN(new_n337));
  AOI21_X1  g0137(.A(G1), .B1(new_n296), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n297), .A2(G274), .A3(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n338), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n297), .ZN(new_n341));
  INV_X1    g0141(.A(G226), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n339), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n282), .B1(new_n279), .B2(new_n280), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n344), .A2(G223), .B1(new_n275), .B2(G77), .ZN(new_n345));
  INV_X1    g0145(.A(G222), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n281), .A2(new_n282), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n343), .B1(new_n348), .B2(new_n289), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(G190), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT71), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(KEYINPUT10), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n335), .A2(KEYINPUT9), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n336), .A2(new_n350), .A3(new_n352), .A4(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(G200), .ZN(new_n355));
  OR3_X1    g0155(.A1(new_n349), .A2(KEYINPUT70), .A3(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(KEYINPUT70), .B1(new_n349), .B2(new_n355), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n351), .A2(KEYINPUT10), .ZN(new_n359));
  OR3_X1    g0159(.A1(new_n354), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n359), .B1(new_n354), .B2(new_n358), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n349), .A2(G169), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT66), .ZN(new_n363));
  OR3_X1    g0163(.A1(new_n362), .A2(new_n363), .A3(new_n335), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n363), .B1(new_n362), .B2(new_n335), .ZN(new_n365));
  INV_X1    g0165(.A(G179), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n349), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n364), .A2(new_n365), .A3(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n360), .A2(new_n361), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n319), .A2(new_n222), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(new_n322), .B2(new_n222), .ZN(new_n371));
  XOR2_X1   g0171(.A(KEYINPUT8), .B(G58), .Z(new_n372));
  AOI22_X1  g0172(.A1(new_n372), .A2(new_n332), .B1(G20), .B2(G77), .ZN(new_n373));
  XNOR2_X1  g0173(.A(KEYINPUT15), .B(G87), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n209), .A2(G33), .ZN(new_n375));
  OR2_X1    g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n258), .B1(new_n373), .B2(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n371), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(G232), .ZN(new_n379));
  OAI22_X1  g0179(.A1(new_n347), .A2(new_n379), .B1(new_n224), .B2(new_n281), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n344), .A2(G238), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n289), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n339), .B1(new_n341), .B2(new_n223), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(KEYINPUT67), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT67), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n339), .B(new_n386), .C1(new_n341), .C2(new_n223), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n383), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(KEYINPUT68), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT68), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n383), .A2(new_n390), .A3(new_n385), .A4(new_n387), .ZN(new_n391));
  AND2_X1   g0191(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(G169), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n378), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n389), .A2(new_n391), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT69), .B1(new_n395), .B2(new_n366), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT69), .ZN(new_n397));
  AOI211_X1 g0197(.A(new_n397), .B(G179), .C1(new_n389), .C2(new_n391), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n394), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n395), .A2(G190), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n389), .A2(new_n391), .A3(G200), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n400), .A2(new_n378), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n369), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT79), .ZN(new_n405));
  INV_X1    g0205(.A(G190), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n339), .B1(new_n341), .B2(new_n379), .ZN(new_n407));
  OAI211_X1 g0207(.A(G223), .B(new_n282), .C1(new_n273), .C2(new_n274), .ZN(new_n408));
  OAI211_X1 g0208(.A(G226), .B(G1698), .C1(new_n273), .C2(new_n274), .ZN(new_n409));
  NAND2_X1  g0209(.A1(G33), .A2(G87), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n297), .B1(new_n411), .B2(KEYINPUT78), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT78), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n408), .A2(new_n409), .A3(new_n413), .A4(new_n410), .ZN(new_n414));
  AOI211_X1 g0214(.A(new_n406), .B(new_n407), .C1(new_n412), .C2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n411), .A2(KEYINPUT78), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n416), .A2(new_n289), .A3(new_n414), .ZN(new_n417));
  INV_X1    g0217(.A(new_n407), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n355), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n405), .B1(new_n415), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n417), .A2(G190), .A3(new_n418), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n407), .B1(new_n412), .B2(new_n414), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n421), .B(KEYINPUT79), .C1(new_n355), .C2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n330), .A2(new_n319), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n425), .B1(new_n330), .B2(new_n322), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT16), .ZN(new_n427));
  INV_X1    g0227(.A(new_n332), .ZN(new_n428));
  INV_X1    g0228(.A(G159), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n201), .B1(new_n329), .B2(G68), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n431), .B1(new_n432), .B2(new_n209), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n279), .A2(new_n209), .A3(new_n280), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT7), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n279), .A2(KEYINPUT7), .A3(new_n209), .A4(new_n280), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n216), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n427), .B1(new_n433), .B2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(KEYINPUT7), .B1(new_n275), .B2(new_n209), .ZN(new_n440));
  INV_X1    g0240(.A(new_n437), .ZN(new_n441));
  OAI21_X1  g0241(.A(G68), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  XNOR2_X1  g0242(.A(KEYINPUT65), .B(G58), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n231), .B1(new_n443), .B2(new_n216), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n430), .B1(new_n444), .B2(G20), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n442), .A2(new_n445), .A3(KEYINPUT16), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n439), .A2(new_n446), .A3(new_n257), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(KEYINPUT77), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT77), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n439), .A2(new_n446), .A3(new_n449), .A4(new_n257), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n426), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n424), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT17), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n422), .A2(new_n393), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n455), .B1(G179), .B2(new_n422), .ZN(new_n456));
  OAI21_X1  g0256(.A(KEYINPUT18), .B1(new_n451), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n448), .A2(new_n450), .ZN(new_n458));
  INV_X1    g0258(.A(new_n426), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT18), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n422), .A2(G179), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n462), .B1(new_n393), .B2(new_n422), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n460), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n424), .A2(KEYINPUT17), .A3(new_n451), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n454), .A2(new_n457), .A3(new_n464), .A4(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n216), .A2(G20), .ZN(new_n468));
  INV_X1    g0268(.A(new_n253), .ZN(new_n469));
  AOI211_X1 g0269(.A(new_n468), .B(new_n469), .C1(KEYINPUT75), .C2(KEYINPUT12), .ZN(new_n470));
  OR2_X1    g0270(.A1(KEYINPUT75), .A2(KEYINPUT12), .ZN(new_n471));
  AND2_X1   g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR3_X1   g0272(.A1(new_n470), .A2(KEYINPUT75), .A3(KEYINPUT12), .ZN(new_n473));
  AOI211_X1 g0273(.A(new_n472), .B(new_n473), .C1(G68), .C2(new_n321), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT13), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n339), .B1(new_n341), .B2(new_n217), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n281), .A2(G226), .A3(new_n282), .ZN(new_n478));
  NAND2_X1  g0278(.A1(G33), .A2(G97), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI211_X1 g0280(.A(G232), .B(G1698), .C1(new_n273), .C2(new_n274), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT72), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n281), .A2(KEYINPUT72), .A3(G232), .A4(G1698), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n480), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n475), .B(new_n477), .C1(new_n485), .C2(new_n297), .ZN(new_n486));
  INV_X1    g0286(.A(new_n479), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n275), .A2(G1698), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n487), .B1(new_n488), .B2(G226), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n483), .A2(new_n484), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n297), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(KEYINPUT13), .B1(new_n491), .B2(new_n476), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n486), .A2(new_n492), .A3(G190), .ZN(new_n493));
  OAI221_X1 g0293(.A(new_n468), .B1(new_n375), .B2(new_n222), .C1(new_n428), .C2(new_n202), .ZN(new_n494));
  XNOR2_X1  g0294(.A(KEYINPUT73), .B(KEYINPUT11), .ZN(new_n495));
  AND3_X1   g0295(.A1(new_n494), .A2(new_n257), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n495), .B1(new_n494), .B2(new_n257), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OR2_X1    g0298(.A1(new_n498), .A2(KEYINPUT74), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(KEYINPUT74), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n474), .A2(new_n493), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n355), .B1(new_n486), .B2(new_n492), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n486), .A2(new_n492), .A3(G179), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(KEYINPUT76), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT76), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n486), .A2(new_n492), .A3(new_n506), .A4(G179), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n492), .ZN(new_n509));
  NOR3_X1   g0309(.A1(new_n491), .A2(KEYINPUT13), .A3(new_n476), .ZN(new_n510));
  OAI21_X1  g0310(.A(G169), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(KEYINPUT14), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT14), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n513), .B(G169), .C1(new_n509), .C2(new_n510), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n508), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n474), .A2(new_n499), .A3(new_n500), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n503), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n404), .A2(new_n467), .A3(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n315), .A2(new_n307), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n269), .B1(new_n520), .B2(G200), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n521), .B1(new_n406), .B2(new_n520), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n209), .B(G87), .C1(new_n273), .C2(new_n274), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(KEYINPUT22), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT22), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n281), .A2(new_n525), .A3(new_n209), .A4(G87), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n224), .A2(G20), .ZN(new_n528));
  INV_X1    g0328(.A(G116), .ZN(new_n529));
  OAI22_X1  g0329(.A1(KEYINPUT23), .A2(new_n528), .B1(new_n375), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT84), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n531), .B(KEYINPUT23), .C1(new_n209), .C2(G107), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n531), .B1(new_n528), .B2(KEYINPUT23), .ZN(new_n534));
  NOR3_X1   g0334(.A1(new_n530), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT24), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n527), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n536), .B1(new_n527), .B2(new_n535), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n257), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT25), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(new_n254), .B2(G107), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n319), .A2(KEYINPUT25), .A3(new_n224), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n261), .A2(G107), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n295), .A2(new_n299), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n546), .A2(G264), .A3(new_n297), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n219), .A2(new_n282), .ZN(new_n548));
  INV_X1    g0348(.A(G257), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G1698), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n548), .B(new_n550), .C1(new_n273), .C2(new_n274), .ZN(new_n551));
  NAND2_X1  g0351(.A1(G33), .A2(G294), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n297), .B1(new_n553), .B2(KEYINPUT85), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT85), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n551), .A2(new_n555), .A3(new_n552), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n547), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n557), .A2(new_n366), .A3(new_n300), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n300), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n393), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n545), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(G200), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n557), .A2(G190), .A3(new_n300), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n562), .A2(new_n540), .A3(new_n544), .A4(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n297), .A2(KEYINPUT80), .A3(G250), .A4(new_n298), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n297), .A2(G274), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n565), .B1(new_n566), .B2(new_n298), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT80), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n297), .A2(G250), .A3(new_n298), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  OAI211_X1 g0370(.A(G244), .B(G1698), .C1(new_n273), .C2(new_n274), .ZN(new_n571));
  OAI211_X1 g0371(.A(G238), .B(new_n282), .C1(new_n273), .C2(new_n274), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n571), .B(new_n572), .C1(new_n259), .C2(new_n529), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n289), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n570), .A2(new_n366), .A3(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n281), .A2(new_n209), .A3(G68), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT19), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n209), .B1(new_n479), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(G87), .B2(new_n206), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n577), .B1(new_n375), .B2(new_n264), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n576), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n581), .A2(new_n257), .B1(new_n319), .B2(new_n374), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(new_n260), .B2(new_n374), .ZN(new_n583));
  INV_X1    g0383(.A(new_n574), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n569), .A2(new_n568), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n585), .B(new_n565), .C1(new_n566), .C2(new_n298), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n575), .B(new_n583), .C1(G169), .C2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(G190), .ZN(new_n589));
  OAI21_X1  g0389(.A(G200), .B1(new_n584), .B2(new_n586), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n261), .A2(G87), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n589), .A2(new_n590), .A3(new_n582), .A4(new_n591), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n561), .A2(new_n564), .A3(new_n588), .A4(new_n592), .ZN(new_n593));
  OAI211_X1 g0393(.A(G244), .B(new_n282), .C1(new_n273), .C2(new_n274), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT4), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n344), .A2(G250), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n281), .A2(KEYINPUT4), .A3(G244), .A4(new_n282), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n596), .A2(new_n597), .A3(new_n598), .A4(new_n263), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n289), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n546), .A2(new_n297), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n300), .B1(new_n601), .B2(new_n549), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(G200), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n602), .B1(new_n289), .B2(new_n599), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(G190), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT6), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n264), .A2(new_n224), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n608), .B1(new_n609), .B2(new_n205), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n224), .A2(KEYINPUT6), .A3(G97), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n612), .A2(G20), .B1(G77), .B2(new_n332), .ZN(new_n613));
  OAI21_X1  g0413(.A(G107), .B1(new_n440), .B2(new_n441), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n257), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n254), .A2(G97), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n617), .B1(new_n261), .B2(G97), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n605), .A2(new_n607), .A3(new_n616), .A4(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n616), .A2(new_n618), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n604), .A2(new_n393), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n606), .A2(new_n366), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n593), .A2(new_n624), .ZN(new_n625));
  AND4_X1   g0425(.A1(new_n318), .A2(new_n519), .A3(new_n522), .A4(new_n625), .ZN(G372));
  INV_X1    g0426(.A(new_n368), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n515), .A2(new_n516), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n399), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n424), .A2(KEYINPUT17), .A3(new_n451), .ZN(new_n630));
  AOI21_X1  g0430(.A(KEYINPUT17), .B1(new_n424), .B2(new_n451), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n503), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n629), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n464), .A2(new_n457), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n360), .A2(new_n361), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n627), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n573), .A2(KEYINPUT86), .A3(new_n289), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(KEYINPUT86), .B1(new_n573), .B2(new_n289), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n570), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n393), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n644), .A2(new_n575), .A3(new_n583), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n582), .A2(new_n591), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT87), .ZN(new_n647));
  XNOR2_X1  g0447(.A(new_n646), .B(new_n647), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n643), .A2(G200), .B1(new_n587), .B2(G190), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n575), .A2(new_n583), .ZN(new_n650));
  AOI22_X1  g0450(.A1(new_n648), .A2(new_n649), .B1(new_n650), .B2(new_n644), .ZN(new_n651));
  INV_X1    g0451(.A(new_n623), .ZN(new_n652));
  AOI21_X1  g0452(.A(KEYINPUT26), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n592), .A2(new_n588), .ZN(new_n654));
  XOR2_X1   g0454(.A(KEYINPUT90), .B(KEYINPUT26), .Z(new_n655));
  NOR3_X1   g0455(.A1(new_n654), .A2(new_n623), .A3(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n645), .B1(new_n653), .B2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n624), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n658), .A2(new_n564), .A3(new_n651), .ZN(new_n659));
  INV_X1    g0459(.A(new_n270), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n660), .B1(new_n304), .B2(new_n308), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(new_n271), .ZN(new_n662));
  AOI211_X1 g0462(.A(new_n301), .B(new_n547), .C1(new_n554), .C2(new_n556), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n558), .B1(new_n663), .B2(G169), .ZN(new_n664));
  INV_X1    g0464(.A(new_n544), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n527), .A2(new_n535), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(KEYINPUT24), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n537), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n665), .B1(new_n668), .B2(new_n257), .ZN(new_n669));
  OAI21_X1  g0469(.A(KEYINPUT88), .B1(new_n664), .B2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT88), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n545), .A2(new_n671), .A3(new_n558), .A4(new_n560), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n312), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n674), .B1(new_n520), .B2(new_n272), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n662), .A2(new_n673), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT89), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n659), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n662), .A2(new_n673), .A3(new_n675), .A4(KEYINPUT89), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n657), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n639), .B1(new_n518), .B2(new_n680), .ZN(G369));
  OR3_X1    g0481(.A1(new_n469), .A2(KEYINPUT27), .A3(G20), .ZN(new_n682));
  OAI21_X1  g0482(.A(KEYINPUT27), .B1(new_n469), .B2(G20), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(G213), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(G343), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n318), .A2(new_n686), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n561), .A2(new_n564), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n670), .A2(new_n672), .ZN(new_n690));
  INV_X1    g0490(.A(new_n686), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(G330), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n269), .A2(new_n686), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n318), .A2(new_n522), .A3(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n317), .A2(new_n269), .A3(new_n686), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n694), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n688), .B1(new_n669), .B2(new_n691), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n561), .B2(new_n691), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n693), .A2(new_n701), .ZN(G399));
  INV_X1    g0502(.A(new_n212), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(G41), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR3_X1   g0505(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n705), .A2(G1), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n707), .B1(new_n232), .B2(new_n705), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n708), .B(KEYINPUT28), .ZN(new_n709));
  XNOR2_X1  g0509(.A(new_n646), .B(KEYINPUT87), .ZN(new_n710));
  INV_X1    g0510(.A(new_n642), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n586), .B1(new_n711), .B2(new_n640), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n589), .B1(new_n712), .B2(new_n355), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n645), .B1(new_n710), .B2(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n564), .A2(new_n623), .A3(new_n619), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n561), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n716), .B1(new_n317), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n645), .A2(KEYINPUT93), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT93), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n650), .A2(new_n720), .A3(new_n644), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n651), .A2(KEYINPUT26), .A3(new_n652), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n655), .B1(new_n654), .B2(new_n623), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n722), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n686), .B1(new_n718), .B2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT29), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n677), .B1(new_n317), .B2(new_n690), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n729), .A2(new_n679), .A3(new_n716), .ZN(new_n730));
  INV_X1    g0530(.A(new_n657), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n686), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n728), .B1(new_n727), .B2(new_n732), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n663), .A2(G179), .A3(new_n606), .ZN(new_n734));
  OAI211_X1 g0534(.A(new_n643), .B(new_n734), .C1(new_n304), .C2(new_n308), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT30), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n606), .B1(new_n305), .B2(new_n306), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n587), .A2(new_n311), .A3(new_n557), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  AND4_X1   g0539(.A1(new_n311), .A2(new_n557), .A3(new_n574), .A4(new_n570), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n740), .A2(KEYINPUT30), .A3(new_n294), .A4(new_n606), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n735), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT31), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n691), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(KEYINPUT91), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n741), .A2(new_n739), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n643), .A2(new_n559), .A3(new_n366), .A4(new_n604), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n747), .B1(new_n315), .B2(new_n307), .ZN(new_n748));
  OAI211_X1 g0548(.A(KEYINPUT91), .B(new_n744), .C1(new_n746), .C2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n745), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(KEYINPUT92), .B1(new_n746), .B2(new_n748), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT92), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n735), .A2(new_n753), .A3(new_n739), .A4(new_n741), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n752), .A2(new_n754), .A3(new_n686), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(new_n743), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n318), .A2(new_n625), .A3(new_n522), .A4(new_n691), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n751), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G330), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n733), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n709), .B1(new_n761), .B2(G1), .ZN(G364));
  NOR2_X1   g0562(.A1(new_n252), .A2(G20), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n208), .B1(new_n763), .B2(G45), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n704), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n698), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n696), .A2(new_n694), .A3(new_n697), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n703), .A2(new_n275), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n770), .A2(G355), .B1(new_n529), .B2(new_n703), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n250), .A2(new_n337), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n703), .A2(new_n281), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n773), .B1(G45), .B2(new_n232), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n771), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  AND2_X1   g0575(.A1(new_n775), .A2(KEYINPUT94), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G13), .A2(G33), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G20), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n228), .B1(G20), .B2(new_n393), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(new_n775), .B2(KEYINPUT94), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n766), .B1(new_n776), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n366), .A2(new_n355), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT96), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n209), .A2(G190), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n787), .A2(KEYINPUT97), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(KEYINPUT97), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G329), .ZN(new_n792));
  NAND3_X1  g0592(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n406), .ZN(new_n794));
  INV_X1    g0594(.A(KEYINPUT95), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NOR3_X1   g0596(.A1(new_n793), .A2(KEYINPUT95), .A3(new_n406), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(G326), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n785), .A2(G190), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n209), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(G294), .ZN(new_n804));
  INV_X1    g0604(.A(G283), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n355), .A2(G179), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n786), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n366), .A2(G200), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n786), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(G311), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n805), .A2(new_n807), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n209), .A2(new_n406), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(new_n806), .ZN(new_n813));
  INV_X1    g0613(.A(G303), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n793), .A2(G190), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  XOR2_X1   g0616(.A(KEYINPUT33), .B(G317), .Z(new_n817));
  OAI221_X1 g0617(.A(new_n275), .B1(new_n813), .B2(new_n814), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n812), .A2(new_n808), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n811), .B(new_n818), .C1(G322), .C2(new_n820), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n792), .A2(new_n800), .A3(new_n804), .A4(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n790), .A2(new_n429), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT98), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(KEYINPUT32), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n803), .A2(G97), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(new_n202), .B2(new_n798), .ZN(new_n827));
  INV_X1    g0627(.A(new_n807), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n329), .A2(new_n820), .B1(new_n828), .B2(G107), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n829), .B1(new_n222), .B2(new_n809), .C1(new_n216), .C2(new_n816), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n281), .B1(new_n813), .B2(new_n218), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT99), .ZN(new_n832));
  NOR3_X1   g0632(.A1(new_n827), .A2(new_n830), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n825), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n824), .A2(KEYINPUT32), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n822), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n783), .B1(new_n836), .B2(new_n780), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n696), .A2(new_n697), .A3(new_n779), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n769), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(G396));
  INV_X1    g0641(.A(new_n766), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n730), .A2(new_n731), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n399), .A2(new_n402), .A3(new_n691), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n691), .A2(new_n378), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n399), .A2(new_n402), .A3(new_n848), .ZN(new_n849));
  OAI22_X1  g0649(.A1(new_n395), .A2(G169), .B1(new_n377), .B2(new_n371), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n397), .B1(new_n392), .B2(G179), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n395), .A2(KEYINPUT69), .A3(new_n366), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n847), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n849), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n846), .B1(new_n732), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n842), .B1(new_n856), .B2(new_n759), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n857), .A2(KEYINPUT100), .B1(new_n759), .B2(new_n856), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(KEYINPUT100), .B2(new_n857), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n780), .A2(new_n777), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n766), .B1(G77), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n813), .ZN(new_n863));
  AOI22_X1  g0663(.A1(G107), .A2(new_n863), .B1(new_n828), .B2(G87), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n864), .B1(new_n529), .B2(new_n809), .ZN(new_n865));
  INV_X1    g0665(.A(G294), .ZN(new_n866));
  OAI221_X1 g0666(.A(new_n275), .B1(new_n819), .B2(new_n866), .C1(new_n805), .C2(new_n816), .ZN(new_n867));
  AOI211_X1 g0667(.A(new_n865), .B(new_n867), .C1(G97), .C2(new_n803), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n868), .B1(new_n814), .B2(new_n798), .C1(new_n810), .C2(new_n790), .ZN(new_n869));
  INV_X1    g0669(.A(new_n809), .ZN(new_n870));
  AOI22_X1  g0670(.A1(G143), .A2(new_n820), .B1(new_n870), .B2(G159), .ZN(new_n871));
  INV_X1    g0671(.A(G150), .ZN(new_n872));
  INV_X1    g0672(.A(G137), .ZN(new_n873));
  OAI221_X1 g0673(.A(new_n871), .B1(new_n872), .B2(new_n816), .C1(new_n798), .C2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT34), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n874), .A2(new_n875), .ZN(new_n877));
  OAI221_X1 g0677(.A(new_n281), .B1(new_n807), .B2(new_n216), .C1(new_n202), .C2(new_n813), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n878), .B1(new_n803), .B2(new_n329), .ZN(new_n879));
  INV_X1    g0679(.A(G132), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n877), .B(new_n879), .C1(new_n880), .C2(new_n790), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n869), .B1(new_n876), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n862), .B1(new_n882), .B2(new_n780), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(new_n855), .B2(new_n778), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n859), .A2(new_n884), .ZN(G384));
  AND2_X1   g0685(.A1(new_n612), .A2(KEYINPUT35), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n612), .A2(KEYINPUT35), .ZN(new_n887));
  NOR4_X1   g0687(.A1(new_n886), .A2(new_n887), .A3(new_n529), .A4(new_n230), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n888), .B(KEYINPUT36), .ZN(new_n889));
  INV_X1    g0689(.A(new_n232), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n890), .B(G77), .C1(new_n216), .C2(new_n443), .ZN(new_n891));
  AOI211_X1 g0691(.A(new_n208), .B(G13), .C1(new_n891), .C2(new_n246), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n447), .A2(new_n459), .ZN(new_n894));
  INV_X1    g0694(.A(new_n684), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n466), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n684), .B(KEYINPUT102), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT37), .B1(new_n460), .B2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT101), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n460), .A2(new_n902), .A3(new_n463), .ZN(new_n903));
  OAI21_X1  g0703(.A(KEYINPUT101), .B1(new_n451), .B2(new_n456), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n901), .A2(new_n903), .A3(new_n452), .A4(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n894), .B1(new_n463), .B2(new_n895), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n452), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(KEYINPUT37), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  AND3_X1   g0709(.A1(new_n898), .A2(KEYINPUT38), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT38), .B1(new_n898), .B2(new_n909), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT39), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n898), .A2(KEYINPUT38), .A3(new_n909), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n451), .A2(new_n899), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n424), .A2(new_n451), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n451), .B1(new_n456), .B2(new_n899), .ZN(new_n917));
  OAI21_X1  g0717(.A(KEYINPUT37), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n466), .A2(new_n915), .B1(new_n918), .B2(new_n905), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n914), .B1(new_n919), .B2(KEYINPUT38), .ZN(new_n920));
  XNOR2_X1  g0720(.A(KEYINPUT103), .B(KEYINPUT39), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  OAI22_X1  g0722(.A1(new_n912), .A2(new_n913), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n515), .A2(new_n516), .A3(new_n691), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n635), .A2(new_n900), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n516), .A2(new_n686), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n628), .A2(new_n633), .A3(new_n928), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n516), .B(new_n686), .C1(new_n515), .C2(new_n503), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n399), .A2(new_n686), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n931), .B1(new_n846), .B2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT38), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n896), .B1(new_n635), .B2(new_n632), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT37), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(new_n452), .B2(new_n906), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n902), .B1(new_n460), .B2(new_n463), .ZN(new_n939));
  NOR3_X1   g0739(.A1(new_n451), .A2(new_n456), .A3(KEYINPUT101), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n937), .B1(new_n451), .B2(new_n899), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n916), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n938), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n935), .B1(new_n936), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n914), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n927), .B1(new_n934), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n926), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n732), .A2(new_n727), .ZN(new_n949));
  INV_X1    g0749(.A(new_n728), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n518), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n639), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n948), .B(new_n953), .ZN(new_n954));
  NAND4_X1  g0754(.A1(new_n752), .A2(new_n754), .A3(KEYINPUT31), .A4(new_n686), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n756), .A2(new_n757), .A3(new_n955), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n929), .A2(new_n930), .B1(new_n849), .B2(new_n854), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT40), .ZN(new_n958));
  AND3_X1   g0758(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n946), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n466), .A2(new_n915), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n918), .A2(new_n905), .ZN(new_n962));
  AOI21_X1  g0762(.A(KEYINPUT38), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n910), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n956), .A2(new_n957), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n960), .B1(new_n966), .B2(new_n958), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n519), .A2(new_n956), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n967), .A2(new_n968), .ZN(new_n970));
  NOR3_X1   g0770(.A1(new_n969), .A2(new_n970), .A3(new_n694), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n954), .A2(new_n971), .B1(new_n208), .B2(new_n763), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n954), .A2(new_n971), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n893), .B1(new_n972), .B2(new_n973), .ZN(G367));
  NAND2_X1  g0774(.A1(new_n620), .A2(new_n686), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n658), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n652), .A2(new_n686), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n689), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT42), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n648), .A2(new_n691), .ZN(new_n982));
  INV_X1    g0782(.A(new_n645), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n984), .B1(new_n714), .B2(new_n982), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n985), .A2(KEYINPUT43), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n623), .B1(new_n976), .B2(new_n561), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n691), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n981), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT104), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n981), .A2(KEYINPUT104), .A3(new_n986), .A4(new_n988), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n981), .A2(new_n988), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n985), .A2(KEYINPUT43), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n985), .A2(KEYINPUT43), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n994), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n993), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n701), .B2(new_n979), .ZN(new_n999));
  INV_X1    g0799(.A(new_n701), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n993), .A2(new_n1000), .A3(new_n978), .A4(new_n997), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n704), .B(KEYINPUT41), .Z(new_n1002));
  INV_X1    g0802(.A(KEYINPUT44), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n693), .B2(new_n978), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n689), .A2(new_n692), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1005), .A2(KEYINPUT44), .A3(new_n979), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1005), .A2(new_n979), .ZN(new_n1008));
  AND2_X1   g0808(.A1(new_n1008), .A2(KEYINPUT45), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1008), .A2(KEYINPUT45), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1007), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n1000), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n689), .B1(new_n700), .B2(new_n687), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(new_n698), .ZN(new_n1014));
  AND2_X1   g0814(.A1(new_n761), .A2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1008), .B(KEYINPUT45), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1016), .A2(new_n701), .A3(new_n1007), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1012), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1002), .B1(new_n1018), .B2(new_n761), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n999), .B(new_n1001), .C1(new_n1019), .C2(new_n765), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n781), .B1(new_n212), .B2(new_n374), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(new_n773), .B2(new_n241), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n791), .A2(G137), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n802), .A2(new_n216), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n799), .A2(G143), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n813), .A2(new_n443), .B1(new_n809), .B2(new_n202), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n281), .B1(new_n819), .B2(new_n872), .C1(new_n429), .C2(new_n816), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n1027), .B(new_n1028), .C1(G77), .C2(new_n828), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1023), .A2(new_n1025), .A3(new_n1026), .A4(new_n1029), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n802), .A2(new_n224), .B1(new_n805), .B2(new_n809), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT105), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT46), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n813), .B2(new_n529), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n816), .B2(new_n866), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n275), .B1(new_n807), .B2(new_n264), .C1(new_n814), .C2(new_n819), .ZN(new_n1036));
  NOR3_X1   g0836(.A1(new_n813), .A2(new_n1033), .A3(new_n529), .ZN(new_n1037));
  NOR3_X1   g0837(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(G317), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1038), .B1(new_n810), .B2(new_n798), .C1(new_n790), .C2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1030), .B1(new_n1032), .B2(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT47), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n842), .B(new_n1022), .C1(new_n1042), .C2(new_n780), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n779), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n985), .A2(new_n1044), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1020), .A2(new_n1047), .ZN(G387));
  NAND2_X1  g0848(.A1(new_n1014), .A2(new_n765), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT106), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n802), .A2(new_n374), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(new_n799), .B2(G159), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n791), .A2(G150), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n330), .A2(new_n815), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n281), .B1(new_n807), .B2(new_n264), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n202), .A2(new_n819), .B1(new_n813), .B2(new_n222), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n1055), .B(new_n1056), .C1(G68), .C2(new_n870), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .A4(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n791), .A2(G326), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n281), .B1(new_n828), .B2(G116), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n802), .A2(new_n805), .B1(new_n866), .B2(new_n813), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n819), .A2(new_n1039), .B1(new_n809), .B2(new_n814), .ZN(new_n1062));
  XOR2_X1   g0862(.A(new_n1062), .B(KEYINPUT107), .Z(new_n1063));
  INV_X1    g0863(.A(G322), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n1063), .B1(new_n810), .B2(new_n816), .C1(new_n1064), .C2(new_n798), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT48), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1061), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n1066), .B2(new_n1065), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT49), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1059), .B(new_n1060), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1070));
  AND2_X1   g0870(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1058), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n780), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n706), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n770), .A2(new_n1074), .B1(new_n224), .B2(new_n703), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n238), .A2(new_n337), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n372), .A2(new_n202), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT50), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n706), .B(new_n337), .C1(new_n216), .C2(new_n222), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n773), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1075), .B1(new_n1076), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n842), .B1(new_n1081), .B2(new_n781), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1073), .B(new_n1082), .C1(new_n700), .C2(new_n1044), .ZN(new_n1083));
  AND2_X1   g0883(.A1(new_n1050), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n761), .A2(new_n1014), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n704), .B(KEYINPUT108), .Z(new_n1086));
  NOR2_X1   g0886(.A1(new_n761), .A2(new_n1014), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1085), .B(new_n1086), .C1(new_n1087), .C2(KEYINPUT109), .ZN(new_n1088));
  AND2_X1   g0888(.A1(new_n1087), .A2(KEYINPUT109), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1084), .B1(new_n1088), .B2(new_n1089), .ZN(G393));
  INV_X1    g0890(.A(KEYINPUT110), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1012), .A2(new_n1091), .A3(new_n1017), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1016), .A2(KEYINPUT110), .A3(new_n701), .A4(new_n1007), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1018), .B(new_n1086), .C1(new_n1094), .C2(new_n1015), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n281), .B1(new_n807), .B2(new_n218), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n372), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n1097), .A2(new_n809), .B1(new_n216), .B2(new_n813), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n1096), .B(new_n1098), .C1(G50), .C2(new_n815), .ZN(new_n1099));
  INV_X1    g0899(.A(G143), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n1099), .B1(new_n222), .B2(new_n802), .C1(new_n1100), .C2(new_n790), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n798), .A2(new_n872), .B1(new_n429), .B2(new_n819), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT51), .Z(new_n1103));
  OAI21_X1  g0903(.A(new_n275), .B1(new_n807), .B2(new_n224), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n813), .A2(new_n805), .B1(new_n809), .B2(new_n866), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n1104), .B(new_n1105), .C1(G303), .C2(new_n815), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n1106), .B1(new_n529), .B2(new_n802), .C1(new_n790), .C2(new_n1064), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n798), .A2(new_n1039), .B1(new_n810), .B2(new_n819), .ZN(new_n1108));
  XOR2_X1   g0908(.A(new_n1108), .B(KEYINPUT52), .Z(new_n1109));
  OAI22_X1  g0909(.A1(new_n1101), .A2(new_n1103), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n780), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n773), .ZN(new_n1112));
  OAI221_X1 g0912(.A(new_n781), .B1(new_n264), .B2(new_n212), .C1(new_n1112), .C2(new_n245), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1111), .A2(new_n766), .A3(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(new_n979), .B2(new_n779), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(new_n1094), .B2(new_n765), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1095), .A2(new_n1116), .ZN(G390));
  AOI21_X1  g0917(.A(new_n932), .B1(new_n726), .B2(new_n855), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n920), .B(new_n924), .C1(new_n1118), .C2(new_n931), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n929), .A2(new_n930), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n758), .A2(G330), .A3(new_n855), .A4(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n933), .B1(new_n680), .B2(new_n844), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n925), .B1(new_n1122), .B2(new_n1120), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1119), .B(new_n1121), .C1(new_n923), .C2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n924), .B1(new_n910), .B2(new_n963), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n718), .A2(new_n725), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1126), .A2(new_n855), .A3(new_n691), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n931), .B1(new_n1127), .B2(new_n933), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1125), .A2(new_n1128), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n964), .A2(new_n921), .B1(new_n946), .B2(KEYINPUT39), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n844), .B1(new_n730), .B2(new_n731), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1120), .B1(new_n1131), .B2(new_n932), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n924), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1129), .B1(new_n1130), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n956), .A2(new_n957), .A3(G330), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1124), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n956), .A2(G330), .A3(new_n855), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n931), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1138), .A2(new_n1118), .A3(new_n1121), .ZN(new_n1139));
  AND2_X1   g0939(.A1(new_n956), .A2(G330), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n758), .A2(G330), .A3(new_n855), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n957), .A2(new_n1140), .B1(new_n1141), .B2(new_n931), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1122), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1139), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n519), .A2(G330), .A3(new_n956), .ZN(new_n1145));
  NOR3_X1   g0945(.A1(new_n951), .A2(new_n1145), .A3(new_n952), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(KEYINPUT111), .B1(new_n1136), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1140), .A2(new_n519), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1149), .B(new_n639), .C1(new_n733), .C2(new_n518), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n1141), .A2(new_n931), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1135), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1122), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1150), .B1(new_n1153), .B2(new_n1139), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT111), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1119), .B1(new_n923), .B2(new_n1123), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(new_n1152), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1154), .A2(new_n1155), .A3(new_n1157), .A4(new_n1124), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1148), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1086), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(new_n1136), .B2(new_n1147), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT114), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1136), .A2(new_n764), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1130), .A2(new_n777), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n766), .B1(new_n330), .B2(new_n861), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n802), .A2(new_n222), .B1(new_n529), .B2(new_n819), .ZN(new_n1167));
  XOR2_X1   g0967(.A(new_n1167), .B(KEYINPUT113), .Z(new_n1168));
  AOI22_X1  g0968(.A1(new_n870), .A2(G97), .B1(G107), .B2(new_n815), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1169), .B1(new_n798), .B2(new_n805), .ZN(new_n1170));
  XOR2_X1   g0970(.A(new_n1170), .B(KEYINPUT112), .Z(new_n1171));
  OAI221_X1 g0971(.A(new_n275), .B1(new_n807), .B2(new_n216), .C1(new_n218), .C2(new_n813), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(new_n791), .B2(G294), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1168), .A2(new_n1171), .A3(new_n1173), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n803), .A2(G159), .B1(G128), .B2(new_n799), .ZN(new_n1175));
  OR3_X1    g0975(.A1(new_n813), .A2(KEYINPUT53), .A3(new_n872), .ZN(new_n1176));
  OAI21_X1  g0976(.A(KEYINPUT53), .B1(new_n813), .B2(new_n872), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1176), .B(new_n1177), .C1(new_n816), .C2(new_n873), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(KEYINPUT54), .B(G143), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n281), .B1(new_n809), .B2(new_n1179), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n819), .A2(new_n880), .B1(new_n807), .B2(new_n202), .ZN(new_n1181));
  NOR3_X1   g0981(.A1(new_n1178), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(G125), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1175), .B(new_n1182), .C1(new_n1183), .C2(new_n790), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1174), .A2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1166), .B1(new_n1185), .B2(new_n780), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1164), .B1(new_n1165), .B2(new_n1186), .ZN(new_n1187));
  AND3_X1   g0987(.A1(new_n1162), .A2(new_n1163), .A3(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1163), .B1(new_n1162), .B2(new_n1187), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1188), .A2(new_n1189), .ZN(G378));
  NOR2_X1   g0990(.A1(new_n335), .A2(new_n684), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1191), .B(KEYINPUT115), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n369), .B(new_n1192), .ZN(new_n1193));
  XOR2_X1   g0993(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1194));
  XNOR2_X1  g0994(.A(new_n1193), .B(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n964), .A2(new_n921), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n946), .A2(KEYINPUT39), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n924), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n1132), .A2(new_n912), .B1(new_n635), .B2(new_n900), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n967), .B(G330), .C1(new_n1198), .C2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n920), .A2(new_n956), .A3(new_n957), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1201), .A2(KEYINPUT40), .B1(new_n959), .B2(new_n946), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n926), .B(new_n947), .C1(new_n1202), .C2(new_n694), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1195), .B1(new_n1200), .B2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1200), .A2(new_n1203), .A3(new_n1195), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n1159), .A2(new_n1146), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1160), .B1(new_n1207), .B2(KEYINPUT57), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT57), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1150), .B1(new_n1148), .B2(new_n1158), .ZN(new_n1210));
  AND3_X1   g1010(.A1(new_n1200), .A2(new_n1203), .A3(new_n1195), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1211), .A2(new_n1204), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1209), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(KEYINPUT116), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT116), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1215), .B(new_n1209), .C1(new_n1210), .C2(new_n1212), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1208), .A2(new_n1214), .A3(new_n1216), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n765), .B1(new_n1211), .B2(new_n1204), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n281), .A2(G41), .ZN(new_n1219));
  AOI211_X1 g1019(.A(G50), .B(new_n1219), .C1(new_n259), .C2(new_n296), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1219), .B1(new_n222), .B2(new_n813), .C1(new_n816), .C2(new_n264), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n809), .A2(new_n374), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n819), .A2(new_n224), .B1(new_n807), .B2(new_n443), .ZN(new_n1223));
  NOR4_X1   g1023(.A1(new_n1024), .A2(new_n1221), .A3(new_n1222), .A4(new_n1223), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1224), .B1(new_n529), .B2(new_n798), .C1(new_n805), .C2(new_n790), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT58), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1220), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n809), .A2(new_n873), .ZN(new_n1228));
  INV_X1    g1028(.A(G128), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n1229), .A2(new_n819), .B1(new_n813), .B2(new_n1179), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n1228), .B(new_n1230), .C1(G132), .C2(new_n815), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1231), .B1(new_n1183), .B2(new_n798), .C1(new_n872), .C2(new_n802), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1232), .A2(KEYINPUT59), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(KEYINPUT59), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n259), .B(new_n296), .C1(new_n807), .C2(new_n429), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(new_n791), .B2(G124), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1234), .A2(new_n1236), .ZN(new_n1237));
  OAI221_X1 g1037(.A(new_n1227), .B1(new_n1226), .B2(new_n1225), .C1(new_n1233), .C2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(new_n780), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n842), .B1(new_n202), .B2(new_n860), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1195), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1239), .B(new_n1240), .C1(new_n1241), .C2(new_n778), .ZN(new_n1242));
  AND2_X1   g1042(.A1(new_n1218), .A2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1217), .A2(new_n1243), .ZN(G375));
  XOR2_X1   g1044(.A(new_n764), .B(KEYINPUT118), .Z(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1144), .A2(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n766), .B1(G68), .B2(new_n861), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n802), .A2(new_n202), .ZN(new_n1249));
  OAI221_X1 g1049(.A(new_n281), .B1(new_n807), .B2(new_n443), .C1(new_n816), .C2(new_n1179), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n819), .A2(new_n873), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n813), .A2(new_n429), .B1(new_n809), .B2(new_n872), .ZN(new_n1252));
  NOR4_X1   g1052(.A1(new_n1249), .A2(new_n1250), .A3(new_n1251), .A4(new_n1252), .ZN(new_n1253));
  OAI221_X1 g1053(.A(new_n1253), .B1(new_n1229), .B2(new_n790), .C1(new_n880), .C2(new_n798), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n790), .A2(new_n814), .B1(new_n264), .B2(new_n813), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(new_n1255), .B(KEYINPUT119), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(G283), .A2(new_n820), .B1(new_n870), .B2(G107), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n281), .B1(new_n828), .B2(G77), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1257), .B(new_n1258), .C1(new_n529), .C2(new_n816), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1051), .A2(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1260), .B1(new_n866), .B2(new_n798), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1254), .B1(new_n1256), .B2(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1248), .B1(new_n1262), .B2(new_n780), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1263), .B1(new_n1120), .B2(new_n778), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1247), .A2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(KEYINPUT120), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT120), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1247), .A2(new_n1267), .A3(new_n1264), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1266), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT117), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1270), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1153), .A2(new_n1150), .A3(KEYINPUT117), .A4(new_n1139), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  OR2_X1    g1073(.A1(new_n1154), .A2(new_n1002), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1269), .B1(new_n1273), .B2(new_n1274), .ZN(G381));
  AND2_X1   g1075(.A1(new_n1095), .A2(new_n1116), .ZN(new_n1276));
  INV_X1    g1076(.A(G384), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1084), .B(new_n840), .C1(new_n1089), .C2(new_n1088), .ZN(new_n1279));
  NOR4_X1   g1079(.A1(new_n1278), .A2(G381), .A3(G387), .A4(new_n1279), .ZN(new_n1280));
  AND2_X1   g1080(.A1(new_n1162), .A2(new_n1187), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1280), .A2(new_n1281), .A3(new_n1217), .A4(new_n1243), .ZN(G407));
  NAND2_X1  g1082(.A1(new_n685), .A2(G213), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1281), .A2(new_n1284), .ZN(new_n1285));
  OAI211_X1 g1085(.A(G407), .B(G213), .C1(G375), .C2(new_n1285), .ZN(G409));
  NAND3_X1  g1086(.A1(new_n1217), .A2(G378), .A3(new_n1243), .ZN(new_n1287));
  NOR3_X1   g1087(.A1(new_n1210), .A2(new_n1212), .A3(new_n1002), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1242), .B1(new_n1212), .B2(new_n1245), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1281), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1287), .A2(new_n1290), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1153), .A2(new_n1150), .A3(KEYINPUT60), .A4(new_n1139), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT60), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1154), .A2(new_n1293), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1086), .B(new_n1292), .C1(new_n1273), .C2(new_n1294), .ZN(new_n1295));
  AND3_X1   g1095(.A1(new_n1295), .A2(G384), .A3(new_n1269), .ZN(new_n1296));
  AOI21_X1  g1096(.A(G384), .B1(new_n1295), .B2(new_n1269), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1291), .A2(new_n1283), .A3(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(KEYINPUT62), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1291), .A2(new_n1283), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1295), .A2(new_n1269), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n1277), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1295), .A2(G384), .A3(new_n1269), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  OAI211_X1 g1105(.A(G2897), .B(new_n1284), .C1(new_n1305), .C2(KEYINPUT122), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT123), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1307), .B1(new_n1305), .B2(KEYINPUT122), .ZN(new_n1308));
  OAI211_X1 g1108(.A(KEYINPUT122), .B(new_n1307), .C1(new_n1296), .C2(new_n1297), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1306), .B1(new_n1308), .B2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT122), .ZN(new_n1312));
  OAI21_X1  g1112(.A(KEYINPUT123), .B1(new_n1298), .B2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1284), .A2(G2897), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1314), .B1(new_n1298), .B2(new_n1312), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1313), .A2(new_n1315), .A3(new_n1309), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1311), .A2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1301), .A2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT61), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1284), .B1(new_n1287), .B2(new_n1290), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT62), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1320), .A2(new_n1321), .A3(new_n1298), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1300), .A2(new_n1318), .A3(new_n1319), .A4(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(G387), .A2(new_n1276), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(G390), .A2(new_n1020), .A3(new_n1047), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1324), .A2(KEYINPUT124), .A3(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(G393), .A2(G396), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1327), .A2(new_n1279), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT124), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(G390), .A2(new_n1330), .A3(new_n1020), .A4(new_n1047), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1326), .A2(new_n1329), .A3(new_n1331), .ZN(new_n1332));
  AND2_X1   g1132(.A1(new_n1325), .A2(new_n1328), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT125), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1324), .A2(new_n1334), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(G387), .A2(new_n1276), .A3(KEYINPUT125), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1333), .A2(new_n1335), .A3(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1332), .A2(new_n1337), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1323), .A2(new_n1339), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT121), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1301), .A2(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1320), .A2(KEYINPUT121), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1342), .A2(new_n1317), .A3(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1338), .A2(new_n1319), .ZN(new_n1345));
  INV_X1    g1145(.A(KEYINPUT63), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1345), .B1(new_n1299), .B2(new_n1346), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1320), .A2(KEYINPUT63), .A3(new_n1298), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1344), .A2(new_n1347), .A3(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1340), .A2(new_n1349), .ZN(G405));
  XNOR2_X1  g1150(.A(new_n1338), .B(new_n1298), .ZN(new_n1351));
  AND3_X1   g1151(.A1(G375), .A2(KEYINPUT126), .A3(new_n1281), .ZN(new_n1352));
  AOI21_X1  g1152(.A(KEYINPUT126), .B1(G375), .B2(new_n1281), .ZN(new_n1353));
  INV_X1    g1153(.A(new_n1287), .ZN(new_n1354));
  NOR3_X1   g1154(.A1(new_n1352), .A2(new_n1353), .A3(new_n1354), .ZN(new_n1355));
  XNOR2_X1  g1155(.A(new_n1351), .B(new_n1355), .ZN(G402));
endmodule


