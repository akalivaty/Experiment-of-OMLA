//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 0 0 1 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 0 0 1 0 1 1 1 1 1 1 1 1 1 0 1 1 1 1 1 1 1 1 0 1 0 1 1 0 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:27 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n554, new_n555, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n568, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n600, new_n601, new_n604,
    new_n606, new_n607, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1067, new_n1068, new_n1069;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT67), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n453), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(G567), .A2(new_n456), .B1(new_n453), .B2(G2106), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G101), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(new_n460), .ZN(new_n465));
  INV_X1    g040(.A(G137), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n464), .A2(G125), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n460), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n467), .A2(new_n470), .ZN(G160));
  OAI21_X1  g046(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n472));
  INV_X1    g047(.A(G112), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n472), .B1(new_n473), .B2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n464), .A2(G2105), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT68), .ZN(new_n478));
  INV_X1    g053(.A(new_n465), .ZN(new_n479));
  AOI211_X1 g054(.A(new_n474), .B(new_n478), .C1(G136), .C2(new_n479), .ZN(G162));
  AND2_X1   g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  NOR2_X1   g056(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n482));
  OAI211_X1 g057(.A(G138), .B(new_n460), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(KEYINPUT4), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n485));
  NAND4_X1  g060(.A1(new_n464), .A2(new_n485), .A3(G138), .A4(new_n460), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g062(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(G114), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n488), .B1(new_n489), .B2(G2105), .ZN(new_n490));
  AND2_X1   g065(.A1(G126), .A2(G2105), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n491), .B1(new_n481), .B2(new_n482), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT69), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT69), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n494), .B(new_n491), .C1(new_n481), .C2(new_n482), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n490), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n487), .B1(new_n496), .B2(KEYINPUT70), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT70), .ZN(new_n498));
  AOI211_X1 g073(.A(new_n498), .B(new_n490), .C1(new_n493), .C2(new_n495), .ZN(new_n499));
  OAI21_X1  g074(.A(KEYINPUT71), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n490), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n494), .B1(new_n464), .B2(new_n491), .ZN(new_n502));
  INV_X1    g077(.A(new_n495), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(new_n498), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n496), .A2(KEYINPUT70), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT71), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n505), .A2(new_n506), .A3(new_n507), .A4(new_n487), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n500), .A2(new_n508), .ZN(G164));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT5), .B(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n510), .A2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G50), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n516), .A2(new_n519), .ZN(G166));
  NAND3_X1  g095(.A1(new_n511), .A2(G63), .A3(G651), .ZN(new_n521));
  INV_X1    g096(.A(new_n514), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G51), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT72), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  INV_X1    g101(.A(G89), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n526), .B1(new_n527), .B2(new_n512), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT73), .ZN(new_n529));
  OAI211_X1 g104(.A(new_n521), .B(new_n523), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  AND2_X1   g105(.A1(new_n528), .A2(new_n529), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n530), .A2(new_n531), .ZN(G168));
  NAND2_X1  g107(.A1(G77), .A2(G543), .ZN(new_n533));
  INV_X1    g108(.A(new_n511), .ZN(new_n534));
  INV_X1    g109(.A(G64), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT74), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n518), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n538), .B1(new_n537), .B2(new_n536), .ZN(new_n539));
  INV_X1    g114(.A(new_n512), .ZN(new_n540));
  AOI22_X1  g115(.A1(G90), .A2(new_n540), .B1(new_n522), .B2(G52), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n539), .A2(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  AND2_X1   g118(.A1(new_n511), .A2(G56), .ZN(new_n544));
  AND2_X1   g119(.A1(G68), .A2(G543), .ZN(new_n545));
  OAI21_X1  g120(.A(G651), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(KEYINPUT75), .ZN(new_n547));
  AOI22_X1  g122(.A1(G81), .A2(new_n540), .B1(new_n522), .B2(G43), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n546), .A2(KEYINPUT75), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  NAND2_X1  g131(.A1(new_n522), .A2(G53), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT9), .ZN(new_n558));
  XNOR2_X1  g133(.A(KEYINPUT76), .B(G65), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n511), .A2(new_n559), .B1(G78), .B2(G543), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT77), .ZN(new_n561));
  OR2_X1    g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n518), .B1(new_n560), .B2(new_n561), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n562), .A2(new_n563), .B1(G91), .B2(new_n540), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n558), .A2(new_n564), .ZN(G299));
  INV_X1    g140(.A(G168), .ZN(G286));
  INV_X1    g141(.A(G166), .ZN(G303));
  NAND2_X1  g142(.A1(new_n540), .A2(G87), .ZN(new_n568));
  XOR2_X1   g143(.A(new_n568), .B(KEYINPUT78), .Z(new_n569));
  OR2_X1    g144(.A1(new_n511), .A2(G74), .ZN(new_n570));
  AOI22_X1  g145(.A1(G49), .A2(new_n522), .B1(new_n570), .B2(G651), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n571), .ZN(G288));
  AOI21_X1  g147(.A(KEYINPUT79), .B1(new_n511), .B2(G61), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n573), .B1(G73), .B2(G543), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n511), .A2(KEYINPUT79), .A3(G61), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n518), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(G86), .ZN(new_n577));
  INV_X1    g152(.A(G48), .ZN(new_n578));
  OAI22_X1  g153(.A1(new_n512), .A2(new_n577), .B1(new_n514), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G305));
  INV_X1    g156(.A(G85), .ZN(new_n582));
  INV_X1    g157(.A(G47), .ZN(new_n583));
  OAI22_X1  g158(.A1(new_n512), .A2(new_n582), .B1(new_n514), .B2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n585), .A2(new_n518), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G290));
  NAND2_X1  g163(.A1(G301), .A2(G868), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n540), .A2(G92), .ZN(new_n590));
  XOR2_X1   g165(.A(new_n590), .B(KEYINPUT10), .Z(new_n591));
  NAND2_X1  g166(.A1(G79), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G66), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n534), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n594), .A2(G651), .B1(new_n522), .B2(G54), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n589), .B1(new_n597), .B2(G868), .ZN(G321));
  XNOR2_X1  g173(.A(G321), .B(KEYINPUT80), .ZN(G284));
  INV_X1    g174(.A(G868), .ZN(new_n600));
  NAND2_X1  g175(.A1(G299), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(G168), .B2(new_n600), .ZN(G297));
  OAI21_X1  g177(.A(new_n601), .B1(G168), .B2(new_n600), .ZN(G280));
  INV_X1    g178(.A(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n597), .B1(new_n604), .B2(G860), .ZN(G148));
  INV_X1    g180(.A(new_n551), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(new_n600), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n596), .A2(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(new_n600), .ZN(G323));
  XNOR2_X1  g184(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g185(.A1(new_n476), .A2(G123), .ZN(new_n611));
  XOR2_X1   g186(.A(new_n611), .B(KEYINPUT81), .Z(new_n612));
  NAND2_X1  g187(.A1(new_n479), .A2(G135), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n460), .A2(G111), .ZN(new_n614));
  OAI21_X1  g189(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n615));
  OAI211_X1 g190(.A(new_n612), .B(new_n613), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT82), .Z(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(G2096), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n464), .A2(new_n462), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT13), .B(G2100), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n618), .A2(new_n622), .ZN(G156));
  XOR2_X1   g198(.A(G2451), .B(G2454), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT16), .ZN(new_n625));
  XNOR2_X1  g200(.A(G1341), .B(G1348), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(KEYINPUT14), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2427), .B(G2438), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2430), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT15), .B(G2435), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n628), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(new_n631), .B2(new_n630), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n627), .B(new_n633), .Z(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2443), .B(G2446), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  OAI21_X1  g212(.A(G14), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n638), .B1(new_n637), .B2(new_n635), .ZN(G401));
  XNOR2_X1  g214(.A(G2084), .B(G2090), .ZN(new_n640));
  XOR2_X1   g215(.A(G2072), .B(G2078), .Z(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT83), .Z(new_n642));
  XNOR2_X1  g217(.A(G2067), .B(G2678), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n642), .B(KEYINPUT17), .Z(new_n645));
  INV_X1    g220(.A(new_n643), .ZN(new_n646));
  OAI211_X1 g221(.A(new_n640), .B(new_n644), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n646), .A2(new_n640), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n642), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT18), .Z(new_n650));
  NOR2_X1   g225(.A1(new_n643), .A2(new_n640), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n645), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n647), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2096), .B(G2100), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(G227));
  XNOR2_X1  g231(.A(G1971), .B(G1976), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT19), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1956), .B(G2474), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1961), .B(G1966), .ZN(new_n660));
  NOR3_X1   g235(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT84), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n662), .A2(KEYINPUT20), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(KEYINPUT20), .ZN(new_n664));
  AND2_X1   g239(.A1(new_n659), .A2(new_n660), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n659), .A2(new_n660), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n665), .B1(new_n658), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n658), .A2(KEYINPUT85), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n663), .A2(new_n664), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G1991), .B(G1996), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G1981), .B(G1986), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT86), .ZN(new_n674));
  XOR2_X1   g249(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n672), .B(new_n676), .ZN(G229));
  INV_X1    g252(.A(G16), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(G22), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT89), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(G303), .B2(G16), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(G1971), .Z(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT33), .B(G1976), .ZN(new_n683));
  NOR2_X1   g258(.A1(G16), .A2(G23), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT88), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n685), .B1(G288), .B2(new_n678), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n682), .B1(new_n683), .B2(new_n686), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(new_n683), .B2(new_n686), .ZN(new_n688));
  NOR2_X1   g263(.A1(G6), .A2(G16), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(new_n580), .B2(G16), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT32), .B(G1981), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT90), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT34), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n694), .A2(new_n695), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n587), .A2(new_n678), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(new_n678), .B2(G24), .ZN(new_n699));
  INV_X1    g274(.A(G1986), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n699), .A2(new_n700), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n479), .A2(G131), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n476), .A2(G119), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n460), .A2(G107), .ZN(new_n705));
  OAI21_X1  g280(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n703), .B(new_n704), .C1(new_n705), .C2(new_n706), .ZN(new_n707));
  MUX2_X1   g282(.A(G25), .B(new_n707), .S(G29), .Z(new_n708));
  XOR2_X1   g283(.A(KEYINPUT35), .B(G1991), .Z(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n708), .B(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT87), .ZN(new_n712));
  OAI211_X1 g287(.A(new_n701), .B(new_n702), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(new_n712), .B2(new_n711), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n696), .A2(new_n697), .A3(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT91), .B(KEYINPUT36), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G29), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G27), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT96), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G164), .B2(new_n718), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT97), .Z(new_n722));
  INV_X1    g297(.A(G2078), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n479), .A2(G139), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT95), .Z(new_n726));
  XOR2_X1   g301(.A(KEYINPUT94), .B(KEYINPUT25), .Z(new_n727));
  NAND3_X1  g302(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n726), .B(new_n729), .C1(new_n460), .C2(new_n730), .ZN(new_n731));
  MUX2_X1   g306(.A(G33), .B(new_n731), .S(G29), .Z(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(G2072), .Z(new_n733));
  NAND2_X1  g308(.A1(new_n718), .A2(G26), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT28), .ZN(new_n735));
  OR2_X1    g310(.A1(G104), .A2(G2105), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n736), .B(G2104), .C1(G116), .C2(new_n460), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT93), .Z(new_n738));
  AOI22_X1  g313(.A1(G128), .A2(new_n476), .B1(new_n479), .B2(G140), .ZN(new_n739));
  AND2_X1   g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n735), .B1(new_n740), .B2(new_n718), .ZN(new_n741));
  INV_X1    g316(.A(G2067), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(G4), .A2(G16), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(new_n597), .B2(G16), .ZN(new_n745));
  OAI211_X1 g320(.A(new_n733), .B(new_n743), .C1(G1348), .C2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n678), .A2(G19), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT92), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(new_n606), .B2(G16), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(G1341), .Z(new_n750));
  INV_X1    g325(.A(KEYINPUT30), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n751), .A2(G28), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n718), .B1(new_n751), .B2(G28), .ZN(new_n753));
  AND2_X1   g328(.A1(KEYINPUT31), .A2(G11), .ZN(new_n754));
  NOR2_X1   g329(.A1(KEYINPUT31), .A2(G11), .ZN(new_n755));
  OAI22_X1  g330(.A1(new_n752), .A2(new_n753), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT24), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n718), .B1(new_n757), .B2(G34), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n757), .B2(G34), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G160), .B2(G29), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n756), .B1(new_n760), .B2(G2084), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G2084), .B2(new_n760), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n745), .A2(G1348), .ZN(new_n763));
  INV_X1    g338(.A(new_n617), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n764), .B2(new_n718), .ZN(new_n765));
  NOR4_X1   g340(.A1(new_n746), .A2(new_n750), .A3(new_n762), .A4(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n722), .A2(new_n723), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n718), .A2(G35), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G162), .B2(new_n718), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT29), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G2090), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n479), .A2(G141), .B1(G105), .B2(new_n462), .ZN(new_n772));
  NAND3_X1  g347(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT26), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n476), .B2(G129), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  MUX2_X1   g351(.A(G32), .B(new_n776), .S(G29), .Z(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT27), .ZN(new_n778));
  INV_X1    g353(.A(G1996), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n678), .A2(G5), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G171), .B2(new_n678), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G1961), .ZN(new_n783));
  NOR3_X1   g358(.A1(new_n771), .A2(new_n780), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n678), .A2(G21), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G168), .B2(new_n678), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G1966), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n678), .A2(G20), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT23), .Z(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G299), .B2(G16), .ZN(new_n790));
  INV_X1    g365(.A(G1956), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n787), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n766), .A2(new_n767), .A3(new_n784), .A4(new_n793), .ZN(new_n794));
  NOR3_X1   g369(.A1(new_n717), .A2(new_n724), .A3(new_n794), .ZN(G311));
  INV_X1    g370(.A(G311), .ZN(G150));
  AOI22_X1  g371(.A1(G93), .A2(new_n540), .B1(new_n522), .B2(G55), .ZN(new_n797));
  AOI22_X1  g372(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n798), .A2(new_n518), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n606), .B1(KEYINPUT98), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(KEYINPUT98), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n801), .B(new_n802), .Z(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT38), .Z(new_n804));
  NAND2_X1  g379(.A1(new_n597), .A2(G559), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n806), .A2(KEYINPUT39), .ZN(new_n807));
  INV_X1    g382(.A(G860), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n806), .A2(KEYINPUT39), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n807), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n800), .A2(new_n808), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT37), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n810), .A2(new_n812), .ZN(G145));
  XOR2_X1   g388(.A(new_n707), .B(KEYINPUT100), .Z(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(new_n620), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n476), .A2(G130), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n460), .A2(G118), .ZN(new_n817));
  OAI21_X1  g392(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n816), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(G142), .B2(new_n479), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n815), .B(new_n820), .Z(new_n821));
  NOR2_X1   g396(.A1(new_n487), .A2(KEYINPUT99), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT99), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(new_n484), .B2(new_n486), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n496), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n740), .B(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(new_n776), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(new_n731), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n821), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT101), .ZN(new_n830));
  OAI211_X1 g405(.A(new_n830), .B(KEYINPUT102), .C1(new_n821), .C2(new_n828), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n617), .B(G160), .Z(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(G162), .ZN(new_n833));
  AOI21_X1  g408(.A(G37), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(new_n833), .B2(new_n831), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g411(.A(new_n803), .B(new_n608), .Z(new_n837));
  INV_X1    g412(.A(G299), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n596), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n839), .B(KEYINPUT41), .Z(new_n842));
  OAI21_X1  g417(.A(new_n841), .B1(new_n837), .B2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(G288), .B(new_n580), .ZN(new_n844));
  XOR2_X1   g419(.A(G166), .B(new_n587), .Z(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT42), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n846), .B(KEYINPUT103), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n848), .B1(new_n849), .B2(new_n847), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n843), .B(new_n850), .Z(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(G868), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(G868), .B2(new_n800), .ZN(G331));
  XNOR2_X1  g428(.A(G331), .B(KEYINPUT104), .ZN(G295));
  INV_X1    g429(.A(KEYINPUT44), .ZN(new_n855));
  XNOR2_X1  g430(.A(G168), .B(G171), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n803), .A2(new_n856), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n857), .B(KEYINPUT105), .Z(new_n858));
  NOR2_X1   g433(.A1(new_n803), .A2(new_n856), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n859), .A2(new_n840), .ZN(new_n860));
  INV_X1    g435(.A(new_n859), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(new_n857), .ZN(new_n862));
  AOI22_X1  g437(.A1(new_n858), .A2(new_n860), .B1(new_n842), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(G37), .B1(new_n863), .B2(new_n849), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n858), .A2(new_n861), .ZN(new_n865));
  AOI22_X1  g440(.A1(new_n865), .A2(new_n842), .B1(new_n857), .B2(new_n860), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n864), .B1(new_n849), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n855), .B1(new_n867), .B2(KEYINPUT43), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n863), .A2(new_n849), .ZN(new_n869));
  AND2_X1   g444(.A1(new_n869), .A2(new_n864), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n868), .B1(new_n871), .B2(KEYINPUT43), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT106), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(KEYINPUT43), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n874), .B1(KEYINPUT43), .B2(new_n867), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(new_n855), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n873), .A2(new_n876), .ZN(G397));
  INV_X1    g452(.A(G1384), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n825), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n880), .A2(KEYINPUT45), .ZN(new_n881));
  NAND2_X1  g456(.A1(G160), .A2(G40), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n740), .B(G2067), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n885), .B1(new_n776), .B2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT46), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n889), .B1(new_n885), .B2(new_n779), .ZN(new_n890));
  NOR3_X1   g465(.A1(new_n884), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n888), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  XOR2_X1   g467(.A(new_n892), .B(KEYINPUT47), .Z(new_n893));
  XNOR2_X1  g468(.A(new_n776), .B(new_n779), .ZN(new_n894));
  OR2_X1    g469(.A1(new_n707), .A2(new_n710), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n707), .A2(new_n710), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n886), .A2(new_n894), .A3(new_n895), .A4(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n885), .A2(new_n897), .ZN(new_n898));
  XOR2_X1   g473(.A(new_n898), .B(KEYINPUT125), .Z(new_n899));
  NOR3_X1   g474(.A1(new_n884), .A2(G1986), .A3(G290), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(KEYINPUT48), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n886), .A2(new_n894), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n902), .A2(new_n895), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n903), .B1(new_n742), .B2(new_n740), .ZN(new_n904));
  OAI22_X1  g479(.A1(new_n899), .A2(new_n901), .B1(new_n884), .B2(new_n904), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n893), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT45), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n907), .A2(G1384), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n500), .A2(new_n508), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT113), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n500), .A2(new_n508), .A3(KEYINPUT113), .A4(new_n908), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n882), .B1(new_n879), .B2(new_n907), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT114), .ZN(new_n915));
  INV_X1    g490(.A(G1966), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT50), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n882), .B1(new_n880), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(G2084), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n500), .A2(new_n878), .A3(new_n508), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT50), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n919), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n917), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n915), .B1(new_n914), .B2(new_n916), .ZN(new_n925));
  OAI21_X1  g500(.A(KEYINPUT119), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(G8), .ZN(new_n927));
  NOR2_X1   g502(.A1(G168), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n914), .A2(new_n916), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(KEYINPUT114), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT119), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n930), .A2(new_n931), .A3(new_n923), .A4(new_n917), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n926), .A2(new_n928), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(G8), .B1(new_n924), .B2(new_n925), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT51), .ZN(new_n935));
  OAI211_X1 g510(.A(new_n934), .B(new_n935), .C1(new_n927), .C2(G168), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n936), .B(KEYINPUT122), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n926), .A2(G8), .A3(new_n932), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n928), .B1(new_n938), .B2(KEYINPUT120), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT120), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n926), .A2(new_n932), .A3(new_n940), .A4(G8), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n935), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT121), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n937), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AOI211_X1 g519(.A(KEYINPUT121), .B(new_n935), .C1(new_n939), .C2(new_n941), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n933), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(KEYINPUT62), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT62), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n948), .B(new_n933), .C1(new_n944), .C2(new_n945), .ZN(new_n949));
  NAND2_X1  g524(.A1(G303), .A2(G8), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n950), .B(KEYINPUT55), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n825), .A2(new_n908), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT107), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n953), .B(new_n954), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n955), .A2(new_n882), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n921), .A2(new_n907), .ZN(new_n957));
  AOI21_X1  g532(.A(G1971), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n919), .A2(new_n922), .ZN(new_n959));
  OAI22_X1  g534(.A1(new_n958), .A2(KEYINPUT108), .B1(new_n959), .B2(G2090), .ZN(new_n960));
  AND2_X1   g535(.A1(new_n958), .A2(KEYINPUT108), .ZN(new_n961));
  OAI211_X1 g536(.A(G8), .B(new_n952), .C1(new_n960), .C2(new_n961), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n879), .A2(new_n882), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n963), .A2(new_n927), .ZN(new_n964));
  INV_X1    g539(.A(G1981), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n574), .A2(new_n575), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(G651), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT110), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n965), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n969), .B(new_n580), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT111), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n970), .A2(new_n971), .A3(KEYINPUT49), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n971), .B1(new_n970), .B2(KEYINPUT49), .ZN(new_n973));
  OAI221_X1 g548(.A(new_n964), .B1(KEYINPUT49), .B2(new_n970), .C1(new_n972), .C2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(G288), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n975), .A2(G1976), .ZN(new_n976));
  AOI21_X1  g551(.A(KEYINPUT52), .B1(new_n976), .B2(new_n964), .ZN(new_n977));
  INV_X1    g552(.A(G1976), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n964), .B(KEYINPUT109), .C1(new_n978), .C2(G288), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n977), .B(new_n979), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n974), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n882), .B1(new_n879), .B2(KEYINPUT50), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n982), .B1(KEYINPUT50), .B2(new_n921), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n983), .A2(G2090), .ZN(new_n984));
  OAI21_X1  g559(.A(G8), .B1(new_n958), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(new_n951), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n962), .A2(new_n981), .A3(new_n986), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n956), .A2(new_n957), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT53), .B1(new_n988), .B2(new_n723), .ZN(new_n989));
  XNOR2_X1  g564(.A(KEYINPUT123), .B(G1961), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n989), .B1(new_n959), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n723), .A2(KEYINPUT53), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n991), .B1(new_n914), .B2(new_n992), .ZN(new_n993));
  AND3_X1   g568(.A1(new_n987), .A2(G171), .A3(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n947), .A2(new_n949), .A3(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n962), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n974), .A2(new_n978), .A3(new_n975), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n580), .A2(new_n965), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n998), .B(KEYINPUT112), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  AOI22_X1  g575(.A1(new_n996), .A2(new_n981), .B1(new_n1000), .B2(new_n964), .ZN(new_n1001));
  OR2_X1    g576(.A1(new_n934), .A2(G286), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT63), .B1(new_n987), .B2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(G8), .B1(new_n960), .B2(new_n961), .ZN(new_n1005));
  AND2_X1   g580(.A1(new_n1005), .A2(new_n951), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n962), .A2(KEYINPUT63), .A3(new_n981), .ZN(new_n1007));
  NOR3_X1   g582(.A1(new_n1006), .A2(new_n1007), .A3(new_n1002), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1001), .B1(new_n1004), .B2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g584(.A(G301), .B(KEYINPUT54), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n955), .A2(new_n992), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1010), .B1(new_n1011), .B2(new_n913), .ZN(new_n1012));
  AOI22_X1  g587(.A1(new_n993), .A2(new_n1010), .B1(new_n991), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n987), .ZN(new_n1014));
  XNOR2_X1  g589(.A(KEYINPUT56), .B(G2072), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n988), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT115), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n564), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT57), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n1020), .B(G299), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n983), .A2(new_n791), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1016), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1022), .B1(new_n1016), .B2(new_n1023), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G1348), .ZN(new_n1028));
  AOI22_X1  g603(.A1(new_n959), .A2(new_n1028), .B1(new_n742), .B2(new_n963), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n596), .A2(KEYINPUT60), .ZN(new_n1030));
  AOI22_X1  g605(.A1(new_n1027), .A2(KEYINPUT61), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1026), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n1024), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT61), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n1029), .B(new_n596), .ZN(new_n1035));
  AOI22_X1  g610(.A1(new_n1033), .A2(new_n1034), .B1(new_n1035), .B2(KEYINPUT60), .ZN(new_n1036));
  XNOR2_X1  g611(.A(KEYINPUT58), .B(G1341), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n963), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n988), .A2(new_n779), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1038), .B1(new_n1039), .B2(KEYINPUT116), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1040), .B1(KEYINPUT116), .B2(new_n1039), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT118), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n606), .B1(new_n1042), .B2(KEYINPUT59), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1042), .B1(KEYINPUT117), .B2(KEYINPUT59), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1045), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1041), .A2(new_n1047), .A3(new_n1043), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1031), .A2(new_n1036), .A3(new_n1046), .A4(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1029), .A2(new_n596), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1026), .B1(new_n1024), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1014), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1009), .B1(new_n1052), .B2(new_n946), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n995), .A2(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g629(.A(new_n587), .B(new_n700), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n885), .B1(new_n897), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(KEYINPUT124), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT124), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1056), .ZN(new_n1059));
  AOI211_X1 g634(.A(new_n1058), .B(new_n1059), .C1(new_n995), .C2(new_n1053), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n906), .B1(new_n1057), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(KEYINPUT126), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT126), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1063), .B(new_n906), .C1(new_n1057), .C2(new_n1060), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1062), .A2(new_n1064), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g640(.A1(new_n655), .A2(G319), .ZN(new_n1067));
  NOR3_X1   g641(.A1(G229), .A2(G401), .A3(new_n1067), .ZN(new_n1068));
  XOR2_X1   g642(.A(new_n1068), .B(KEYINPUT127), .Z(new_n1069));
  NAND3_X1  g643(.A1(new_n875), .A2(new_n835), .A3(new_n1069), .ZN(G225));
  INV_X1    g644(.A(G225), .ZN(G308));
endmodule


