

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X2 U548 ( .A(n703), .ZN(n706) );
  AND2_X1 U549 ( .A1(n740), .A2(n516), .ZN(n741) );
  AND2_X1 U550 ( .A1(n750), .A2(n749), .ZN(n751) );
  NOR2_X2 U551 ( .A1(n534), .A2(n533), .ZN(G160) );
  NOR2_X1 U552 ( .A1(n728), .A2(n678), .ZN(n515) );
  OR2_X1 U553 ( .A1(G1971), .A2(G303), .ZN(n516) );
  OR2_X1 U554 ( .A1(G1966), .A2(n758), .ZN(n517) );
  INV_X1 U555 ( .A(G8), .ZN(n678) );
  NAND2_X1 U556 ( .A1(n517), .A2(n515), .ZN(n679) );
  NAND2_X1 U557 ( .A1(n706), .A2(G8), .ZN(n758) );
  NAND2_X1 U558 ( .A1(G160), .A2(G40), .ZN(n783) );
  NOR2_X2 U559 ( .A1(G2105), .A2(n522), .ZN(n850) );
  NOR2_X1 U560 ( .A1(G651), .A2(n623), .ZN(n646) );
  BUF_X1 U561 ( .A(n675), .Z(G164) );
  INV_X1 U562 ( .A(G2104), .ZN(n522) );
  NAND2_X1 U563 ( .A1(G102), .A2(n850), .ZN(n521) );
  NOR2_X1 U564 ( .A1(G2104), .A2(G2105), .ZN(n518) );
  XOR2_X1 U565 ( .A(KEYINPUT66), .B(n518), .Z(n519) );
  XNOR2_X2 U566 ( .A(n519), .B(KEYINPUT17), .ZN(n851) );
  NAND2_X1 U567 ( .A1(n851), .A2(G138), .ZN(n520) );
  NAND2_X1 U568 ( .A1(n521), .A2(n520), .ZN(n527) );
  AND2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n854) );
  NAND2_X1 U570 ( .A1(G114), .A2(n854), .ZN(n525) );
  NAND2_X1 U571 ( .A1(n522), .A2(G2105), .ZN(n523) );
  XNOR2_X2 U572 ( .A(n523), .B(KEYINPUT65), .ZN(n855) );
  NAND2_X1 U573 ( .A1(G126), .A2(n855), .ZN(n524) );
  NAND2_X1 U574 ( .A1(n525), .A2(n524), .ZN(n526) );
  NOR2_X1 U575 ( .A1(n527), .A2(n526), .ZN(n675) );
  NAND2_X1 U576 ( .A1(n854), .A2(G113), .ZN(n530) );
  NAND2_X1 U577 ( .A1(G101), .A2(n850), .ZN(n528) );
  XOR2_X1 U578 ( .A(KEYINPUT23), .B(n528), .Z(n529) );
  NAND2_X1 U579 ( .A1(n530), .A2(n529), .ZN(n534) );
  NAND2_X1 U580 ( .A1(n855), .A2(G125), .ZN(n532) );
  NAND2_X1 U581 ( .A1(G137), .A2(n851), .ZN(n531) );
  NAND2_X1 U582 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U583 ( .A(KEYINPUT0), .B(G543), .Z(n623) );
  INV_X1 U584 ( .A(G651), .ZN(n539) );
  NOR2_X1 U585 ( .A1(n623), .A2(n539), .ZN(n642) );
  NAND2_X1 U586 ( .A1(n642), .A2(G77), .ZN(n535) );
  XOR2_X1 U587 ( .A(KEYINPUT69), .B(n535), .Z(n537) );
  NOR2_X1 U588 ( .A1(G651), .A2(G543), .ZN(n638) );
  NAND2_X1 U589 ( .A1(n638), .A2(G90), .ZN(n536) );
  NAND2_X1 U590 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U591 ( .A(n538), .B(KEYINPUT9), .ZN(n542) );
  NOR2_X1 U592 ( .A1(G543), .A2(n539), .ZN(n540) );
  XOR2_X1 U593 ( .A(KEYINPUT1), .B(n540), .Z(n637) );
  NAND2_X1 U594 ( .A1(G64), .A2(n637), .ZN(n541) );
  NAND2_X1 U595 ( .A1(n542), .A2(n541), .ZN(n545) );
  NAND2_X1 U596 ( .A1(n646), .A2(G52), .ZN(n543) );
  XOR2_X1 U597 ( .A(KEYINPUT68), .B(n543), .Z(n544) );
  NOR2_X1 U598 ( .A1(n545), .A2(n544), .ZN(G171) );
  AND2_X1 U599 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U600 ( .A(G69), .ZN(G235) );
  INV_X1 U601 ( .A(G108), .ZN(G238) );
  INV_X1 U602 ( .A(G82), .ZN(G220) );
  NAND2_X1 U603 ( .A1(G89), .A2(n638), .ZN(n546) );
  XOR2_X1 U604 ( .A(KEYINPUT4), .B(n546), .Z(n547) );
  XNOR2_X1 U605 ( .A(n547), .B(KEYINPUT77), .ZN(n549) );
  NAND2_X1 U606 ( .A1(G76), .A2(n642), .ZN(n548) );
  NAND2_X1 U607 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U608 ( .A(KEYINPUT5), .B(n550), .ZN(n556) );
  NAND2_X1 U609 ( .A1(G63), .A2(n637), .ZN(n552) );
  NAND2_X1 U610 ( .A1(G51), .A2(n646), .ZN(n551) );
  NAND2_X1 U611 ( .A1(n552), .A2(n551), .ZN(n554) );
  XOR2_X1 U612 ( .A(KEYINPUT6), .B(KEYINPUT78), .Z(n553) );
  XNOR2_X1 U613 ( .A(n554), .B(n553), .ZN(n555) );
  NAND2_X1 U614 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U615 ( .A(KEYINPUT7), .B(n557), .ZN(G168) );
  XOR2_X1 U616 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U617 ( .A1(G7), .A2(G661), .ZN(n558) );
  XNOR2_X1 U618 ( .A(n558), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U619 ( .A(G223), .B(KEYINPUT72), .Z(n824) );
  NAND2_X1 U620 ( .A1(n824), .A2(G567), .ZN(n559) );
  XOR2_X1 U621 ( .A(KEYINPUT11), .B(n559), .Z(G234) );
  XOR2_X1 U622 ( .A(KEYINPUT12), .B(KEYINPUT74), .Z(n561) );
  NAND2_X1 U623 ( .A1(G81), .A2(n638), .ZN(n560) );
  XNOR2_X1 U624 ( .A(n561), .B(n560), .ZN(n564) );
  NAND2_X1 U625 ( .A1(n642), .A2(G68), .ZN(n562) );
  XNOR2_X1 U626 ( .A(KEYINPUT75), .B(n562), .ZN(n563) );
  NOR2_X1 U627 ( .A1(n564), .A2(n563), .ZN(n566) );
  XNOR2_X1 U628 ( .A(KEYINPUT76), .B(KEYINPUT13), .ZN(n565) );
  XNOR2_X1 U629 ( .A(n566), .B(n565), .ZN(n570) );
  NAND2_X1 U630 ( .A1(G56), .A2(n637), .ZN(n567) );
  XNOR2_X1 U631 ( .A(n567), .B(KEYINPUT14), .ZN(n568) );
  XNOR2_X1 U632 ( .A(n568), .B(KEYINPUT73), .ZN(n569) );
  NOR2_X1 U633 ( .A1(n570), .A2(n569), .ZN(n572) );
  NAND2_X1 U634 ( .A1(n646), .A2(G43), .ZN(n571) );
  NAND2_X1 U635 ( .A1(n572), .A2(n571), .ZN(n986) );
  INV_X1 U636 ( .A(G860), .ZN(n613) );
  OR2_X1 U637 ( .A1(n986), .A2(n613), .ZN(G153) );
  INV_X1 U638 ( .A(G171), .ZN(G301) );
  NAND2_X1 U639 ( .A1(G868), .A2(G301), .ZN(n581) );
  NAND2_X1 U640 ( .A1(G92), .A2(n638), .ZN(n574) );
  NAND2_X1 U641 ( .A1(G79), .A2(n642), .ZN(n573) );
  NAND2_X1 U642 ( .A1(n574), .A2(n573), .ZN(n578) );
  NAND2_X1 U643 ( .A1(G66), .A2(n637), .ZN(n576) );
  NAND2_X1 U644 ( .A1(G54), .A2(n646), .ZN(n575) );
  NAND2_X1 U645 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U646 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U647 ( .A(KEYINPUT15), .B(n579), .Z(n987) );
  OR2_X1 U648 ( .A1(n987), .A2(G868), .ZN(n580) );
  NAND2_X1 U649 ( .A1(n581), .A2(n580), .ZN(G284) );
  NAND2_X1 U650 ( .A1(G65), .A2(n637), .ZN(n583) );
  NAND2_X1 U651 ( .A1(G53), .A2(n646), .ZN(n582) );
  NAND2_X1 U652 ( .A1(n583), .A2(n582), .ZN(n587) );
  NAND2_X1 U653 ( .A1(G91), .A2(n638), .ZN(n585) );
  NAND2_X1 U654 ( .A1(G78), .A2(n642), .ZN(n584) );
  NAND2_X1 U655 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U656 ( .A1(n587), .A2(n586), .ZN(n990) );
  INV_X1 U657 ( .A(n990), .ZN(G299) );
  INV_X1 U658 ( .A(G868), .ZN(n658) );
  NOR2_X1 U659 ( .A1(G286), .A2(n658), .ZN(n589) );
  NOR2_X1 U660 ( .A1(G868), .A2(G299), .ZN(n588) );
  NOR2_X1 U661 ( .A1(n589), .A2(n588), .ZN(G297) );
  NAND2_X1 U662 ( .A1(n613), .A2(G559), .ZN(n590) );
  NAND2_X1 U663 ( .A1(n590), .A2(n987), .ZN(n591) );
  XNOR2_X1 U664 ( .A(n591), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U665 ( .A1(G868), .A2(n986), .ZN(n594) );
  NAND2_X1 U666 ( .A1(G868), .A2(n987), .ZN(n592) );
  NOR2_X1 U667 ( .A1(G559), .A2(n592), .ZN(n593) );
  NOR2_X1 U668 ( .A1(n594), .A2(n593), .ZN(G282) );
  NAND2_X1 U669 ( .A1(G99), .A2(n850), .ZN(n596) );
  NAND2_X1 U670 ( .A1(G111), .A2(n854), .ZN(n595) );
  NAND2_X1 U671 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U672 ( .A(KEYINPUT80), .B(n597), .ZN(n603) );
  NAND2_X1 U673 ( .A1(G123), .A2(n855), .ZN(n598) );
  XOR2_X1 U674 ( .A(KEYINPUT18), .B(n598), .Z(n599) );
  XNOR2_X1 U675 ( .A(n599), .B(KEYINPUT79), .ZN(n601) );
  NAND2_X1 U676 ( .A1(G135), .A2(n851), .ZN(n600) );
  NAND2_X1 U677 ( .A1(n601), .A2(n600), .ZN(n602) );
  NOR2_X1 U678 ( .A1(n603), .A2(n602), .ZN(n959) );
  XNOR2_X1 U679 ( .A(n959), .B(G2096), .ZN(n605) );
  INV_X1 U680 ( .A(G2100), .ZN(n604) );
  NAND2_X1 U681 ( .A1(n605), .A2(n604), .ZN(G156) );
  NAND2_X1 U682 ( .A1(G67), .A2(n637), .ZN(n607) );
  NAND2_X1 U683 ( .A1(G55), .A2(n646), .ZN(n606) );
  NAND2_X1 U684 ( .A1(n607), .A2(n606), .ZN(n611) );
  NAND2_X1 U685 ( .A1(G93), .A2(n638), .ZN(n609) );
  NAND2_X1 U686 ( .A1(G80), .A2(n642), .ZN(n608) );
  NAND2_X1 U687 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U688 ( .A1(n611), .A2(n610), .ZN(n657) );
  NAND2_X1 U689 ( .A1(G559), .A2(n987), .ZN(n612) );
  XOR2_X1 U690 ( .A(n986), .B(n612), .Z(n655) );
  NAND2_X1 U691 ( .A1(n613), .A2(n655), .ZN(n614) );
  XNOR2_X1 U692 ( .A(n614), .B(KEYINPUT81), .ZN(n615) );
  XNOR2_X1 U693 ( .A(n657), .B(n615), .ZN(G145) );
  NAND2_X1 U694 ( .A1(G60), .A2(n637), .ZN(n617) );
  NAND2_X1 U695 ( .A1(G47), .A2(n646), .ZN(n616) );
  NAND2_X1 U696 ( .A1(n617), .A2(n616), .ZN(n621) );
  NAND2_X1 U697 ( .A1(G85), .A2(n638), .ZN(n619) );
  NAND2_X1 U698 ( .A1(G72), .A2(n642), .ZN(n618) );
  NAND2_X1 U699 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U700 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U701 ( .A(n622), .B(KEYINPUT67), .ZN(G290) );
  NAND2_X1 U702 ( .A1(G74), .A2(G651), .ZN(n628) );
  NAND2_X1 U703 ( .A1(G49), .A2(n646), .ZN(n625) );
  NAND2_X1 U704 ( .A1(G87), .A2(n623), .ZN(n624) );
  NAND2_X1 U705 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U706 ( .A1(n637), .A2(n626), .ZN(n627) );
  NAND2_X1 U707 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U708 ( .A(n629), .B(KEYINPUT82), .ZN(G288) );
  NAND2_X1 U709 ( .A1(G62), .A2(n637), .ZN(n631) );
  NAND2_X1 U710 ( .A1(G50), .A2(n646), .ZN(n630) );
  NAND2_X1 U711 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U712 ( .A(KEYINPUT84), .B(n632), .ZN(n636) );
  NAND2_X1 U713 ( .A1(G88), .A2(n638), .ZN(n634) );
  NAND2_X1 U714 ( .A1(G75), .A2(n642), .ZN(n633) );
  NAND2_X1 U715 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U716 ( .A1(n636), .A2(n635), .ZN(G166) );
  INV_X1 U717 ( .A(G166), .ZN(G303) );
  NAND2_X1 U718 ( .A1(n637), .A2(G61), .ZN(n640) );
  NAND2_X1 U719 ( .A1(n638), .A2(G86), .ZN(n639) );
  NAND2_X1 U720 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U721 ( .A(KEYINPUT83), .B(n641), .Z(n645) );
  NAND2_X1 U722 ( .A1(G73), .A2(n642), .ZN(n643) );
  XOR2_X1 U723 ( .A(KEYINPUT2), .B(n643), .Z(n644) );
  NOR2_X1 U724 ( .A1(n645), .A2(n644), .ZN(n648) );
  NAND2_X1 U725 ( .A1(n646), .A2(G48), .ZN(n647) );
  NAND2_X1 U726 ( .A1(n648), .A2(n647), .ZN(G305) );
  XOR2_X1 U727 ( .A(KEYINPUT19), .B(KEYINPUT85), .Z(n649) );
  XNOR2_X1 U728 ( .A(G290), .B(n649), .ZN(n650) );
  XOR2_X1 U729 ( .A(n650), .B(n657), .Z(n652) );
  XNOR2_X1 U730 ( .A(G288), .B(n990), .ZN(n651) );
  XNOR2_X1 U731 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U732 ( .A(n653), .B(G303), .ZN(n654) );
  XNOR2_X1 U733 ( .A(n654), .B(G305), .ZN(n876) );
  XNOR2_X1 U734 ( .A(n655), .B(n876), .ZN(n656) );
  NAND2_X1 U735 ( .A1(n656), .A2(G868), .ZN(n660) );
  NAND2_X1 U736 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U737 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U738 ( .A(KEYINPUT86), .B(n661), .Z(G295) );
  NAND2_X1 U739 ( .A1(G2084), .A2(G2078), .ZN(n662) );
  XOR2_X1 U740 ( .A(KEYINPUT20), .B(n662), .Z(n663) );
  NAND2_X1 U741 ( .A1(G2090), .A2(n663), .ZN(n664) );
  XNOR2_X1 U742 ( .A(KEYINPUT21), .B(n664), .ZN(n665) );
  NAND2_X1 U743 ( .A1(n665), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U744 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U745 ( .A(KEYINPUT71), .B(G132), .ZN(G219) );
  XOR2_X1 U746 ( .A(KEYINPUT70), .B(G57), .Z(G237) );
  NOR2_X1 U747 ( .A1(G220), .A2(G219), .ZN(n666) );
  XOR2_X1 U748 ( .A(KEYINPUT22), .B(n666), .Z(n667) );
  NOR2_X1 U749 ( .A1(G218), .A2(n667), .ZN(n668) );
  NAND2_X1 U750 ( .A1(G96), .A2(n668), .ZN(n831) );
  NAND2_X1 U751 ( .A1(n831), .A2(G2106), .ZN(n673) );
  NOR2_X1 U752 ( .A1(G237), .A2(G238), .ZN(n669) );
  NAND2_X1 U753 ( .A1(G120), .A2(n669), .ZN(n670) );
  NOR2_X1 U754 ( .A1(n670), .A2(G235), .ZN(n671) );
  XNOR2_X1 U755 ( .A(n671), .B(KEYINPUT87), .ZN(n832) );
  NAND2_X1 U756 ( .A1(n832), .A2(G567), .ZN(n672) );
  NAND2_X1 U757 ( .A1(n673), .A2(n672), .ZN(n899) );
  NAND2_X1 U758 ( .A1(G483), .A2(G661), .ZN(n674) );
  NOR2_X1 U759 ( .A1(n899), .A2(n674), .ZN(n828) );
  NAND2_X1 U760 ( .A1(n828), .A2(G36), .ZN(G176) );
  NOR2_X2 U761 ( .A1(n675), .A2(G1384), .ZN(n784) );
  INV_X1 U762 ( .A(n784), .ZN(n676) );
  NOR2_X2 U763 ( .A1(n676), .A2(n783), .ZN(n677) );
  XNOR2_X2 U764 ( .A(n677), .B(KEYINPUT64), .ZN(n703) );
  INV_X1 U765 ( .A(n758), .ZN(n745) );
  NOR2_X1 U766 ( .A1(n706), .A2(G2084), .ZN(n728) );
  XNOR2_X1 U767 ( .A(KEYINPUT30), .B(n679), .ZN(n680) );
  NOR2_X1 U768 ( .A1(G168), .A2(n680), .ZN(n684) );
  XNOR2_X1 U769 ( .A(KEYINPUT25), .B(G2078), .ZN(n909) );
  NAND2_X1 U770 ( .A1(n703), .A2(n909), .ZN(n682) );
  INV_X1 U771 ( .A(G1961), .ZN(n996) );
  NAND2_X1 U772 ( .A1(n706), .A2(n996), .ZN(n681) );
  NAND2_X1 U773 ( .A1(n682), .A2(n681), .ZN(n691) );
  NOR2_X1 U774 ( .A1(G171), .A2(n691), .ZN(n683) );
  NOR2_X1 U775 ( .A1(n684), .A2(n683), .ZN(n686) );
  INV_X1 U776 ( .A(KEYINPUT31), .ZN(n685) );
  XNOR2_X1 U777 ( .A(n686), .B(n685), .ZN(n725) );
  NOR2_X1 U778 ( .A1(n706), .A2(G2090), .ZN(n688) );
  NOR2_X1 U779 ( .A1(G1971), .A2(n758), .ZN(n687) );
  NOR2_X1 U780 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U781 ( .A1(n689), .A2(G303), .ZN(n690) );
  OR2_X1 U782 ( .A1(n678), .A2(n690), .ZN(n719) );
  AND2_X1 U783 ( .A1(n725), .A2(n719), .ZN(n718) );
  NAND2_X1 U784 ( .A1(n691), .A2(G171), .ZN(n717) );
  NAND2_X1 U785 ( .A1(n703), .A2(G1996), .ZN(n692) );
  XNOR2_X1 U786 ( .A(n692), .B(KEYINPUT26), .ZN(n694) );
  NAND2_X1 U787 ( .A1(n706), .A2(G1341), .ZN(n693) );
  NAND2_X1 U788 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U789 ( .A1(n986), .A2(n695), .ZN(n700) );
  NAND2_X1 U790 ( .A1(n700), .A2(n987), .ZN(n699) );
  NAND2_X1 U791 ( .A1(G2067), .A2(n703), .ZN(n697) );
  NAND2_X1 U792 ( .A1(n706), .A2(G1348), .ZN(n696) );
  NAND2_X1 U793 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U794 ( .A1(n699), .A2(n698), .ZN(n702) );
  OR2_X1 U795 ( .A1(n700), .A2(n987), .ZN(n701) );
  NAND2_X1 U796 ( .A1(n702), .A2(n701), .ZN(n710) );
  NAND2_X1 U797 ( .A1(n703), .A2(G2072), .ZN(n705) );
  XNOR2_X1 U798 ( .A(KEYINPUT92), .B(KEYINPUT27), .ZN(n704) );
  XNOR2_X1 U799 ( .A(n705), .B(n704), .ZN(n708) );
  AND2_X1 U800 ( .A1(n706), .A2(G1956), .ZN(n707) );
  NOR2_X1 U801 ( .A1(n708), .A2(n707), .ZN(n711) );
  NAND2_X1 U802 ( .A1(n711), .A2(n990), .ZN(n709) );
  NAND2_X1 U803 ( .A1(n710), .A2(n709), .ZN(n714) );
  NOR2_X1 U804 ( .A1(n711), .A2(n990), .ZN(n712) );
  XOR2_X1 U805 ( .A(n712), .B(KEYINPUT28), .Z(n713) );
  NAND2_X1 U806 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U807 ( .A(n715), .B(KEYINPUT29), .Z(n716) );
  NAND2_X1 U808 ( .A1(n717), .A2(n716), .ZN(n726) );
  NAND2_X1 U809 ( .A1(n718), .A2(n726), .ZN(n723) );
  INV_X1 U810 ( .A(n719), .ZN(n721) );
  AND2_X1 U811 ( .A1(G286), .A2(G8), .ZN(n720) );
  OR2_X1 U812 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U813 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U814 ( .A(KEYINPUT32), .B(n724), .Z(n733) );
  NAND2_X1 U815 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U816 ( .A(n727), .B(KEYINPUT93), .ZN(n731) );
  NAND2_X1 U817 ( .A1(G8), .A2(n728), .ZN(n729) );
  NAND2_X1 U818 ( .A1(n729), .A2(n517), .ZN(n730) );
  NOR2_X1 U819 ( .A1(n731), .A2(n730), .ZN(n732) );
  NOR2_X1 U820 ( .A1(n733), .A2(n732), .ZN(n737) );
  NAND2_X1 U821 ( .A1(G166), .A2(G8), .ZN(n734) );
  NOR2_X1 U822 ( .A1(G2090), .A2(n734), .ZN(n735) );
  NOR2_X1 U823 ( .A1(n737), .A2(n735), .ZN(n736) );
  NOR2_X1 U824 ( .A1(n745), .A2(n736), .ZN(n754) );
  INV_X1 U825 ( .A(n737), .ZN(n742) );
  NOR2_X1 U826 ( .A1(G288), .A2(G1976), .ZN(n738) );
  XOR2_X1 U827 ( .A(n738), .B(KEYINPUT94), .Z(n995) );
  OR2_X1 U828 ( .A1(n995), .A2(n758), .ZN(n739) );
  NAND2_X1 U829 ( .A1(n739), .A2(KEYINPUT33), .ZN(n743) );
  AND2_X1 U830 ( .A1(n995), .A2(n743), .ZN(n740) );
  NAND2_X1 U831 ( .A1(n742), .A2(n741), .ZN(n750) );
  INV_X1 U832 ( .A(n743), .ZN(n748) );
  INV_X1 U833 ( .A(KEYINPUT33), .ZN(n744) );
  NAND2_X1 U834 ( .A1(G1976), .A2(G288), .ZN(n991) );
  AND2_X1 U835 ( .A1(n744), .A2(n991), .ZN(n746) );
  AND2_X1 U836 ( .A1(n746), .A2(n745), .ZN(n747) );
  OR2_X1 U837 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U838 ( .A(n751), .B(KEYINPUT95), .ZN(n752) );
  XNOR2_X1 U839 ( .A(G1981), .B(G305), .ZN(n1007) );
  NOR2_X1 U840 ( .A1(n752), .A2(n1007), .ZN(n753) );
  NOR2_X1 U841 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U842 ( .A(KEYINPUT96), .B(n755), .ZN(n788) );
  NOR2_X1 U843 ( .A1(G1981), .A2(G305), .ZN(n756) );
  XOR2_X1 U844 ( .A(n756), .B(KEYINPUT24), .Z(n757) );
  NOR2_X1 U845 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U846 ( .A(KEYINPUT91), .B(n759), .ZN(n786) );
  INV_X1 U847 ( .A(G1996), .ZN(n776) );
  NAND2_X1 U848 ( .A1(n854), .A2(G117), .ZN(n761) );
  NAND2_X1 U849 ( .A1(G141), .A2(n851), .ZN(n760) );
  NAND2_X1 U850 ( .A1(n761), .A2(n760), .ZN(n767) );
  NAND2_X1 U851 ( .A1(G129), .A2(n855), .ZN(n762) );
  XNOR2_X1 U852 ( .A(n762), .B(KEYINPUT90), .ZN(n765) );
  NAND2_X1 U853 ( .A1(G105), .A2(n850), .ZN(n763) );
  XNOR2_X1 U854 ( .A(n763), .B(KEYINPUT38), .ZN(n764) );
  NAND2_X1 U855 ( .A1(n765), .A2(n764), .ZN(n766) );
  NOR2_X1 U856 ( .A1(n767), .A2(n766), .ZN(n865) );
  AND2_X1 U857 ( .A1(n776), .A2(n865), .ZN(n768) );
  XOR2_X1 U858 ( .A(KEYINPUT97), .B(n768), .Z(n971) );
  NAND2_X1 U859 ( .A1(G95), .A2(n850), .ZN(n770) );
  NAND2_X1 U860 ( .A1(G107), .A2(n854), .ZN(n769) );
  NAND2_X1 U861 ( .A1(n770), .A2(n769), .ZN(n774) );
  NAND2_X1 U862 ( .A1(n855), .A2(G119), .ZN(n772) );
  NAND2_X1 U863 ( .A1(G131), .A2(n851), .ZN(n771) );
  NAND2_X1 U864 ( .A1(n772), .A2(n771), .ZN(n773) );
  OR2_X1 U865 ( .A1(n774), .A2(n773), .ZN(n862) );
  NAND2_X1 U866 ( .A1(G1991), .A2(n862), .ZN(n775) );
  XNOR2_X1 U867 ( .A(n775), .B(KEYINPUT89), .ZN(n778) );
  NOR2_X1 U868 ( .A1(n776), .A2(n865), .ZN(n777) );
  NOR2_X1 U869 ( .A1(n778), .A2(n777), .ZN(n800) );
  INV_X1 U870 ( .A(n800), .ZN(n965) );
  NOR2_X1 U871 ( .A1(G1986), .A2(G290), .ZN(n779) );
  NOR2_X1 U872 ( .A1(G1991), .A2(n862), .ZN(n960) );
  NOR2_X1 U873 ( .A1(n779), .A2(n960), .ZN(n780) );
  NOR2_X1 U874 ( .A1(n965), .A2(n780), .ZN(n781) );
  NOR2_X1 U875 ( .A1(n971), .A2(n781), .ZN(n782) );
  XNOR2_X1 U876 ( .A(KEYINPUT39), .B(n782), .ZN(n785) );
  NOR2_X1 U877 ( .A1(n784), .A2(n783), .ZN(n809) );
  NAND2_X1 U878 ( .A1(n785), .A2(n809), .ZN(n799) );
  AND2_X1 U879 ( .A1(n786), .A2(n799), .ZN(n787) );
  NAND2_X1 U880 ( .A1(n788), .A2(n787), .ZN(n807) );
  NAND2_X1 U881 ( .A1(G116), .A2(n854), .ZN(n790) );
  NAND2_X1 U882 ( .A1(G128), .A2(n855), .ZN(n789) );
  NAND2_X1 U883 ( .A1(n790), .A2(n789), .ZN(n792) );
  XOR2_X1 U884 ( .A(KEYINPUT88), .B(KEYINPUT35), .Z(n791) );
  XNOR2_X1 U885 ( .A(n792), .B(n791), .ZN(n797) );
  NAND2_X1 U886 ( .A1(G104), .A2(n850), .ZN(n794) );
  NAND2_X1 U887 ( .A1(G140), .A2(n851), .ZN(n793) );
  NAND2_X1 U888 ( .A1(n794), .A2(n793), .ZN(n795) );
  XNOR2_X1 U889 ( .A(KEYINPUT34), .B(n795), .ZN(n796) );
  NOR2_X1 U890 ( .A1(n797), .A2(n796), .ZN(n798) );
  XOR2_X1 U891 ( .A(KEYINPUT36), .B(n798), .Z(n871) );
  XOR2_X1 U892 ( .A(G2067), .B(KEYINPUT37), .Z(n808) );
  AND2_X1 U893 ( .A1(n871), .A2(n808), .ZN(n958) );
  NAND2_X1 U894 ( .A1(n958), .A2(n809), .ZN(n805) );
  INV_X1 U895 ( .A(n799), .ZN(n803) );
  XOR2_X1 U896 ( .A(G1986), .B(G290), .Z(n988) );
  NAND2_X1 U897 ( .A1(n988), .A2(n800), .ZN(n801) );
  NAND2_X1 U898 ( .A1(n801), .A2(n809), .ZN(n802) );
  OR2_X1 U899 ( .A1(n803), .A2(n802), .ZN(n804) );
  AND2_X1 U900 ( .A1(n805), .A2(n804), .ZN(n806) );
  NAND2_X1 U901 ( .A1(n807), .A2(n806), .ZN(n811) );
  NOR2_X1 U902 ( .A1(n871), .A2(n808), .ZN(n968) );
  NAND2_X1 U903 ( .A1(n968), .A2(n809), .ZN(n810) );
  NAND2_X1 U904 ( .A1(n811), .A2(n810), .ZN(n812) );
  XNOR2_X1 U905 ( .A(n812), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U906 ( .A(G2427), .B(G2451), .ZN(n822) );
  XOR2_X1 U907 ( .A(G2430), .B(G2443), .Z(n814) );
  XNOR2_X1 U908 ( .A(G2435), .B(KEYINPUT99), .ZN(n813) );
  XNOR2_X1 U909 ( .A(n814), .B(n813), .ZN(n818) );
  XOR2_X1 U910 ( .A(G2438), .B(G2454), .Z(n816) );
  XNOR2_X1 U911 ( .A(G1348), .B(G1341), .ZN(n815) );
  XNOR2_X1 U912 ( .A(n816), .B(n815), .ZN(n817) );
  XOR2_X1 U913 ( .A(n818), .B(n817), .Z(n820) );
  XNOR2_X1 U914 ( .A(KEYINPUT98), .B(G2446), .ZN(n819) );
  XNOR2_X1 U915 ( .A(n820), .B(n819), .ZN(n821) );
  XNOR2_X1 U916 ( .A(n822), .B(n821), .ZN(n823) );
  NAND2_X1 U917 ( .A1(n823), .A2(G14), .ZN(n902) );
  XOR2_X1 U918 ( .A(KEYINPUT100), .B(n902), .Z(G401) );
  NAND2_X1 U919 ( .A1(G2106), .A2(n824), .ZN(G217) );
  NAND2_X1 U920 ( .A1(G15), .A2(G2), .ZN(n825) );
  XNOR2_X1 U921 ( .A(KEYINPUT101), .B(n825), .ZN(n826) );
  NAND2_X1 U922 ( .A1(n826), .A2(G661), .ZN(G259) );
  NAND2_X1 U923 ( .A1(G3), .A2(G1), .ZN(n827) );
  XNOR2_X1 U924 ( .A(KEYINPUT102), .B(n827), .ZN(n829) );
  NAND2_X1 U925 ( .A1(n829), .A2(n828), .ZN(n830) );
  XOR2_X1 U926 ( .A(KEYINPUT103), .B(n830), .Z(G188) );
  INV_X1 U928 ( .A(G96), .ZN(G221) );
  NOR2_X1 U929 ( .A1(n832), .A2(n831), .ZN(G325) );
  INV_X1 U930 ( .A(G325), .ZN(G261) );
  NAND2_X1 U931 ( .A1(G100), .A2(n850), .ZN(n834) );
  NAND2_X1 U932 ( .A1(G112), .A2(n854), .ZN(n833) );
  NAND2_X1 U933 ( .A1(n834), .A2(n833), .ZN(n839) );
  NAND2_X1 U934 ( .A1(G124), .A2(n855), .ZN(n835) );
  XNOR2_X1 U935 ( .A(n835), .B(KEYINPUT44), .ZN(n837) );
  NAND2_X1 U936 ( .A1(G136), .A2(n851), .ZN(n836) );
  NAND2_X1 U937 ( .A1(n837), .A2(n836), .ZN(n838) );
  NOR2_X1 U938 ( .A1(n839), .A2(n838), .ZN(G162) );
  XNOR2_X1 U939 ( .A(n959), .B(KEYINPUT48), .ZN(n840) );
  XNOR2_X1 U940 ( .A(n840), .B(KEYINPUT46), .ZN(n841) );
  XNOR2_X1 U941 ( .A(G164), .B(n841), .ZN(n869) );
  NAND2_X1 U942 ( .A1(G106), .A2(n850), .ZN(n843) );
  NAND2_X1 U943 ( .A1(G142), .A2(n851), .ZN(n842) );
  NAND2_X1 U944 ( .A1(n843), .A2(n842), .ZN(n844) );
  XNOR2_X1 U945 ( .A(n844), .B(KEYINPUT45), .ZN(n846) );
  NAND2_X1 U946 ( .A1(G130), .A2(n855), .ZN(n845) );
  NAND2_X1 U947 ( .A1(n846), .A2(n845), .ZN(n849) );
  NAND2_X1 U948 ( .A1(n854), .A2(G118), .ZN(n847) );
  XOR2_X1 U949 ( .A(KEYINPUT106), .B(n847), .Z(n848) );
  NOR2_X1 U950 ( .A1(n849), .A2(n848), .ZN(n864) );
  NAND2_X1 U951 ( .A1(G103), .A2(n850), .ZN(n853) );
  NAND2_X1 U952 ( .A1(G139), .A2(n851), .ZN(n852) );
  NAND2_X1 U953 ( .A1(n853), .A2(n852), .ZN(n860) );
  NAND2_X1 U954 ( .A1(G115), .A2(n854), .ZN(n857) );
  NAND2_X1 U955 ( .A1(G127), .A2(n855), .ZN(n856) );
  NAND2_X1 U956 ( .A1(n857), .A2(n856), .ZN(n858) );
  XOR2_X1 U957 ( .A(KEYINPUT47), .B(n858), .Z(n859) );
  NOR2_X1 U958 ( .A1(n860), .A2(n859), .ZN(n975) );
  XOR2_X1 U959 ( .A(G162), .B(n975), .Z(n861) );
  XNOR2_X1 U960 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U961 ( .A(n864), .B(n863), .Z(n867) );
  XNOR2_X1 U962 ( .A(G160), .B(n865), .ZN(n866) );
  XNOR2_X1 U963 ( .A(n867), .B(n866), .ZN(n868) );
  XNOR2_X1 U964 ( .A(n869), .B(n868), .ZN(n870) );
  XNOR2_X1 U965 ( .A(n871), .B(n870), .ZN(n872) );
  NOR2_X1 U966 ( .A1(G37), .A2(n872), .ZN(n873) );
  XOR2_X1 U967 ( .A(KEYINPUT107), .B(n873), .Z(G395) );
  XNOR2_X1 U968 ( .A(n986), .B(KEYINPUT108), .ZN(n875) );
  XNOR2_X1 U969 ( .A(G171), .B(n987), .ZN(n874) );
  XNOR2_X1 U970 ( .A(n875), .B(n874), .ZN(n878) );
  XOR2_X1 U971 ( .A(G286), .B(n876), .Z(n877) );
  XNOR2_X1 U972 ( .A(n878), .B(n877), .ZN(n879) );
  NOR2_X1 U973 ( .A1(G37), .A2(n879), .ZN(G397) );
  XOR2_X1 U974 ( .A(KEYINPUT41), .B(G1991), .Z(n881) );
  XNOR2_X1 U975 ( .A(G1981), .B(G1996), .ZN(n880) );
  XNOR2_X1 U976 ( .A(n881), .B(n880), .ZN(n882) );
  XOR2_X1 U977 ( .A(n882), .B(KEYINPUT105), .Z(n884) );
  XNOR2_X1 U978 ( .A(G1976), .B(G1971), .ZN(n883) );
  XNOR2_X1 U979 ( .A(n884), .B(n883), .ZN(n888) );
  XOR2_X1 U980 ( .A(G1986), .B(G1956), .Z(n886) );
  XNOR2_X1 U981 ( .A(G1966), .B(G1961), .ZN(n885) );
  XNOR2_X1 U982 ( .A(n886), .B(n885), .ZN(n887) );
  XOR2_X1 U983 ( .A(n888), .B(n887), .Z(n890) );
  XNOR2_X1 U984 ( .A(KEYINPUT104), .B(G2474), .ZN(n889) );
  XNOR2_X1 U985 ( .A(n890), .B(n889), .ZN(G229) );
  XOR2_X1 U986 ( .A(G2100), .B(G2096), .Z(n892) );
  XNOR2_X1 U987 ( .A(KEYINPUT42), .B(G2678), .ZN(n891) );
  XNOR2_X1 U988 ( .A(n892), .B(n891), .ZN(n896) );
  XOR2_X1 U989 ( .A(KEYINPUT43), .B(G2090), .Z(n894) );
  XNOR2_X1 U990 ( .A(G2067), .B(G2072), .ZN(n893) );
  XNOR2_X1 U991 ( .A(n894), .B(n893), .ZN(n895) );
  XOR2_X1 U992 ( .A(n896), .B(n895), .Z(n898) );
  XNOR2_X1 U993 ( .A(G2084), .B(G2078), .ZN(n897) );
  XNOR2_X1 U994 ( .A(n898), .B(n897), .ZN(G227) );
  INV_X1 U995 ( .A(n899), .ZN(G319) );
  NOR2_X1 U996 ( .A1(G395), .A2(G397), .ZN(n900) );
  XNOR2_X1 U997 ( .A(n900), .B(KEYINPUT110), .ZN(n901) );
  NAND2_X1 U998 ( .A1(n902), .A2(n901), .ZN(n906) );
  NOR2_X1 U999 ( .A1(G229), .A2(G227), .ZN(n903) );
  XOR2_X1 U1000 ( .A(KEYINPUT109), .B(n903), .Z(n904) );
  XNOR2_X1 U1001 ( .A(n904), .B(KEYINPUT49), .ZN(n905) );
  NOR2_X1 U1002 ( .A1(n906), .A2(n905), .ZN(n907) );
  NAND2_X1 U1003 ( .A1(n907), .A2(G319), .ZN(n908) );
  XOR2_X1 U1004 ( .A(KEYINPUT111), .B(n908), .Z(G225) );
  XOR2_X1 U1005 ( .A(KEYINPUT112), .B(G225), .Z(G308) );
  INV_X1 U1006 ( .A(G120), .ZN(G236) );
  XNOR2_X1 U1007 ( .A(G1991), .B(G25), .ZN(n919) );
  XOR2_X1 U1008 ( .A(G2072), .B(G33), .Z(n914) );
  XOR2_X1 U1009 ( .A(n909), .B(G27), .Z(n911) );
  XNOR2_X1 U1010 ( .A(G32), .B(G1996), .ZN(n910) );
  NOR2_X1 U1011 ( .A1(n911), .A2(n910), .ZN(n912) );
  XNOR2_X1 U1012 ( .A(KEYINPUT118), .B(n912), .ZN(n913) );
  NAND2_X1 U1013 ( .A1(n914), .A2(n913), .ZN(n916) );
  XNOR2_X1 U1014 ( .A(G26), .B(G2067), .ZN(n915) );
  NOR2_X1 U1015 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1016 ( .A(KEYINPUT119), .B(n917), .ZN(n918) );
  NOR2_X1 U1017 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1018 ( .A1(G28), .A2(n920), .ZN(n921) );
  XNOR2_X1 U1019 ( .A(KEYINPUT53), .B(n921), .ZN(n925) );
  XOR2_X1 U1020 ( .A(KEYINPUT120), .B(G34), .Z(n923) );
  XNOR2_X1 U1021 ( .A(G2084), .B(KEYINPUT54), .ZN(n922) );
  XNOR2_X1 U1022 ( .A(n923), .B(n922), .ZN(n924) );
  NAND2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n927) );
  XNOR2_X1 U1024 ( .A(G35), .B(G2090), .ZN(n926) );
  NOR2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n928) );
  XOR2_X1 U1026 ( .A(KEYINPUT55), .B(n928), .Z(n929) );
  NOR2_X1 U1027 ( .A1(G29), .A2(n929), .ZN(n930) );
  XNOR2_X1 U1028 ( .A(KEYINPUT121), .B(n930), .ZN(n1018) );
  XOR2_X1 U1029 ( .A(G16), .B(KEYINPUT124), .Z(n955) );
  XNOR2_X1 U1030 ( .A(KEYINPUT59), .B(KEYINPUT126), .ZN(n931) );
  XNOR2_X1 U1031 ( .A(n931), .B(G4), .ZN(n932) );
  XNOR2_X1 U1032 ( .A(G1348), .B(n932), .ZN(n939) );
  XNOR2_X1 U1033 ( .A(G1956), .B(G20), .ZN(n937) );
  XNOR2_X1 U1034 ( .A(G1981), .B(G6), .ZN(n934) );
  XNOR2_X1 U1035 ( .A(G1341), .B(G19), .ZN(n933) );
  NOR2_X1 U1036 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1037 ( .A(KEYINPUT125), .B(n935), .ZN(n936) );
  NOR2_X1 U1038 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1039 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1040 ( .A(n940), .B(KEYINPUT60), .ZN(n952) );
  XNOR2_X1 U1041 ( .A(G1986), .B(G24), .ZN(n945) );
  XNOR2_X1 U1042 ( .A(G1976), .B(G23), .ZN(n942) );
  XNOR2_X1 U1043 ( .A(G22), .B(G1971), .ZN(n941) );
  NOR2_X1 U1044 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1045 ( .A(KEYINPUT127), .B(n943), .ZN(n944) );
  NOR2_X1 U1046 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1047 ( .A(KEYINPUT58), .B(n946), .ZN(n950) );
  XNOR2_X1 U1048 ( .A(G1966), .B(G21), .ZN(n948) );
  XNOR2_X1 U1049 ( .A(G1961), .B(G5), .ZN(n947) );
  NOR2_X1 U1050 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1051 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1052 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1053 ( .A(n953), .B(KEYINPUT61), .ZN(n954) );
  NAND2_X1 U1054 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1055 ( .A1(G11), .A2(n956), .ZN(n1016) );
  XOR2_X1 U1056 ( .A(G2084), .B(G160), .Z(n957) );
  NOR2_X1 U1057 ( .A1(n958), .A2(n957), .ZN(n963) );
  NOR2_X1 U1058 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1059 ( .A(KEYINPUT113), .B(n961), .Z(n962) );
  NAND2_X1 U1060 ( .A1(n963), .A2(n962), .ZN(n964) );
  NOR2_X1 U1061 ( .A1(n965), .A2(n964), .ZN(n966) );
  XOR2_X1 U1062 ( .A(KEYINPUT114), .B(n966), .Z(n967) );
  NOR2_X1 U1063 ( .A1(n968), .A2(n967), .ZN(n974) );
  XNOR2_X1 U1064 ( .A(G2090), .B(G162), .ZN(n969) );
  XNOR2_X1 U1065 ( .A(n969), .B(KEYINPUT115), .ZN(n970) );
  NOR2_X1 U1066 ( .A1(n971), .A2(n970), .ZN(n972) );
  XOR2_X1 U1067 ( .A(KEYINPUT51), .B(n972), .Z(n973) );
  NAND2_X1 U1068 ( .A1(n974), .A2(n973), .ZN(n980) );
  XOR2_X1 U1069 ( .A(G2072), .B(n975), .Z(n977) );
  XOR2_X1 U1070 ( .A(G164), .B(G2078), .Z(n976) );
  NOR2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1072 ( .A(n978), .B(KEYINPUT50), .Z(n979) );
  NOR2_X1 U1073 ( .A1(n980), .A2(n979), .ZN(n981) );
  XOR2_X1 U1074 ( .A(KEYINPUT52), .B(n981), .Z(n982) );
  XNOR2_X1 U1075 ( .A(n982), .B(KEYINPUT116), .ZN(n983) );
  NOR2_X1 U1076 ( .A1(KEYINPUT55), .A2(n983), .ZN(n984) );
  XNOR2_X1 U1077 ( .A(n984), .B(KEYINPUT117), .ZN(n985) );
  NAND2_X1 U1078 ( .A1(n985), .A2(G29), .ZN(n1014) );
  XNOR2_X1 U1079 ( .A(KEYINPUT56), .B(G16), .ZN(n1012) );
  XNOR2_X1 U1080 ( .A(n986), .B(G1341), .ZN(n1005) );
  XNOR2_X1 U1081 ( .A(G1348), .B(n987), .ZN(n989) );
  NAND2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n1002) );
  XNOR2_X1 U1083 ( .A(G1956), .B(n990), .ZN(n992) );
  NAND2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n994) );
  XNOR2_X1 U1085 ( .A(G1971), .B(G303), .ZN(n993) );
  NOR2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n1000) );
  XOR2_X1 U1087 ( .A(n995), .B(KEYINPUT122), .Z(n998) );
  XNOR2_X1 U1088 ( .A(n996), .B(G171), .ZN(n997) );
  NOR2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NOR2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1092 ( .A(KEYINPUT123), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1010) );
  XOR2_X1 U1094 ( .A(G1966), .B(G168), .Z(n1006) );
  NOR2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1096 ( .A(KEYINPUT57), .B(n1008), .Z(n1009) );
  NAND2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1098 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1099 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NOR2_X1 U1100 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1101 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1102 ( .A(KEYINPUT62), .B(n1019), .Z(G311) );
  INV_X1 U1103 ( .A(G311), .ZN(G150) );
endmodule

