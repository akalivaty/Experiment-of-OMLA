//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 1 1 0 0 0 0 0 1 0 1 0 1 1 0 0 1 0 1 1 0 1 0 0 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 0 0 0 1 1 0 0 0 0 1 0 0 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:46 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1292, new_n1293, new_n1295, new_n1296, new_n1297,
    new_n1298, new_n1299, new_n1300, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357;
  INV_X1    g0000(.A(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G58), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT0), .ZN(new_n212));
  AND2_X1   g0012(.A1(KEYINPUT64), .A2(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(KEYINPUT64), .A2(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(G58), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(new_n201), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G50), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(new_n211), .A2(new_n212), .B1(new_n217), .B2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n222), .B1(new_n212), .B2(new_n211), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT65), .Z(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n225));
  INV_X1    g0025(.A(G244), .ZN(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT66), .B(G68), .ZN(new_n227));
  INV_X1    g0027(.A(G238), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n225), .B1(new_n202), .B2(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(KEYINPUT67), .ZN(new_n230));
  AOI22_X1  g0030(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n231));
  AOI22_X1  g0031(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n232));
  NAND3_X1  g0032(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n229), .A2(KEYINPUT67), .ZN(new_n234));
  OAI21_X1  g0034(.A(new_n209), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  OAI21_X1  g0035(.A(new_n224), .B1(KEYINPUT1), .B2(new_n235), .ZN(new_n236));
  AOI21_X1  g0036(.A(new_n236), .B1(KEYINPUT1), .B2(new_n235), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G264), .B(G270), .Z(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  NAND2_X1  g0045(.A1(G68), .A2(G77), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n203), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT68), .ZN(new_n248));
  XOR2_X1   g0048(.A(G50), .B(G58), .Z(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G87), .B(G97), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G107), .B(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n250), .B(new_n253), .ZN(G351));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(new_n216), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n215), .A2(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n218), .A2(KEYINPUT8), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT8), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G58), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n257), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G150), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G20), .A2(G33), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NOR3_X1   g0066(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n267));
  OAI22_X1  g0067(.A1(new_n264), .A2(new_n266), .B1(new_n267), .B2(new_n207), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n256), .B1(new_n263), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G50), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n270), .A2(new_n216), .A3(new_n255), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n206), .A2(G20), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G50), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n269), .B(new_n273), .C1(new_n274), .C2(new_n276), .ZN(new_n277));
  XNOR2_X1  g0077(.A(new_n277), .B(KEYINPUT9), .ZN(new_n278));
  AND2_X1   g0078(.A1(G33), .A2(G41), .ZN(new_n279));
  OAI21_X1  g0079(.A(G274), .B1(new_n279), .B2(new_n216), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n281));
  NOR3_X1   g0081(.A1(new_n280), .A2(KEYINPUT69), .A3(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT69), .ZN(new_n283));
  INV_X1    g0083(.A(G274), .ZN(new_n284));
  AND2_X1   g0084(.A1(G1), .A2(G13), .ZN(new_n285));
  NAND2_X1  g0085(.A1(G33), .A2(G41), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n281), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n283), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n282), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n286), .A2(G1), .A3(G13), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(new_n281), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n290), .B1(G226), .B2(new_n293), .ZN(new_n294));
  OR2_X1    g0094(.A1(KEYINPUT3), .A2(G33), .ZN(new_n295));
  NAND2_X1  g0095(.A1(KEYINPUT3), .A2(G33), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G1698), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n297), .A2(G222), .A3(new_n298), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n299), .B(KEYINPUT70), .ZN(new_n300));
  AND2_X1   g0100(.A1(KEYINPUT3), .A2(G33), .ZN(new_n301));
  NOR2_X1   g0101(.A1(KEYINPUT3), .A2(G33), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n303), .A2(new_n298), .ZN(new_n304));
  AOI22_X1  g0104(.A1(new_n304), .A2(G223), .B1(G77), .B2(new_n303), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n300), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n294), .B1(new_n306), .B2(new_n291), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G200), .ZN(new_n308));
  OAI211_X1 g0108(.A(G190), .B(new_n294), .C1(new_n306), .C2(new_n291), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n278), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT10), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT10), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n278), .A2(new_n308), .A3(new_n312), .A4(new_n309), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  OR2_X1    g0114(.A1(new_n307), .A2(G179), .ZN(new_n315));
  INV_X1    g0115(.A(G169), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n307), .A2(new_n316), .ZN(new_n317));
  AND3_X1   g0117(.A1(new_n315), .A2(new_n277), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n314), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n261), .A2(new_n275), .ZN(new_n321));
  OAI22_X1  g0121(.A1(new_n321), .A2(new_n274), .B1(new_n270), .B2(new_n261), .ZN(new_n322));
  XNOR2_X1  g0122(.A(new_n322), .B(KEYINPUT74), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT7), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n215), .A2(new_n303), .A3(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n295), .A2(new_n207), .A3(new_n296), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(KEYINPUT7), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n325), .A2(new_n327), .A3(G68), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n219), .B1(new_n227), .B2(new_n218), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(G20), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n265), .A2(G159), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n328), .A2(KEYINPUT16), .A3(new_n330), .A4(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n256), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n329), .A2(G20), .B1(G159), .B2(new_n265), .ZN(new_n334));
  OR2_X1    g0134(.A1(KEYINPUT64), .A2(G20), .ZN(new_n335));
  NAND2_X1  g0135(.A1(KEYINPUT64), .A2(G20), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(KEYINPUT7), .B1(new_n337), .B2(new_n297), .ZN(new_n338));
  INV_X1    g0138(.A(new_n227), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n303), .A2(new_n324), .A3(new_n207), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(KEYINPUT16), .B1(new_n334), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n323), .B1(new_n333), .B2(new_n342), .ZN(new_n343));
  AND3_X1   g0143(.A1(new_n291), .A2(G232), .A3(new_n281), .ZN(new_n344));
  NAND2_X1  g0144(.A1(G33), .A2(G87), .ZN(new_n345));
  INV_X1    g0145(.A(G226), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G1698), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n347), .B1(G223), .B2(G1698), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n345), .B1(new_n348), .B2(new_n303), .ZN(new_n349));
  INV_X1    g0149(.A(new_n291), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n344), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(G179), .ZN(new_n352));
  OAI21_X1  g0152(.A(KEYINPUT69), .B1(new_n280), .B2(new_n281), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n287), .A2(new_n283), .A3(new_n288), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AND3_X1   g0155(.A1(new_n351), .A2(new_n352), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(G169), .B1(new_n351), .B2(new_n355), .ZN(new_n357));
  NOR3_X1   g0157(.A1(new_n356), .A2(new_n357), .A3(KEYINPUT75), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT75), .ZN(new_n359));
  NOR2_X1   g0159(.A1(G223), .A2(G1698), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n360), .B1(new_n346), .B2(G1698), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n361), .A2(new_n297), .B1(G33), .B2(G87), .ZN(new_n362));
  INV_X1    g0162(.A(G232), .ZN(new_n363));
  OAI22_X1  g0163(.A1(new_n362), .A2(new_n291), .B1(new_n363), .B2(new_n292), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n316), .B1(new_n364), .B2(new_n290), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n351), .A2(new_n352), .A3(new_n355), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n359), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n343), .B1(new_n358), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT18), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT18), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n370), .B(new_n343), .C1(new_n358), .C2(new_n367), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT17), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n351), .A2(new_n355), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(G200), .ZN(new_n374));
  INV_X1    g0174(.A(G190), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n374), .B1(new_n375), .B2(new_n373), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n372), .B1(new_n343), .B2(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n373), .A2(new_n375), .ZN(new_n378));
  INV_X1    g0178(.A(G200), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n379), .B1(new_n351), .B2(new_n355), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n334), .A2(new_n341), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT16), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n384), .A2(new_n256), .A3(new_n332), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n381), .A2(new_n385), .A3(KEYINPUT17), .A4(new_n323), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n369), .A2(new_n371), .A3(new_n377), .A4(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT72), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n201), .A2(KEYINPUT66), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT66), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(G68), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n389), .A2(new_n391), .A3(G20), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT12), .ZN(new_n394));
  INV_X1    g0194(.A(G13), .ZN(new_n395));
  NOR3_X1   g0195(.A1(new_n394), .A2(new_n395), .A3(G1), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n395), .A2(G1), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n397), .A2(G20), .A3(new_n201), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n393), .A2(new_n396), .B1(new_n398), .B2(new_n394), .ZN(new_n399));
  INV_X1    g0199(.A(new_n256), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n201), .B1(new_n206), .B2(G20), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n400), .A2(new_n270), .A3(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n388), .B1(new_n399), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n398), .A2(new_n394), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n227), .A2(new_n396), .A3(G20), .ZN(new_n405));
  AND4_X1   g0205(.A1(new_n388), .A2(new_n402), .A3(new_n404), .A4(new_n405), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n335), .A2(G33), .A3(G77), .A4(new_n336), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n265), .A2(G50), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n407), .A2(new_n392), .A3(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT11), .ZN(new_n410));
  AND3_X1   g0210(.A1(new_n409), .A2(new_n410), .A3(new_n256), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n410), .B1(new_n409), .B2(new_n256), .ZN(new_n412));
  OAI22_X1  g0212(.A1(new_n403), .A2(new_n406), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT14), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n346), .A2(new_n298), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n363), .A2(G1698), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n415), .B(new_n416), .C1(new_n301), .C2(new_n302), .ZN(new_n417));
  INV_X1    g0217(.A(G33), .ZN(new_n418));
  INV_X1    g0218(.A(G97), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n417), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n350), .ZN(new_n423));
  XOR2_X1   g0223(.A(KEYINPUT71), .B(KEYINPUT13), .Z(new_n424));
  AND3_X1   g0224(.A1(new_n291), .A2(G238), .A3(new_n281), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  AND4_X1   g0226(.A1(new_n355), .A2(new_n423), .A3(new_n424), .A4(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n425), .B1(new_n422), .B2(new_n350), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n424), .B1(new_n428), .B2(new_n355), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n414), .B(G169), .C1(new_n427), .C2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n428), .A2(new_n355), .A3(new_n424), .ZN(new_n431));
  NOR2_X1   g0231(.A1(G226), .A2(G1698), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n432), .B1(new_n363), .B2(G1698), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n420), .B1(new_n433), .B2(new_n297), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n426), .B1(new_n434), .B2(new_n291), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n435), .A2(new_n290), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT13), .ZN(new_n437));
  OAI211_X1 g0237(.A(G179), .B(new_n431), .C1(new_n436), .C2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n430), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n424), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(new_n435), .B2(new_n290), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n431), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n414), .B1(new_n442), .B2(G169), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n413), .B1(new_n439), .B2(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n437), .B1(new_n428), .B2(new_n355), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n427), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n413), .B1(new_n446), .B2(G190), .ZN(new_n447));
  OAI21_X1  g0247(.A(G200), .B1(new_n427), .B2(new_n429), .ZN(new_n448));
  AOI21_X1  g0248(.A(KEYINPUT73), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n413), .ZN(new_n450));
  OAI211_X1 g0250(.A(G190), .B(new_n431), .C1(new_n436), .C2(new_n437), .ZN(new_n451));
  AND4_X1   g0251(.A1(KEYINPUT73), .A2(new_n450), .A3(new_n451), .A4(new_n448), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n444), .B1(new_n449), .B2(new_n452), .ZN(new_n453));
  OAI22_X1  g0253(.A1(new_n262), .A2(new_n266), .B1(new_n215), .B2(new_n202), .ZN(new_n454));
  XNOR2_X1  g0254(.A(KEYINPUT15), .B(G87), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n257), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n256), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n274), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n202), .B1(new_n206), .B2(G20), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n458), .A2(new_n459), .B1(new_n202), .B2(new_n271), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(G232), .A2(G1698), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n298), .A2(G238), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n297), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n464), .B(new_n350), .C1(G107), .C2(new_n297), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n293), .A2(G244), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n465), .A2(new_n355), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n461), .B1(G200), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n468), .B1(new_n375), .B2(new_n467), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n467), .A2(new_n316), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n465), .A2(new_n355), .A3(new_n352), .A4(new_n466), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n470), .A2(new_n471), .A3(new_n461), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  NOR4_X1   g0273(.A1(new_n320), .A2(new_n387), .A3(new_n453), .A4(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT19), .ZN(new_n476));
  AND2_X1   g0276(.A1(new_n476), .A2(KEYINPUT80), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n476), .A2(KEYINPUT80), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n335), .A2(G33), .A3(G97), .A4(new_n336), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n297), .A2(new_n215), .A3(G68), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NOR3_X1   g0283(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n420), .B1(new_n477), .B2(new_n478), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n484), .B1(new_n485), .B2(new_n215), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n256), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n455), .A2(new_n271), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n206), .A2(G33), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n458), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n455), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n487), .A2(new_n488), .A3(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(G45), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n495), .A2(G1), .ZN(new_n496));
  INV_X1    g0296(.A(G250), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n291), .A2(new_n498), .B1(new_n287), .B2(new_n496), .ZN(new_n499));
  NOR2_X1   g0299(.A1(G238), .A2(G1698), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n500), .B1(new_n226), .B2(G1698), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n501), .A2(new_n297), .B1(G33), .B2(G116), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n499), .B1(new_n502), .B2(new_n291), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n352), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n503), .A2(new_n316), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n494), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n504), .A2(new_n379), .ZN(new_n508));
  INV_X1    g0308(.A(G87), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n490), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n499), .B(G190), .C1(new_n502), .C2(new_n291), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n487), .A2(new_n511), .A3(new_n488), .A4(new_n512), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n507), .B1(new_n508), .B2(new_n513), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n338), .A2(G107), .A3(new_n340), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT6), .ZN(new_n516));
  NOR3_X1   g0316(.A1(new_n516), .A2(new_n419), .A3(G107), .ZN(new_n517));
  XNOR2_X1  g0317(.A(G97), .B(G107), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n517), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  OAI22_X1  g0319(.A1(new_n519), .A2(new_n215), .B1(new_n202), .B2(new_n266), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n256), .B1(new_n515), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n270), .A2(G97), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n522), .B1(new_n491), .B2(G97), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  AND2_X1   g0324(.A1(KEYINPUT5), .A2(G41), .ZN(new_n525));
  NOR2_X1   g0325(.A1(KEYINPUT5), .A2(G41), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n496), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n527), .A2(G257), .A3(new_n291), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(KEYINPUT78), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n527), .A2(new_n280), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT78), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n527), .A2(new_n532), .A3(G257), .A4(new_n291), .ZN(new_n533));
  AND3_X1   g0333(.A1(new_n529), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n226), .A2(G1698), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(new_n301), .B2(new_n302), .ZN(new_n536));
  NOR2_X1   g0336(.A1(KEYINPUT76), .A2(KEYINPUT4), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OAI221_X1 g0338(.A(new_n535), .B1(KEYINPUT76), .B2(KEYINPUT4), .C1(new_n301), .C2(new_n302), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n297), .A2(G250), .A3(G1698), .ZN(new_n540));
  NAND2_X1  g0340(.A1(G33), .A2(G283), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n538), .A2(new_n539), .A3(new_n540), .A4(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT77), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n542), .A2(new_n543), .A3(new_n350), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n543), .B1(new_n542), .B2(new_n350), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n534), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n524), .B1(new_n546), .B2(G200), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n542), .A2(new_n350), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n534), .A2(G190), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(KEYINPUT79), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT79), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n534), .A2(new_n551), .A3(G190), .A4(new_n548), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n547), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n534), .A2(new_n548), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n555), .A2(new_n316), .B1(new_n521), .B2(new_n523), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n352), .B(new_n534), .C1(new_n544), .C2(new_n545), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(G107), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n271), .A2(KEYINPUT25), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(KEYINPUT25), .B1(new_n271), .B2(new_n560), .ZN(new_n562));
  OAI22_X1  g0362(.A1(new_n490), .A2(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT22), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n335), .B(new_n336), .C1(new_n301), .C2(new_n302), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n564), .B1(new_n565), .B2(new_n509), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT23), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n560), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n568), .B1(new_n335), .B2(new_n336), .ZN(new_n569));
  AOI21_X1  g0369(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n570));
  OAI22_X1  g0370(.A1(new_n570), .A2(G20), .B1(new_n567), .B2(new_n560), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n297), .A2(new_n215), .A3(KEYINPUT22), .A4(G87), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n566), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(KEYINPUT24), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT24), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n566), .A2(new_n572), .A3(new_n576), .A4(new_n573), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n563), .B1(new_n578), .B2(new_n256), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n497), .A2(G1698), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(new_n301), .B2(new_n302), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT81), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(G33), .A2(G294), .ZN(new_n584));
  OAI211_X1 g0384(.A(G257), .B(G1698), .C1(new_n301), .C2(new_n302), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n580), .B(KEYINPUT81), .C1(new_n302), .C2(new_n301), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n583), .A2(new_n584), .A3(new_n585), .A4(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n350), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n527), .A2(G264), .A3(new_n291), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n588), .A2(new_n375), .A3(new_n531), .A4(new_n590), .ZN(new_n591));
  AOI211_X1 g0391(.A(new_n530), .B(new_n589), .C1(new_n587), .C2(new_n350), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n591), .B1(new_n592), .B2(G200), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n579), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n588), .A2(new_n531), .A3(new_n590), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n316), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n589), .B1(new_n587), .B2(new_n350), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n597), .A2(new_n352), .A3(new_n531), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n400), .B1(new_n575), .B2(new_n577), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n596), .B(new_n598), .C1(new_n599), .C2(new_n563), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n594), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(KEYINPUT82), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT82), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n594), .A2(new_n600), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n206), .A2(G45), .ZN(new_n605));
  OR2_X1    g0405(.A1(KEYINPUT5), .A2(G41), .ZN(new_n606));
  NAND2_X1  g0406(.A1(KEYINPUT5), .A2(G41), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n608), .A2(new_n350), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n530), .B1(new_n609), .B2(G270), .ZN(new_n610));
  OAI211_X1 g0410(.A(G257), .B(new_n298), .C1(new_n301), .C2(new_n302), .ZN(new_n611));
  OAI211_X1 g0411(.A(G264), .B(G1698), .C1(new_n301), .C2(new_n302), .ZN(new_n612));
  INV_X1    g0412(.A(G303), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n611), .B(new_n612), .C1(new_n613), .C2(new_n297), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n350), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(G116), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n271), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n458), .A2(G116), .A3(new_n489), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n418), .A2(G97), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n335), .A2(new_n620), .A3(new_n336), .A4(new_n541), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n255), .A2(new_n216), .B1(G20), .B2(new_n617), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n621), .A2(KEYINPUT20), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(KEYINPUT20), .B1(new_n621), .B2(new_n622), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n618), .B(new_n619), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n616), .A2(KEYINPUT21), .A3(new_n625), .A4(G169), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n625), .A2(G179), .A3(new_n615), .A4(new_n610), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n316), .B1(new_n610), .B2(new_n615), .ZN(new_n629));
  AOI21_X1  g0429(.A(KEYINPUT21), .B1(new_n629), .B2(new_n625), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n625), .B1(new_n616), .B2(G200), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(new_n375), .B2(new_n616), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n602), .A2(new_n604), .A3(new_n634), .ZN(new_n635));
  NOR4_X1   g0435(.A1(new_n475), .A2(new_n514), .A3(new_n559), .A4(new_n635), .ZN(G372));
  AND2_X1   g0436(.A1(new_n369), .A2(new_n371), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n472), .A2(KEYINPUT85), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT85), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n470), .A2(new_n639), .A3(new_n461), .A4(new_n471), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n447), .A2(KEYINPUT73), .A3(new_n448), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n450), .A2(new_n451), .A3(new_n448), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT73), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n641), .B1(new_n642), .B2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n444), .ZN(new_n647));
  OAI21_X1  g0447(.A(KEYINPUT86), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n377), .A2(new_n386), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NOR3_X1   g0450(.A1(new_n646), .A2(new_n647), .A3(KEYINPUT86), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n637), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT87), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OAI211_X1 g0454(.A(KEYINPUT87), .B(new_n637), .C1(new_n650), .C2(new_n651), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(new_n655), .A3(new_n314), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n656), .A2(new_n319), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n556), .A2(new_n557), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n494), .A2(new_n505), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT83), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n660), .B1(new_n502), .B2(new_n291), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n226), .A2(G1698), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n662), .B1(G238), .B2(G1698), .ZN(new_n663));
  OAI22_X1  g0463(.A1(new_n663), .A2(new_n303), .B1(new_n418), .B2(new_n617), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n664), .A2(KEYINPUT83), .A3(new_n350), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n499), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n316), .ZN(new_n668));
  AND4_X1   g0468(.A1(new_n487), .A2(new_n511), .A3(new_n488), .A4(new_n512), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n667), .A2(G200), .ZN(new_n670));
  AOI22_X1  g0470(.A1(new_n659), .A2(new_n668), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT26), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n658), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n659), .A2(new_n668), .ZN(new_n674));
  OAI21_X1  g0474(.A(KEYINPUT26), .B1(new_n558), .B2(new_n514), .ZN(new_n675));
  AND3_X1   g0475(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n596), .A2(new_n598), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(new_n579), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n616), .A2(G169), .A3(new_n625), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT21), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n681), .A2(new_n627), .A3(new_n626), .ZN(new_n682));
  OAI21_X1  g0482(.A(KEYINPUT84), .B1(new_n678), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n494), .A2(new_n505), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n498), .A2(new_n291), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n280), .B2(new_n605), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n686), .B1(new_n661), .B2(new_n665), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(G169), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n379), .ZN(new_n689));
  OAI22_X1  g0489(.A1(new_n684), .A2(new_n688), .B1(new_n689), .B2(new_n513), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n690), .B1(new_n579), .B2(new_n593), .ZN(new_n691));
  AOI22_X1  g0491(.A1(new_n547), .A2(new_n553), .B1(new_n556), .B2(new_n557), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT84), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n631), .A2(new_n693), .A3(new_n600), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n683), .A2(new_n691), .A3(new_n692), .A4(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n676), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n474), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n657), .A2(new_n697), .ZN(G369));
  NAND2_X1  g0498(.A1(new_n215), .A2(new_n397), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n699), .A2(KEYINPUT27), .ZN(new_n700));
  OAI21_X1  g0500(.A(G213), .B1(new_n699), .B2(KEYINPUT27), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(G343), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n704), .A2(new_n625), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n682), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n631), .A2(new_n633), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n706), .B1(new_n707), .B2(new_n705), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(G330), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  OAI211_X1 g0512(.A(new_n602), .B(new_n604), .C1(new_n579), .C2(new_n703), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n678), .A2(new_n704), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n682), .A2(KEYINPUT88), .A3(new_n703), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(KEYINPUT88), .B1(new_n682), .B2(new_n703), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n722), .B1(new_n713), .B2(new_n714), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n723), .B1(new_n678), .B2(new_n703), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n718), .A2(new_n724), .ZN(G399));
  INV_X1    g0525(.A(new_n210), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(G41), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n484), .A2(new_n617), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n728), .A2(G1), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n731), .B1(new_n220), .B2(new_n728), .ZN(new_n732));
  XNOR2_X1  g0532(.A(new_n732), .B(KEYINPUT28), .ZN(new_n733));
  AOI21_X1  g0533(.A(G179), .B1(new_n610), .B2(new_n615), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n546), .A2(new_n595), .A3(new_n667), .A4(new_n734), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n534), .A2(new_n548), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n597), .A2(new_n504), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n610), .A2(new_n615), .A3(G179), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n736), .A2(new_n737), .A3(KEYINPUT30), .A4(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT30), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n534), .A2(new_n597), .A3(new_n504), .A4(new_n548), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n741), .B1(new_n742), .B2(new_n738), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n735), .A2(new_n740), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(new_n704), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT31), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n744), .A2(KEYINPUT31), .A3(new_n704), .ZN(new_n748));
  INV_X1    g0548(.A(new_n508), .ZN(new_n749));
  AOI22_X1  g0549(.A1(new_n659), .A2(new_n506), .B1(new_n749), .B2(new_n669), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n692), .A2(new_n750), .A3(new_n703), .ZN(new_n751));
  OAI211_X1 g0551(.A(new_n747), .B(new_n748), .C1(new_n635), .C2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G330), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n704), .B1(new_n676), .B2(new_n695), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(KEYINPUT29), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n631), .A2(new_n600), .ZN(new_n756));
  AND4_X1   g0556(.A1(new_n692), .A2(new_n594), .A3(new_n756), .A4(new_n671), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n658), .A2(new_n750), .A3(new_n672), .ZN(new_n758));
  OAI21_X1  g0558(.A(KEYINPUT26), .B1(new_n558), .B2(new_n690), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n758), .A2(new_n759), .A3(new_n674), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n703), .B1(new_n757), .B2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT29), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n753), .B1(new_n755), .B2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n733), .B1(new_n765), .B2(G1), .ZN(G364));
  NOR2_X1   g0566(.A1(G13), .A2(G33), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(G20), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n709), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n726), .A2(new_n303), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G355), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(G116), .B2(new_n210), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n250), .A2(G45), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n726), .A2(new_n297), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n776), .B1(new_n495), .B2(new_n221), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n773), .B1(new_n774), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n216), .B1(G20), .B2(new_n316), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n769), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n337), .A2(new_n395), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G45), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n728), .A2(G1), .A3(new_n784), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT89), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n782), .A2(new_n787), .ZN(new_n788));
  NOR3_X1   g0588(.A1(G179), .A2(G190), .A3(G200), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n337), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n297), .B1(new_n791), .B2(G329), .ZN(new_n792));
  INV_X1    g0592(.A(G311), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n215), .A2(new_n352), .ZN(new_n794));
  NOR2_X1   g0594(.A1(G190), .A2(G200), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n792), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n794), .A2(G200), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n375), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n797), .B1(G326), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n798), .A2(G190), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(KEYINPUT91), .B(KEYINPUT33), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n803), .B(G317), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n800), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n379), .A2(G179), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT90), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n207), .A2(new_n375), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n375), .A2(G200), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n794), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(G322), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n809), .A2(new_n613), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n215), .A2(G190), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n807), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(G283), .ZN(new_n816));
  INV_X1    g0616(.A(G294), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n215), .B1(new_n352), .B2(new_n810), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n815), .A2(new_n816), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NOR3_X1   g0619(.A1(new_n805), .A2(new_n813), .A3(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n799), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n297), .B1(new_n560), .B2(new_n815), .C1(new_n821), .C2(new_n272), .ZN(new_n822));
  INV_X1    g0622(.A(G159), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n790), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT32), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(new_n802), .B2(new_n201), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n809), .A2(new_n509), .B1(new_n811), .B2(new_n218), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n796), .A2(new_n202), .B1(new_n818), .B2(new_n419), .ZN(new_n828));
  NOR4_X1   g0628(.A1(new_n822), .A2(new_n826), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  OR2_X1    g0629(.A1(new_n820), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(KEYINPUT92), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(new_n779), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n830), .A2(KEYINPUT92), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n770), .B(new_n788), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n709), .A2(new_n710), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n835), .A2(new_n712), .A3(new_n787), .ZN(new_n836));
  AND2_X1   g0636(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(G396));
  NAND2_X1  g0638(.A1(new_n704), .A2(new_n461), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n469), .A2(new_n472), .A3(new_n839), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n638), .A2(new_n461), .A3(new_n640), .A4(new_n704), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OR2_X1    g0642(.A1(new_n754), .A2(new_n842), .ZN(new_n843));
  AND4_X1   g0643(.A1(new_n692), .A2(new_n683), .A3(new_n691), .A4(new_n694), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n673), .A2(new_n675), .A3(new_n674), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n703), .B(new_n842), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n786), .B1(new_n847), .B2(new_n753), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n753), .B2(new_n847), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n815), .A2(new_n509), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(G311), .B2(new_n791), .ZN(new_n851));
  XOR2_X1   g0651(.A(new_n851), .B(KEYINPUT93), .Z(new_n852));
  OAI22_X1  g0652(.A1(new_n809), .A2(new_n560), .B1(new_n796), .B2(new_n617), .ZN(new_n853));
  INV_X1    g0653(.A(new_n811), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n853), .B1(G294), .B2(new_n854), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n303), .B1(new_n419), .B2(new_n818), .C1(new_n821), .C2(new_n613), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n856), .B1(G283), .B2(new_n801), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n852), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n796), .ZN(new_n859));
  AOI22_X1  g0659(.A1(G159), .A2(new_n859), .B1(new_n854), .B2(G143), .ZN(new_n860));
  INV_X1    g0660(.A(G137), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n860), .B1(new_n802), .B2(new_n264), .C1(new_n861), .C2(new_n821), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n862), .B(KEYINPUT34), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n864), .A2(KEYINPUT94), .ZN(new_n865));
  INV_X1    g0665(.A(G132), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n297), .B1(new_n790), .B2(new_n866), .ZN(new_n867));
  OAI22_X1  g0667(.A1(new_n815), .A2(new_n201), .B1(new_n218), .B2(new_n818), .ZN(new_n868));
  INV_X1    g0668(.A(new_n809), .ZN(new_n869));
  AOI211_X1 g0669(.A(new_n867), .B(new_n868), .C1(G50), .C2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n864), .B2(KEYINPUT94), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n858), .B1(new_n865), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n779), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n779), .A2(new_n767), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n787), .B1(new_n202), .B2(new_n874), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n873), .B(new_n875), .C1(new_n768), .C2(new_n842), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n849), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(G384));
  INV_X1    g0678(.A(new_n519), .ZN(new_n879));
  OR2_X1    g0679(.A1(new_n879), .A2(KEYINPUT35), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(KEYINPUT35), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n880), .A2(G116), .A3(new_n217), .A4(new_n881), .ZN(new_n882));
  XNOR2_X1  g0682(.A(KEYINPUT95), .B(KEYINPUT36), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n882), .B(new_n883), .ZN(new_n884));
  AOI211_X1 g0684(.A(new_n202), .B(new_n220), .C1(new_n339), .C2(G58), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n885), .A2(KEYINPUT96), .B1(new_n272), .B2(G68), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n886), .B1(KEYINPUT96), .B2(new_n885), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n206), .A2(G13), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n884), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT39), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT98), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT37), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n381), .A2(new_n385), .A3(new_n323), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n343), .A2(new_n702), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n368), .A2(new_n892), .A3(new_n893), .A4(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT74), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n322), .B(new_n897), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n332), .A2(new_n256), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n898), .B1(new_n899), .B2(new_n384), .ZN(new_n900));
  INV_X1    g0700(.A(new_n322), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT16), .B1(new_n334), .B2(new_n328), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n901), .B1(new_n333), .B2(new_n902), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n900), .A2(new_n381), .B1(new_n903), .B2(new_n702), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n903), .B1(new_n358), .B2(new_n367), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n892), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n891), .B1(new_n896), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n903), .A2(new_n702), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n387), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n893), .A2(new_n908), .ZN(new_n911));
  INV_X1    g0711(.A(new_n902), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n912), .A2(new_n256), .A3(new_n332), .ZN(new_n913));
  OAI21_X1  g0713(.A(KEYINPUT75), .B1(new_n356), .B2(new_n357), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n365), .A2(new_n359), .A3(new_n366), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n901), .A2(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT37), .B1(new_n911), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n917), .A2(KEYINPUT98), .A3(new_n895), .ZN(new_n918));
  AND4_X1   g0718(.A1(KEYINPUT38), .A2(new_n907), .A3(new_n910), .A4(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n894), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT99), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n377), .A2(new_n386), .A3(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n922), .A2(new_n369), .A3(new_n371), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n921), .B1(new_n377), .B2(new_n386), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n920), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n368), .A2(new_n893), .A3(new_n894), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(KEYINPUT37), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n895), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT38), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n890), .B1(new_n919), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n647), .A2(new_n703), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT38), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n910), .A2(new_n918), .ZN(new_n934));
  AOI21_X1  g0734(.A(KEYINPUT98), .B1(new_n917), .B2(new_n895), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n907), .A2(KEYINPUT38), .A3(new_n910), .A4(new_n918), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n936), .A2(KEYINPUT39), .A3(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n930), .A2(new_n932), .A3(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n637), .A2(new_n702), .ZN(new_n940));
  NOR3_X1   g0740(.A1(new_n450), .A2(KEYINPUT97), .A3(new_n703), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT97), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(new_n413), .B2(new_n704), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n453), .A2(new_n945), .ZN(new_n946));
  OAI211_X1 g0746(.A(new_n944), .B(new_n444), .C1(new_n449), .C2(new_n452), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n472), .A2(new_n704), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n949), .B1(new_n846), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n936), .A2(new_n937), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n940), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT100), .ZN(new_n955));
  AND3_X1   g0755(.A1(new_n939), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n955), .B1(new_n939), .B2(new_n954), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OR3_X1    g0758(.A1(new_n475), .A2(new_n755), .A3(new_n763), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n657), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n958), .B(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n842), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n962), .B1(new_n946), .B2(new_n947), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n752), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT101), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n963), .A2(new_n752), .A3(KEYINPUT101), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n953), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT40), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n919), .A2(new_n929), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n963), .A2(new_n752), .A3(KEYINPUT40), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n970), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n474), .A2(new_n752), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n973), .A2(new_n974), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n975), .A2(G330), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n961), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n206), .B2(new_n783), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n961), .A2(new_n977), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n889), .B1(new_n979), .B2(new_n980), .ZN(G367));
  AOI21_X1  g0781(.A(new_n703), .B1(new_n521), .B2(new_n523), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n559), .A2(new_n982), .B1(new_n558), .B2(new_n703), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT103), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  OAI221_X1 g0785(.A(KEYINPUT103), .B1(new_n558), .B2(new_n703), .C1(new_n559), .C2(new_n982), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n558), .B1(new_n988), .B2(new_n600), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT42), .ZN(new_n990));
  INV_X1    g0790(.A(new_n722), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n715), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n990), .B1(new_n988), .B2(new_n992), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n987), .A2(KEYINPUT42), .A3(new_n723), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n703), .A2(new_n989), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n487), .A2(new_n488), .A3(new_n511), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n704), .A2(new_n996), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n674), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n671), .A2(new_n997), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AND2_X1   g0800(.A1(new_n1000), .A2(KEYINPUT43), .ZN(new_n1001));
  XOR2_X1   g0801(.A(KEYINPUT102), .B(KEYINPUT43), .Z(new_n1002));
  NOR2_X1   g0802(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  OR3_X1    g0803(.A1(new_n995), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n718), .A2(new_n988), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n995), .A2(new_n1003), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1005), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n727), .B(KEYINPUT41), .Z(new_n1011));
  INV_X1    g0811(.A(KEYINPUT44), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1012), .A2(KEYINPUT104), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(KEYINPUT104), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n985), .A2(new_n986), .A3(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1013), .B1(new_n724), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n678), .A2(new_n703), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n992), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1013), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1018), .A2(new_n988), .A3(new_n1019), .A4(new_n1014), .ZN(new_n1020));
  AOI21_X1  g0820(.A(KEYINPUT45), .B1(new_n724), .B2(new_n987), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n992), .A2(new_n987), .A3(new_n1017), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT45), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1016), .B(new_n1020), .C1(new_n1021), .C2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n717), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1022), .B(new_n1023), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1027), .A2(new_n718), .A3(new_n1016), .A4(new_n1020), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1025), .A2(KEYINPUT105), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT106), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n712), .B1(new_n992), .B2(new_n1032), .ZN(new_n1033));
  NOR3_X1   g0833(.A1(new_n723), .A2(new_n711), .A3(KEYINPUT106), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n1033), .A2(new_n1034), .B1(new_n715), .B2(new_n991), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n992), .A2(new_n1032), .A3(new_n712), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n715), .A2(new_n991), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n711), .B1(new_n723), .B2(KEYINPUT106), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n764), .B1(new_n1035), .B2(new_n1039), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT107), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1025), .A2(KEYINPUT105), .A3(new_n718), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1031), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1011), .B1(new_n1043), .B2(new_n765), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n784), .A2(G1), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1010), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n815), .A2(new_n202), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n809), .A2(new_n218), .B1(new_n201), .B2(new_n818), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n1047), .B(new_n1048), .C1(G50), .C2(new_n859), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n297), .B1(new_n861), .B2(new_n790), .C1(new_n811), .C2(new_n264), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(G143), .B2(new_n799), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1049), .B(new_n1051), .C1(new_n823), .C2(new_n802), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n809), .A2(new_n617), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT46), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n817), .A2(new_n802), .B1(new_n821), .B2(new_n793), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n815), .A2(new_n419), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n297), .B1(new_n791), .B2(G317), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n613), .B2(new_n811), .ZN(new_n1058));
  OR4_X1    g0858(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .A4(new_n1058), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n796), .A2(new_n816), .B1(new_n818), .B2(new_n560), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1060), .B(KEYINPUT108), .Z(new_n1061));
  OAI21_X1  g0861(.A(new_n1052), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT47), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n779), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n998), .A2(new_n999), .A3(new_n769), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n780), .B1(new_n210), .B2(new_n455), .C1(new_n776), .C2(new_n244), .ZN(new_n1066));
  AND2_X1   g0866(.A1(new_n786), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1064), .A2(new_n1065), .A3(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1046), .A2(new_n1068), .ZN(G387));
  OAI221_X1 g0869(.A(new_n297), .B1(new_n419), .B2(new_n815), .C1(new_n821), .C2(new_n823), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n261), .B2(new_n801), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n818), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n492), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1073), .B1(new_n811), .B2(new_n272), .C1(new_n201), .C2(new_n796), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n809), .A2(new_n202), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(G150), .B2(new_n791), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1074), .B1(KEYINPUT109), .B2(new_n1076), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1071), .B(new_n1077), .C1(KEYINPUT109), .C2(new_n1076), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n297), .B1(new_n791), .B2(G326), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n809), .A2(new_n817), .B1(new_n816), .B2(new_n818), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(G303), .A2(new_n859), .B1(new_n854), .B2(G317), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n1081), .B1(new_n802), .B2(new_n793), .C1(new_n812), .C2(new_n821), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT48), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1080), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n1083), .B2(new_n1082), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT49), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n1079), .B1(new_n617), .B2(new_n815), .C1(new_n1085), .C2(new_n1086), .ZN(new_n1087));
  AND2_X1   g0887(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1078), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n779), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n716), .A2(new_n769), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n771), .A2(new_n729), .B1(new_n560), .B2(new_n726), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n241), .A2(new_n495), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n261), .A2(new_n272), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT50), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n730), .A2(new_n495), .A3(new_n246), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n775), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1092), .B1(new_n1093), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n787), .B1(new_n1098), .B2(new_n780), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1090), .A2(new_n1091), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1045), .ZN(new_n1101));
  AND2_X1   g0901(.A1(new_n1035), .A2(new_n1039), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1035), .A2(new_n764), .A3(new_n1039), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n728), .B1(new_n1103), .B2(KEYINPUT110), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(KEYINPUT110), .B2(new_n1103), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n1100), .B1(new_n1101), .B2(new_n1102), .C1(new_n1105), .C2(new_n1041), .ZN(G393));
  INV_X1    g0906(.A(KEYINPUT107), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1040), .B(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n728), .B1(new_n1108), .B2(new_n1029), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1043), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n297), .B1(new_n791), .B2(G322), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n1111), .B1(new_n809), .B2(new_n816), .C1(new_n560), .C2(new_n815), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT114), .ZN(new_n1113));
  OR2_X1    g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n796), .A2(new_n817), .B1(new_n818), .B2(new_n617), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(G303), .B2(new_n801), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1114), .A2(new_n1115), .A3(new_n1117), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n799), .A2(G317), .B1(new_n854), .B2(G311), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT52), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n303), .B(new_n850), .C1(G143), .C2(new_n791), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n809), .A2(new_n227), .B1(new_n796), .B2(new_n262), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n818), .A2(new_n202), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1121), .B(new_n1124), .C1(new_n272), .C2(new_n802), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n799), .A2(G150), .B1(new_n854), .B2(G159), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT51), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n1118), .A2(new_n1120), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n1128), .A2(new_n779), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n780), .B1(new_n419), .B2(new_n210), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(new_n775), .B2(new_n253), .ZN(new_n1131));
  XOR2_X1   g0931(.A(new_n1131), .B(KEYINPUT112), .Z(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n786), .ZN(new_n1133));
  XOR2_X1   g0933(.A(new_n1133), .B(KEYINPUT113), .Z(new_n1134));
  AOI211_X1 g0934(.A(new_n1129), .B(new_n1134), .C1(new_n988), .C2(new_n769), .ZN(new_n1135));
  OR2_X1    g0935(.A1(new_n1029), .A2(KEYINPUT111), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1101), .B1(new_n1029), .B2(KEYINPUT111), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1135), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1110), .A2(new_n1138), .ZN(G390));
  INV_X1    g0939(.A(new_n753), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n474), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n657), .A2(new_n959), .A3(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n949), .B1(new_n753), .B2(new_n962), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  NOR3_X1   g0944(.A1(new_n753), .A2(new_n962), .A3(new_n949), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n704), .B(new_n962), .C1(new_n676), .C2(new_n695), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n1144), .A2(new_n1145), .B1(new_n1146), .B2(new_n950), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1145), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n951), .B1(new_n761), .B2(new_n962), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1148), .A2(new_n1150), .A3(new_n1143), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1147), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1142), .A2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n948), .B1(new_n1146), .B2(new_n950), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n930), .A2(new_n938), .B1(new_n1154), .B2(new_n931), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1149), .A2(new_n948), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n925), .A2(new_n928), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n933), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n937), .ZN(new_n1159));
  AND3_X1   g0959(.A1(new_n1156), .A2(new_n1159), .A3(new_n931), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1145), .B1(new_n1155), .B2(new_n1160), .ZN(new_n1161));
  AND3_X1   g0961(.A1(new_n936), .A2(KEYINPUT39), .A3(new_n937), .ZN(new_n1162));
  AOI21_X1  g0962(.A(KEYINPUT39), .B1(new_n1158), .B2(new_n937), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n1162), .A2(new_n1163), .B1(new_n932), .B2(new_n952), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1156), .A2(new_n1159), .A3(new_n931), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1164), .A2(new_n1165), .A3(new_n1148), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1161), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n728), .B1(new_n1153), .B2(new_n1167), .ZN(new_n1168));
  NOR3_X1   g0968(.A1(new_n1155), .A2(new_n1160), .A3(new_n1145), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1148), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1171), .A2(new_n1142), .A3(new_n1152), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1168), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1171), .A2(new_n1045), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n767), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n874), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n786), .B1(new_n261), .B2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1123), .B1(G116), .B2(new_n854), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT115), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n560), .A2(new_n802), .B1(new_n821), .B2(new_n816), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n303), .B1(new_n817), .B2(new_n790), .C1(new_n809), .C2(new_n509), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n815), .A2(new_n201), .B1(new_n796), .B2(new_n419), .ZN(new_n1182));
  NOR4_X1   g0982(.A1(new_n1179), .A2(new_n1180), .A3(new_n1181), .A4(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  OR2_X1    g0984(.A1(new_n1184), .A2(KEYINPUT116), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n303), .B1(new_n791), .B2(G125), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n272), .B2(new_n815), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(G128), .B2(new_n799), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n869), .A2(G150), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n1189), .A2(KEYINPUT53), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n1189), .A2(KEYINPUT53), .B1(G137), .B2(new_n801), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(KEYINPUT54), .B(G143), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n866), .A2(new_n811), .B1(new_n796), .B2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(G159), .B2(new_n1072), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1188), .A2(new_n1190), .A3(new_n1191), .A4(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1184), .A2(KEYINPUT116), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1185), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1177), .B1(new_n1197), .B2(new_n779), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1198), .B(KEYINPUT117), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1175), .A2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1173), .A2(new_n1174), .A3(new_n1200), .ZN(G378));
  AND3_X1   g1001(.A1(new_n963), .A2(new_n752), .A3(KEYINPUT101), .ZN(new_n1202));
  AOI21_X1  g1002(.A(KEYINPUT101), .B1(new_n963), .B2(new_n752), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(KEYINPUT40), .B1(new_n1204), .B2(new_n953), .ZN(new_n1205));
  OAI21_X1  g1005(.A(G330), .B1(new_n971), .B2(new_n972), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n277), .A2(new_n702), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n320), .A2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n314), .A2(new_n319), .A3(new_n1207), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1211), .A2(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1209), .A2(new_n1210), .A3(new_n1212), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  NOR3_X1   g1017(.A1(new_n1205), .A2(new_n1206), .A3(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n972), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n710), .B1(new_n1159), .B2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1216), .B1(new_n970), .B2(new_n1220), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n1218), .A2(new_n1221), .B1(new_n956), .B2(new_n957), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1217), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n939), .A2(new_n954), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(KEYINPUT100), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n939), .A2(new_n954), .A3(new_n955), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n970), .A2(new_n1220), .A3(new_n1216), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1223), .A2(new_n1225), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1222), .A2(new_n1228), .A3(new_n1045), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n787), .B1(new_n272), .B2(new_n874), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n815), .A2(new_n218), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n1075), .B(new_n1231), .C1(new_n492), .C2(new_n859), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n799), .A2(G116), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n297), .A2(G41), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n1234), .B1(new_n790), .B2(new_n816), .C1(new_n818), .C2(new_n201), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(G97), .B2(new_n801), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n811), .A2(new_n560), .ZN(new_n1237));
  XNOR2_X1  g1037(.A(new_n1237), .B(KEYINPUT118), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1232), .A2(new_n1233), .A3(new_n1236), .A4(new_n1238), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(new_n1239), .B(KEYINPUT58), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n809), .A2(new_n1192), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1241), .B(KEYINPUT119), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n859), .A2(G137), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n854), .A2(G128), .B1(new_n1072), .B2(G150), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(G125), .A2(new_n799), .B1(new_n801), .B2(G132), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .A4(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(KEYINPUT59), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n807), .A2(G159), .A3(new_n814), .ZN(new_n1248));
  AOI211_X1 g1048(.A(G33), .B(G41), .C1(new_n791), .C2(G124), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1247), .A2(new_n1248), .A3(new_n1249), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1246), .A2(KEYINPUT59), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n272), .B1(G33), .B2(G41), .ZN(new_n1252));
  OAI221_X1 g1052(.A(new_n1240), .B1(new_n1250), .B2(new_n1251), .C1(new_n1234), .C2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT120), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n779), .ZN(new_n1257));
  OAI221_X1 g1057(.A(new_n1230), .B1(new_n1255), .B2(new_n1257), .C1(new_n1216), .C2(new_n768), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1229), .A2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT121), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1229), .A2(KEYINPUT121), .A3(new_n1258), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT57), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n657), .A2(new_n959), .A3(new_n1141), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(new_n1171), .B2(new_n1152), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1222), .A2(new_n1228), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1264), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1152), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1142), .B1(new_n1167), .B2(new_n1269), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1270), .A2(KEYINPUT57), .A3(new_n1228), .A4(new_n1222), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1268), .A2(new_n727), .A3(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1263), .A2(new_n1272), .ZN(G375));
  XNOR2_X1  g1073(.A(new_n1265), .B(new_n1152), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1011), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  XOR2_X1   g1076(.A(new_n1276), .B(KEYINPUT122), .Z(new_n1277));
  NAND2_X1  g1077(.A1(new_n949), .A2(new_n767), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n786), .B1(G68), .B2(new_n1176), .ZN(new_n1279));
  AOI22_X1  g1079(.A1(new_n854), .A2(G137), .B1(new_n1072), .B2(G50), .ZN(new_n1280));
  OAI221_X1 g1080(.A(new_n1280), .B1(new_n264), .B2(new_n796), .C1(new_n823), .C2(new_n809), .ZN(new_n1281));
  AOI211_X1 g1081(.A(new_n303), .B(new_n1231), .C1(G128), .C2(new_n791), .ZN(new_n1282));
  OAI221_X1 g1082(.A(new_n1282), .B1(new_n866), .B2(new_n821), .C1(new_n802), .C2(new_n1192), .ZN(new_n1283));
  AOI211_X1 g1083(.A(new_n297), .B(new_n1047), .C1(G303), .C2(new_n791), .ZN(new_n1284));
  OAI221_X1 g1084(.A(new_n1284), .B1(new_n617), .B2(new_n802), .C1(new_n817), .C2(new_n821), .ZN(new_n1285));
  AOI22_X1  g1085(.A1(G107), .A2(new_n859), .B1(new_n854), .B2(G283), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n1286), .B(new_n1073), .C1(new_n419), .C2(new_n809), .ZN(new_n1287));
  OAI22_X1  g1087(.A1(new_n1281), .A2(new_n1283), .B1(new_n1285), .B2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1279), .B1(new_n1288), .B2(new_n779), .ZN(new_n1289));
  AOI22_X1  g1089(.A1(new_n1152), .A2(new_n1045), .B1(new_n1278), .B2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1277), .A2(new_n1290), .ZN(G381));
  OR4_X1    g1091(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1292));
  NOR4_X1   g1092(.A1(new_n1292), .A2(G381), .A3(G387), .A4(G378), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1293), .A2(new_n1272), .A3(new_n1263), .ZN(G407));
  NAND2_X1  g1094(.A1(new_n1174), .A2(new_n1200), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1295), .B1(new_n1172), .B2(new_n1168), .ZN(new_n1296));
  INV_X1    g1096(.A(G343), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(G213), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1296), .A2(new_n1299), .ZN(new_n1300));
  OAI211_X1 g1100(.A(G407), .B(G213), .C1(G375), .C2(new_n1300), .ZN(G409));
  XNOR2_X1  g1101(.A(G393), .B(new_n837), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(new_n1303));
  AND3_X1   g1103(.A1(new_n1046), .A2(new_n1068), .A3(G390), .ZN(new_n1304));
  AOI21_X1  g1104(.A(G390), .B1(new_n1046), .B2(new_n1068), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1303), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(G390), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(G387), .A2(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1046), .A2(new_n1068), .A3(G390), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1308), .A2(new_n1302), .A3(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT61), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1306), .A2(new_n1310), .A3(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1263), .A2(G378), .A3(new_n1272), .ZN(new_n1313));
  NOR3_X1   g1113(.A1(new_n1266), .A2(new_n1267), .A3(new_n1011), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1296), .B1(new_n1259), .B2(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1299), .B1(new_n1313), .B2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1269), .A2(new_n1265), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT60), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n728), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1319), .B1(new_n1274), .B2(new_n1318), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1320), .A2(G384), .A3(new_n1290), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(G384), .B1(new_n1320), .B2(new_n1290), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  AND2_X1   g1124(.A1(new_n1316), .A2(new_n1324), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1312), .B1(KEYINPUT63), .B2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1313), .A2(new_n1315), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1327), .A2(KEYINPUT123), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT123), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1313), .A2(new_n1329), .A3(new_n1315), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1328), .A2(new_n1298), .A3(new_n1324), .A4(new_n1330), .ZN(new_n1331));
  XOR2_X1   g1131(.A(KEYINPUT124), .B(KEYINPUT63), .Z(new_n1332));
  NAND2_X1  g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1299), .A2(G2897), .ZN(new_n1334));
  XNOR2_X1  g1134(.A(new_n1324), .B(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1335), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1328), .A2(new_n1298), .A3(new_n1330), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1326), .A2(new_n1333), .A3(new_n1338), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1311), .B1(new_n1335), .B2(new_n1316), .ZN(new_n1340));
  NAND4_X1  g1140(.A1(new_n1327), .A2(KEYINPUT62), .A3(new_n1298), .A4(new_n1324), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1341), .A2(KEYINPUT125), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT125), .ZN(new_n1343));
  NAND4_X1  g1143(.A1(new_n1316), .A2(new_n1343), .A3(KEYINPUT62), .A4(new_n1324), .ZN(new_n1344));
  AND2_X1   g1144(.A1(new_n1342), .A2(new_n1344), .ZN(new_n1345));
  INV_X1    g1145(.A(KEYINPUT62), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1331), .A2(new_n1346), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1340), .B1(new_n1345), .B2(new_n1347), .ZN(new_n1348));
  AND2_X1   g1148(.A1(new_n1306), .A2(new_n1310), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1339), .B1(new_n1348), .B2(new_n1349), .ZN(G405));
  OR2_X1    g1150(.A1(new_n1324), .A2(KEYINPUT126), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1324), .A2(KEYINPUT126), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(G375), .A2(new_n1296), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1353), .A2(new_n1313), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1351), .A2(new_n1352), .A3(new_n1354), .ZN(new_n1355));
  NAND4_X1  g1155(.A1(new_n1353), .A2(new_n1324), .A3(KEYINPUT126), .A4(new_n1313), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1355), .A2(new_n1356), .ZN(new_n1357));
  XNOR2_X1  g1157(.A(new_n1357), .B(new_n1349), .ZN(G402));
endmodule


