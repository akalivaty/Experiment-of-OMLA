//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 1 1 0 0 1 0 0 0 0 0 1 0 0 0 0 0 0 1 1 0 1 0 0 0 1 1 1 1 1 0 0 1 1 0 0 0 0 0 1 1 0 1 0 0 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n806, new_n807,
    new_n808, new_n810, new_n811, new_n812, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963, new_n964, new_n965;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT11), .B(G169gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT83), .B(KEYINPUT12), .ZN(new_n206));
  XOR2_X1   g005(.A(new_n205), .B(new_n206), .Z(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  XOR2_X1   g007(.A(G43gat), .B(G50gat), .Z(new_n209));
  INV_X1    g008(.A(G36gat), .ZN(new_n210));
  AND2_X1   g009(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G29gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n214), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n209), .B1(new_n216), .B2(KEYINPUT15), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n217), .B1(KEYINPUT15), .B2(new_n216), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n216), .A2(KEYINPUT15), .A3(new_n209), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n218), .A2(KEYINPUT17), .A3(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT86), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n218), .A2(KEYINPUT86), .A3(KEYINPUT17), .A4(new_n219), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(G15gat), .B(G22gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT16), .ZN(new_n226));
  AOI21_X1  g025(.A(G1gat), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT84), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n225), .B(new_n228), .C1(new_n226), .C2(G1gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n232), .B1(KEYINPUT85), .B2(G8gat), .ZN(new_n233));
  XNOR2_X1  g032(.A(KEYINPUT85), .B(G8gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n230), .A2(new_n231), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(KEYINPUT17), .B1(new_n218), .B2(new_n219), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n224), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(G229gat), .A2(G233gat), .ZN(new_n240));
  AOI22_X1  g039(.A1(new_n233), .A2(new_n235), .B1(new_n218), .B2(new_n219), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT87), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n243), .A2(KEYINPUT18), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n239), .A2(new_n240), .A3(new_n242), .A4(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n218), .A2(new_n219), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n236), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(KEYINPUT88), .B(KEYINPUT13), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(new_n240), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n246), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n241), .B1(new_n224), .B2(new_n238), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n245), .B1(new_n253), .B2(new_n240), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n208), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n253), .A2(new_n240), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(new_n244), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n257), .A2(new_n207), .A3(new_n251), .A4(new_n246), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(G169gat), .ZN(new_n261));
  INV_X1    g060(.A(G176gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(G169gat), .A2(G176gat), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  OAI211_X1 g064(.A(KEYINPUT69), .B(new_n263), .C1(new_n265), .C2(KEYINPUT26), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n268));
  NOR2_X1   g067(.A1(G169gat), .A2(G176gat), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n266), .B(new_n270), .C1(KEYINPUT26), .C2(new_n263), .ZN(new_n271));
  NAND2_X1  g070(.A1(G183gat), .A2(G190gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT27), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(G183gat), .ZN(new_n275));
  INV_X1    g074(.A(G183gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT27), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT67), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(G190gat), .B1(new_n275), .B2(KEYINPUT67), .ZN(new_n281));
  AOI21_X1  g080(.A(KEYINPUT28), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT28), .ZN(new_n283));
  NOR3_X1   g082(.A1(new_n278), .A2(new_n283), .A3(G190gat), .ZN(new_n284));
  OAI21_X1  g083(.A(KEYINPUT68), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(KEYINPUT27), .B(G183gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n286), .A2(KEYINPUT67), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n275), .A2(KEYINPUT67), .ZN(new_n288));
  INV_X1    g087(.A(G190gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n283), .B1(new_n287), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n284), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT68), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n273), .B1(new_n285), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT24), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n276), .A2(G190gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n289), .A2(G183gat), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n272), .A2(KEYINPUT24), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n269), .A2(KEYINPUT23), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT23), .ZN(new_n304));
  NOR3_X1   g103(.A1(new_n304), .A2(G169gat), .A3(G176gat), .ZN(new_n305));
  NOR3_X1   g104(.A1(new_n303), .A2(new_n305), .A3(new_n265), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT25), .B1(new_n302), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT25), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n309), .B1(new_n263), .B2(new_n304), .ZN(new_n310));
  INV_X1    g109(.A(new_n301), .ZN(new_n311));
  XNOR2_X1  g110(.A(G183gat), .B(G190gat), .ZN(new_n312));
  OAI211_X1 g111(.A(new_n310), .B(new_n311), .C1(new_n297), .C2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT64), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n314), .B1(new_n305), .B2(new_n265), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n261), .A2(new_n262), .A3(KEYINPUT23), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n316), .A2(KEYINPUT64), .A3(new_n264), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NOR3_X1   g117(.A1(new_n313), .A2(new_n318), .A3(KEYINPUT65), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT65), .ZN(new_n320));
  AND3_X1   g119(.A1(new_n316), .A2(KEYINPUT64), .A3(new_n264), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT64), .B1(new_n316), .B2(new_n264), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(KEYINPUT25), .B1(new_n269), .B2(KEYINPUT23), .ZN(new_n324));
  NOR3_X1   g123(.A1(new_n300), .A2(new_n324), .A3(new_n301), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n320), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n308), .B1(new_n319), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n296), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G226gat), .ZN(new_n329));
  INV_X1    g128(.A(G233gat), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n331), .A2(KEYINPUT29), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT66), .ZN(new_n334));
  OAI21_X1  g133(.A(KEYINPUT65), .B1(new_n313), .B2(new_n318), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n323), .A2(new_n325), .A3(new_n320), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n334), .B1(new_n337), .B2(new_n308), .ZN(new_n338));
  AOI211_X1 g137(.A(KEYINPUT66), .B(new_n307), .C1(new_n335), .C2(new_n336), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n331), .B(new_n296), .C1(new_n338), .C2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n333), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(G197gat), .B(G204gat), .ZN(new_n342));
  INV_X1    g141(.A(G211gat), .ZN(new_n343));
  INV_X1    g142(.A(G218gat), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n342), .B1(KEYINPUT22), .B2(new_n345), .ZN(new_n346));
  XOR2_X1   g145(.A(G211gat), .B(G218gat), .Z(new_n347));
  OR2_X1    g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n346), .A2(new_n347), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n341), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n350), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n307), .B1(new_n335), .B2(new_n336), .ZN(new_n353));
  INV_X1    g152(.A(new_n331), .ZN(new_n354));
  NOR3_X1   g153(.A1(new_n295), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n327), .A2(KEYINPUT66), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n353), .A2(new_n334), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n295), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n332), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n352), .B(new_n356), .C1(new_n359), .C2(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(G8gat), .B(G36gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(G64gat), .B(G92gat), .ZN(new_n363));
  XOR2_X1   g162(.A(new_n362), .B(new_n363), .Z(new_n364));
  NAND3_X1  g163(.A1(new_n351), .A2(new_n361), .A3(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT30), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n351), .A2(KEYINPUT30), .A3(new_n361), .A4(new_n364), .ZN(new_n368));
  INV_X1    g167(.A(new_n364), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n296), .B1(new_n338), .B2(new_n339), .ZN(new_n370));
  AOI211_X1 g169(.A(new_n350), .B(new_n355), .C1(new_n370), .C2(new_n332), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n352), .B1(new_n333), .B2(new_n340), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n369), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n367), .A2(KEYINPUT76), .A3(new_n368), .A4(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n371), .A2(new_n372), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT76), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n375), .A2(new_n376), .A3(KEYINPUT30), .A4(new_n364), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  XOR2_X1   g177(.A(G141gat), .B(G148gat), .Z(new_n379));
  INV_X1    g178(.A(G155gat), .ZN(new_n380));
  INV_X1    g179(.A(G162gat), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT2), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT77), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT2), .ZN(new_n385));
  AOI22_X1  g184(.A1(new_n384), .A2(new_n385), .B1(G155gat), .B2(G162gat), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n383), .B(new_n386), .C1(G155gat), .C2(G162gat), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n386), .B1(G155gat), .B2(G162gat), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n388), .A2(new_n382), .A3(new_n379), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(KEYINPUT3), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT3), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n387), .A2(new_n392), .A3(new_n389), .ZN(new_n393));
  INV_X1    g192(.A(G113gat), .ZN(new_n394));
  INV_X1    g193(.A(G120gat), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT1), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(G127gat), .B(G134gat), .ZN(new_n397));
  XOR2_X1   g196(.A(KEYINPUT70), .B(G113gat), .Z(new_n398));
  OAI211_X1 g197(.A(new_n396), .B(new_n397), .C1(new_n398), .C2(new_n395), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n396), .B1(new_n394), .B2(new_n395), .ZN(new_n400));
  INV_X1    g199(.A(new_n397), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n391), .A2(new_n393), .A3(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n390), .ZN(new_n405));
  INV_X1    g204(.A(new_n403), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n405), .A2(KEYINPUT4), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(G225gat), .A2(G233gat), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n387), .A2(new_n389), .A3(new_n402), .A4(new_n399), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT4), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n404), .A2(new_n407), .A3(new_n408), .A4(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n408), .ZN(new_n413));
  INV_X1    g212(.A(new_n409), .ZN(new_n414));
  AOI22_X1  g213(.A1(new_n387), .A2(new_n389), .B1(new_n402), .B2(new_n399), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT5), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n412), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n409), .B(KEYINPUT4), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n419), .A2(KEYINPUT5), .A3(new_n408), .A4(new_n404), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  XNOR2_X1  g220(.A(G1gat), .B(G29gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n422), .B(KEYINPUT0), .ZN(new_n423));
  XNOR2_X1  g222(.A(G57gat), .B(G85gat), .ZN(new_n424));
  XOR2_X1   g223(.A(new_n423), .B(new_n424), .Z(new_n425));
  NAND2_X1  g224(.A1(new_n421), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT6), .ZN(new_n427));
  INV_X1    g226(.A(new_n425), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n418), .A2(new_n428), .A3(new_n420), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n426), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n418), .A2(KEYINPUT6), .A3(new_n420), .A4(new_n428), .ZN(new_n431));
  AND2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n378), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT29), .ZN(new_n435));
  AOI21_X1  g234(.A(KEYINPUT3), .B1(new_n350), .B2(new_n435), .ZN(new_n436));
  OAI211_X1 g235(.A(G228gat), .B(G233gat), .C1(new_n436), .C2(new_n405), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n350), .B1(new_n393), .B2(new_n435), .ZN(new_n438));
  OR2_X1    g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(G22gat), .ZN(new_n440));
  NAND2_X1  g239(.A1(G228gat), .A2(G233gat), .ZN(new_n441));
  XOR2_X1   g240(.A(new_n441), .B(KEYINPUT79), .Z(new_n442));
  NAND3_X1  g241(.A1(new_n346), .A2(KEYINPUT80), .A3(new_n347), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n435), .B(new_n443), .C1(new_n350), .C2(KEYINPUT80), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n405), .B1(new_n444), .B2(new_n392), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n442), .B1(new_n445), .B2(new_n438), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n439), .A2(new_n440), .A3(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n440), .B1(new_n439), .B2(new_n446), .ZN(new_n449));
  OAI21_X1  g248(.A(KEYINPUT81), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n439), .A2(new_n446), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(G22gat), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT81), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n452), .A2(new_n447), .A3(new_n453), .ZN(new_n454));
  XOR2_X1   g253(.A(G78gat), .B(G106gat), .Z(new_n455));
  XNOR2_X1  g254(.A(new_n455), .B(KEYINPUT78), .ZN(new_n456));
  XOR2_X1   g255(.A(KEYINPUT31), .B(G50gat), .Z(new_n457));
  XNOR2_X1  g256(.A(new_n456), .B(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n450), .A2(new_n454), .A3(new_n459), .ZN(new_n460));
  OAI211_X1 g259(.A(KEYINPUT81), .B(new_n458), .C1(new_n448), .C2(new_n449), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NOR3_X1   g261(.A1(new_n434), .A2(KEYINPUT35), .A3(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT74), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT32), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n406), .B(new_n296), .C1(new_n338), .C2(new_n339), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT71), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n357), .A2(new_n358), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT71), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n468), .A2(new_n469), .A3(new_n406), .A4(new_n296), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n370), .A2(new_n403), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n467), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(G227gat), .A2(G233gat), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n465), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(KEYINPUT33), .B1(new_n472), .B2(new_n474), .ZN(new_n476));
  XNOR2_X1  g275(.A(G15gat), .B(G43gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n477), .B(KEYINPUT72), .ZN(new_n478));
  XNOR2_X1  g277(.A(G71gat), .B(G99gat), .ZN(new_n479));
  XOR2_X1   g278(.A(new_n478), .B(new_n479), .Z(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  NOR3_X1   g280(.A1(new_n475), .A2(new_n476), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n472), .A2(new_n474), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT33), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n483), .A2(KEYINPUT32), .A3(new_n486), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n467), .A2(new_n470), .A3(new_n471), .A4(new_n473), .ZN(new_n488));
  XNOR2_X1  g287(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OR2_X1    g289(.A1(new_n488), .A2(KEYINPUT34), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n487), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n464), .B1(new_n482), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n490), .B1(KEYINPUT34), .B2(new_n488), .ZN(new_n494));
  AOI211_X1 g293(.A(new_n465), .B(new_n485), .C1(new_n472), .C2(new_n474), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n475), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n483), .A2(new_n484), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n497), .A2(new_n498), .A3(new_n480), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n496), .A2(KEYINPUT74), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n493), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT75), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n502), .B(new_n494), .C1(new_n482), .C2(new_n495), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n494), .B1(new_n482), .B2(new_n495), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT75), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n463), .A2(new_n501), .A3(new_n503), .A4(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n432), .B1(new_n374), .B2(new_n377), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n460), .A2(new_n461), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n501), .A2(new_n507), .A3(new_n504), .A4(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT35), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  NOR3_X1   g310(.A1(new_n482), .A2(new_n492), .A3(new_n464), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT74), .B1(new_n496), .B2(new_n499), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n504), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT36), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n507), .A2(new_n508), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT40), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n404), .A2(new_n411), .A3(new_n407), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT39), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n518), .A2(new_n519), .A3(new_n413), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(new_n425), .ZN(new_n521));
  INV_X1    g320(.A(new_n415), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n522), .A2(new_n408), .A3(new_n409), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT39), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n524), .B1(new_n518), .B2(new_n413), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n517), .B1(new_n521), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n518), .A2(new_n413), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n527), .A2(KEYINPUT39), .A3(new_n523), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n528), .A2(KEYINPUT40), .A3(new_n425), .A4(new_n520), .ZN(new_n529));
  AND3_X1   g328(.A1(new_n526), .A2(new_n529), .A3(new_n429), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n368), .A2(new_n373), .A3(KEYINPUT76), .ZN(new_n531));
  AOI21_X1  g330(.A(KEYINPUT30), .B1(new_n375), .B2(new_n364), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n377), .B(new_n530), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT82), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n374), .A2(KEYINPUT82), .A3(new_n377), .A4(new_n530), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n430), .A2(new_n431), .A3(new_n365), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n351), .A2(new_n361), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n369), .B1(new_n539), .B2(KEYINPUT37), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT37), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n355), .B1(new_n370), .B2(new_n332), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n542), .B1(new_n543), .B2(new_n350), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n341), .A2(new_n352), .ZN(new_n545));
  AOI21_X1  g344(.A(KEYINPUT38), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n538), .B1(new_n541), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n375), .A2(new_n542), .ZN(new_n548));
  OAI21_X1  g347(.A(KEYINPUT38), .B1(new_n540), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n462), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n516), .B1(new_n537), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT36), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n501), .A2(new_n505), .A3(new_n503), .A4(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n515), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n260), .B1(new_n511), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(G85gat), .A2(G92gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(KEYINPUT7), .ZN(new_n557));
  NOR2_X1   g356(.A1(G85gat), .A2(G92gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(G99gat), .A2(G106gat), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n558), .B1(KEYINPUT8), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(G99gat), .B(G106gat), .Z(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n562), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n564), .A2(new_n557), .A3(new_n560), .ZN(new_n565));
  AND2_X1   g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n237), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n224), .A2(new_n567), .ZN(new_n568));
  AND2_X1   g367(.A1(G232gat), .A2(G233gat), .ZN(new_n569));
  AOI22_X1  g368(.A1(new_n247), .A2(new_n566), .B1(KEYINPUT41), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(G190gat), .B(G218gat), .Z(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n569), .A2(KEYINPUT41), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT92), .ZN(new_n575));
  XNOR2_X1  g374(.A(G134gat), .B(G162gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  OR2_X1    g377(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n573), .A2(new_n578), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT9), .ZN(new_n581));
  INV_X1    g380(.A(G71gat), .ZN(new_n582));
  INV_X1    g381(.A(G78gat), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(KEYINPUT89), .ZN(new_n585));
  XOR2_X1   g384(.A(G57gat), .B(G64gat), .Z(new_n586));
  INV_X1    g385(.A(KEYINPUT89), .ZN(new_n587));
  OAI211_X1 g386(.A(new_n587), .B(new_n581), .C1(new_n582), .C2(new_n583), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n585), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(G71gat), .B(G78gat), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n585), .A2(new_n586), .A3(new_n590), .A4(new_n588), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT21), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  XOR2_X1   g395(.A(KEYINPUT91), .B(KEYINPUT19), .Z(new_n597));
  XOR2_X1   g396(.A(new_n596), .B(new_n597), .Z(new_n598));
  OAI211_X1 g397(.A(new_n233), .B(new_n235), .C1(new_n595), .C2(new_n594), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G127gat), .B(G155gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT20), .ZN(new_n602));
  NAND2_X1  g401(.A1(G231gat), .A2(G233gat), .ZN(new_n603));
  XOR2_X1   g402(.A(new_n603), .B(KEYINPUT90), .Z(new_n604));
  XNOR2_X1  g403(.A(new_n602), .B(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G183gat), .B(G211gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n600), .B(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n563), .A2(new_n565), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT10), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n592), .A2(new_n563), .A3(new_n593), .A4(new_n565), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n566), .A2(KEYINPUT10), .A3(new_n592), .A4(new_n593), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(KEYINPUT93), .ZN(new_n616));
  NAND2_X1  g415(.A1(G230gat), .A2(G233gat), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT93), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n613), .A2(new_n618), .A3(new_n614), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n616), .A2(new_n617), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n610), .A2(new_n612), .ZN(new_n621));
  INV_X1    g420(.A(new_n617), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G120gat), .B(G148gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(G176gat), .B(G204gat), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n624), .B(new_n625), .Z(new_n626));
  NAND3_X1  g425(.A1(new_n620), .A2(new_n623), .A3(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n615), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n623), .B1(new_n628), .B2(new_n622), .ZN(new_n629));
  INV_X1    g428(.A(new_n626), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n579), .A2(new_n580), .A3(new_n608), .A4(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n555), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(new_n432), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(G1gat), .ZN(G1324gat));
  INV_X1    g438(.A(new_n378), .ZN(new_n640));
  XOR2_X1   g439(.A(KEYINPUT16), .B(G8gat), .Z(new_n641));
  NAND3_X1  g440(.A1(new_n637), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  AND3_X1   g441(.A1(new_n642), .A2(KEYINPUT94), .A3(KEYINPUT42), .ZN(new_n643));
  AOI21_X1  g442(.A(KEYINPUT42), .B1(new_n642), .B2(KEYINPUT94), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n637), .A2(new_n640), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT95), .ZN(new_n646));
  AND3_X1   g445(.A1(new_n645), .A2(new_n646), .A3(G8gat), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n646), .B1(new_n645), .B2(G8gat), .ZN(new_n648));
  OAI22_X1  g447(.A1(new_n643), .A2(new_n644), .B1(new_n647), .B2(new_n648), .ZN(G1325gat));
  NAND2_X1  g448(.A1(new_n515), .A2(new_n553), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(G15gat), .B1(new_n636), .B2(new_n651), .ZN(new_n652));
  AND3_X1   g451(.A1(new_n501), .A2(new_n503), .A3(new_n505), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n654), .A2(G15gat), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n652), .B1(new_n636), .B2(new_n655), .ZN(G1326gat));
  NOR2_X1   g455(.A1(new_n636), .A2(new_n508), .ZN(new_n657));
  XOR2_X1   g456(.A(KEYINPUT43), .B(G22gat), .Z(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(G1327gat));
  AND2_X1   g458(.A1(new_n579), .A2(new_n580), .ZN(new_n660));
  INV_X1    g459(.A(new_n608), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(new_n633), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n555), .A2(new_n214), .A3(new_n432), .A4(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT45), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n579), .A2(new_n580), .ZN(new_n666));
  AND2_X1   g465(.A1(new_n666), .A2(KEYINPUT44), .ZN(new_n667));
  AND3_X1   g466(.A1(new_n515), .A2(new_n551), .A3(new_n553), .ZN(new_n668));
  AOI22_X1  g467(.A1(new_n653), .A2(new_n463), .B1(new_n509), .B2(KEYINPUT35), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n246), .A2(new_n251), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n207), .B1(new_n671), .B2(new_n257), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n252), .A2(new_n254), .A3(new_n208), .ZN(new_n673));
  OAI21_X1  g472(.A(KEYINPUT96), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT96), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n255), .A2(new_n258), .A3(new_n675), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n678), .A2(new_n662), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT97), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n434), .A2(new_n680), .A3(new_n462), .ZN(new_n681));
  OAI21_X1  g480(.A(KEYINPUT97), .B1(new_n507), .B2(new_n508), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n537), .A2(new_n550), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n515), .A2(new_n683), .A3(new_n553), .A4(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n660), .B1(new_n511), .B2(new_n685), .ZN(new_n686));
  OAI211_X1 g485(.A(new_n670), .B(new_n679), .C1(new_n686), .C2(KEYINPUT44), .ZN(new_n687));
  OAI21_X1  g486(.A(G29gat), .B1(new_n687), .B2(new_n433), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n665), .A2(new_n688), .ZN(G1328gat));
  NAND2_X1  g488(.A1(new_n555), .A2(new_n663), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n690), .A2(G36gat), .A3(new_n378), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT46), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n687), .A2(KEYINPUT98), .A3(new_n378), .ZN(new_n693));
  OAI21_X1  g492(.A(KEYINPUT98), .B1(new_n687), .B2(new_n378), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(G36gat), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n692), .B1(new_n693), .B2(new_n695), .ZN(G1329gat));
  NOR2_X1   g495(.A1(new_n690), .A2(new_n654), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n650), .A2(G43gat), .ZN(new_n698));
  OAI22_X1  g497(.A1(new_n697), .A2(G43gat), .B1(new_n687), .B2(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g499(.A(G50gat), .B1(new_n687), .B2(new_n508), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(KEYINPUT99), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n508), .A2(G50gat), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n555), .A2(new_n663), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT48), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n702), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  OAI211_X1 g506(.A(new_n701), .B(new_n704), .C1(KEYINPUT99), .C2(KEYINPUT48), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(G1331gat));
  NOR4_X1   g508(.A1(new_n677), .A2(new_n661), .A3(new_n666), .A4(new_n633), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT100), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n711), .B1(new_n511), .B2(new_n685), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(new_n432), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g513(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n712), .A2(new_n640), .A3(new_n715), .ZN(new_n716));
  OR2_X1    g515(.A1(new_n716), .A2(KEYINPUT101), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(KEYINPUT101), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n717), .A2(new_n720), .A3(new_n718), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(G1333gat));
  NAND3_X1  g523(.A1(new_n712), .A2(new_n582), .A3(new_n653), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n712), .A2(new_n650), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n725), .B1(new_n726), .B2(new_n582), .ZN(new_n727));
  XOR2_X1   g526(.A(KEYINPUT102), .B(KEYINPUT50), .Z(new_n728));
  XNOR2_X1  g527(.A(new_n727), .B(new_n728), .ZN(G1334gat));
  NAND2_X1  g528(.A1(new_n712), .A2(new_n462), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g530(.A1(new_n677), .A2(new_n608), .A3(new_n633), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n670), .B(new_n732), .C1(new_n686), .C2(KEYINPUT44), .ZN(new_n733));
  OAI21_X1  g532(.A(G85gat), .B1(new_n733), .B2(new_n433), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n433), .A2(G85gat), .A3(new_n633), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n677), .A2(new_n608), .ZN(new_n736));
  AND3_X1   g535(.A1(new_n686), .A2(KEYINPUT51), .A3(new_n736), .ZN(new_n737));
  AOI21_X1  g536(.A(KEYINPUT51), .B1(new_n686), .B2(new_n736), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n735), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n734), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(KEYINPUT103), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT103), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n734), .A2(new_n739), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n741), .A2(new_n743), .ZN(G1336gat));
  NOR2_X1   g543(.A1(new_n633), .A2(G92gat), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n640), .B(new_n745), .C1(new_n737), .C2(new_n738), .ZN(new_n746));
  OAI21_X1  g545(.A(G92gat), .B1(new_n733), .B2(new_n378), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(KEYINPUT52), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT52), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n746), .A2(new_n747), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n751), .ZN(G1337gat));
  OAI21_X1  g551(.A(G99gat), .B1(new_n733), .B2(new_n651), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n654), .A2(G99gat), .A3(new_n633), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n737), .B2(new_n738), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n755), .ZN(G1338gat));
  OAI21_X1  g555(.A(G106gat), .B1(new_n733), .B2(new_n508), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n508), .A2(G106gat), .A3(new_n633), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n758), .B1(new_n737), .B2(new_n738), .ZN(new_n759));
  XNOR2_X1  g558(.A(KEYINPUT104), .B(KEYINPUT53), .ZN(new_n760));
  AND3_X1   g559(.A1(new_n757), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n760), .B1(new_n757), .B2(new_n759), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n761), .A2(new_n762), .ZN(G1339gat));
  INV_X1    g562(.A(KEYINPUT105), .ZN(new_n764));
  AOI211_X1 g563(.A(KEYINPUT54), .B(new_n622), .C1(new_n613), .C2(new_n614), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n764), .B1(new_n765), .B2(new_n626), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT54), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n615), .A2(new_n767), .A3(new_n617), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n768), .A2(KEYINPUT105), .A3(new_n630), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n767), .B1(new_n628), .B2(new_n622), .ZN(new_n770));
  AOI22_X1  g569(.A1(new_n766), .A2(new_n769), .B1(new_n620), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n627), .B1(new_n771), .B2(KEYINPUT55), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n766), .A2(new_n769), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n620), .A2(new_n770), .ZN(new_n774));
  AND3_X1   g573(.A1(new_n773), .A2(KEYINPUT55), .A3(new_n774), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n674), .A2(new_n776), .A3(new_n676), .ZN(new_n777));
  OAI22_X1  g576(.A1(new_n253), .A2(new_n240), .B1(new_n248), .B2(new_n250), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n778), .A2(new_n205), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n673), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(new_n632), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n666), .B1(new_n777), .B2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n666), .A2(new_n780), .A3(new_n776), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n661), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n677), .A2(new_n634), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n432), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n501), .A2(new_n504), .A3(new_n508), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n789), .A2(new_n640), .A3(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n791), .A2(new_n398), .A3(new_n677), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n640), .A2(new_n433), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n654), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n462), .B1(new_n785), .B2(new_n787), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(G113gat), .B1(new_n797), .B2(new_n260), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n792), .A2(new_n798), .ZN(G1340gat));
  NAND3_X1  g598(.A1(new_n791), .A2(new_n395), .A3(new_n632), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n795), .A2(new_n632), .A3(new_n796), .ZN(new_n801));
  AND3_X1   g600(.A1(new_n801), .A2(KEYINPUT106), .A3(G120gat), .ZN(new_n802));
  AOI21_X1  g601(.A(KEYINPUT106), .B1(new_n801), .B2(G120gat), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n800), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  XOR2_X1   g603(.A(new_n804), .B(KEYINPUT107), .Z(G1341gat));
  INV_X1    g604(.A(G127gat), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n791), .A2(new_n806), .A3(new_n608), .ZN(new_n807));
  OAI21_X1  g606(.A(G127gat), .B1(new_n797), .B2(new_n661), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(G1342gat));
  INV_X1    g608(.A(G134gat), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n791), .A2(new_n810), .A3(new_n666), .ZN(new_n811));
  OR2_X1    g610(.A1(new_n811), .A2(KEYINPUT56), .ZN(new_n812));
  OAI21_X1  g611(.A(G134gat), .B1(new_n797), .B2(new_n660), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(KEYINPUT56), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(G1343gat));
  INV_X1    g614(.A(KEYINPUT108), .ZN(new_n816));
  AOI22_X1  g615(.A1(new_n776), .A2(new_n259), .B1(new_n780), .B2(new_n632), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n783), .B1(new_n817), .B2(new_n666), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n786), .B1(new_n818), .B2(new_n661), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n462), .A2(KEYINPUT57), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n816), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n820), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n773), .A2(new_n774), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT55), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n771), .A2(KEYINPUT55), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n825), .A2(new_n627), .A3(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n781), .B1(new_n260), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n660), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n608), .B1(new_n829), .B2(new_n783), .ZN(new_n830));
  OAI211_X1 g629(.A(KEYINPUT108), .B(new_n822), .C1(new_n830), .C2(new_n786), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n508), .B1(new_n785), .B2(new_n787), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n821), .B(new_n831), .C1(new_n832), .C2(KEYINPUT57), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n650), .A2(new_n794), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n677), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n836), .A2(KEYINPUT58), .A3(G141gat), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n789), .A2(KEYINPUT109), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n378), .A2(new_n462), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n650), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n433), .B1(new_n785), .B2(new_n787), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT109), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AND3_X1   g642(.A1(new_n838), .A2(new_n840), .A3(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(G141gat), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n844), .A2(new_n845), .A3(new_n259), .ZN(new_n846));
  OR2_X1    g645(.A1(KEYINPUT110), .A2(KEYINPUT58), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n833), .A2(new_n259), .A3(new_n834), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(G141gat), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n850), .B1(new_n846), .B2(KEYINPUT110), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT58), .ZN(new_n852));
  AOI22_X1  g651(.A1(new_n837), .A2(new_n848), .B1(new_n851), .B2(new_n852), .ZN(G1344gat));
  INV_X1    g652(.A(G148gat), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n844), .A2(new_n854), .A3(new_n632), .ZN(new_n855));
  AOI211_X1 g654(.A(KEYINPUT59), .B(new_n854), .C1(new_n835), .C2(new_n632), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT59), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n818), .A2(new_n661), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n635), .A2(new_n260), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n858), .B1(new_n861), .B2(new_n508), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n820), .B1(new_n785), .B2(new_n787), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n865), .A2(new_n632), .A3(new_n834), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n857), .B1(new_n866), .B2(G148gat), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n855), .B1(new_n856), .B2(new_n867), .ZN(G1345gat));
  NAND3_X1  g667(.A1(new_n844), .A2(new_n380), .A3(new_n608), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n835), .A2(new_n608), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n869), .B1(new_n870), .B2(new_n380), .ZN(G1346gat));
  NAND2_X1  g670(.A1(new_n821), .A2(new_n831), .ZN(new_n872));
  AOI21_X1  g671(.A(KEYINPUT57), .B1(new_n788), .B2(new_n462), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n666), .B(new_n834), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(KEYINPUT112), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT112), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n833), .A2(new_n876), .A3(new_n666), .A4(new_n834), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n875), .A2(G162gat), .A3(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n660), .A2(G162gat), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n838), .A2(new_n840), .A3(new_n843), .A4(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT111), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI211_X1 g681(.A(new_n839), .B(new_n650), .C1(new_n841), .C2(new_n842), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n883), .A2(KEYINPUT111), .A3(new_n838), .A4(new_n879), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n878), .A2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT113), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n878), .A2(new_n885), .A3(KEYINPUT113), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(G1347gat));
  NOR2_X1   g689(.A1(new_n790), .A2(new_n378), .ZN(new_n891));
  OR2_X1    g690(.A1(new_n891), .A2(KEYINPUT114), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n432), .B1(new_n785), .B2(new_n787), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n891), .A2(KEYINPUT114), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(KEYINPUT115), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT115), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n892), .A2(new_n897), .A3(new_n893), .A4(new_n894), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n899), .A2(new_n261), .A3(new_n677), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n640), .A2(new_n433), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n654), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n796), .ZN(new_n903));
  OAI21_X1  g702(.A(G169gat), .B1(new_n903), .B2(new_n260), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n904), .B(KEYINPUT116), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n900), .A2(new_n905), .ZN(G1348gat));
  NAND3_X1  g705(.A1(new_n899), .A2(new_n262), .A3(new_n632), .ZN(new_n907));
  OAI21_X1  g706(.A(G176gat), .B1(new_n903), .B2(new_n633), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(G1349gat));
  OAI21_X1  g708(.A(G183gat), .B1(new_n903), .B2(new_n661), .ZN(new_n910));
  XNOR2_X1  g709(.A(KEYINPUT117), .B(KEYINPUT60), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n608), .A2(new_n286), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n910), .B(new_n911), .C1(new_n895), .C2(new_n912), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n913), .A2(KEYINPUT118), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n913), .A2(KEYINPUT118), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n910), .B1(new_n895), .B2(new_n912), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(KEYINPUT60), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n914), .B1(new_n915), .B2(new_n917), .ZN(G1350gat));
  NAND4_X1  g717(.A1(new_n896), .A2(new_n289), .A3(new_n666), .A4(new_n898), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT61), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n902), .A2(new_n666), .A3(new_n796), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n920), .B1(new_n921), .B2(G190gat), .ZN(new_n922));
  AND3_X1   g721(.A1(new_n921), .A2(new_n920), .A3(G190gat), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n919), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT119), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OAI211_X1 g725(.A(new_n919), .B(KEYINPUT119), .C1(new_n922), .C2(new_n923), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(G1351gat));
  NOR2_X1   g727(.A1(new_n650), .A2(new_n901), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(new_n832), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n930), .A2(G197gat), .A3(new_n678), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT120), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n862), .A2(new_n932), .A3(new_n864), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n929), .A2(KEYINPUT121), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT121), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n935), .B1(new_n650), .B2(new_n901), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n859), .A2(new_n860), .ZN(new_n938));
  AOI21_X1  g737(.A(KEYINPUT57), .B1(new_n938), .B2(new_n462), .ZN(new_n939));
  OAI21_X1  g738(.A(KEYINPUT120), .B1(new_n939), .B2(new_n863), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n933), .A2(new_n937), .A3(new_n940), .A4(new_n259), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n931), .B1(new_n941), .B2(G197gat), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n942), .B(KEYINPUT122), .ZN(G1352gat));
  XNOR2_X1  g742(.A(KEYINPUT123), .B(G204gat), .ZN(new_n944));
  NAND4_X1  g743(.A1(new_n933), .A2(new_n937), .A3(new_n940), .A4(new_n632), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT125), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n947), .B1(new_n946), .B2(new_n945), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT62), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n944), .B1(KEYINPUT124), .B2(new_n949), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n930), .A2(new_n633), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(KEYINPUT124), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n951), .B(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n948), .A2(new_n953), .ZN(G1353gat));
  AOI21_X1  g753(.A(new_n661), .B1(new_n862), .B2(new_n864), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n343), .B1(new_n955), .B2(new_n937), .ZN(new_n956));
  OR3_X1    g755(.A1(new_n956), .A2(KEYINPUT126), .A3(KEYINPUT63), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n929), .A2(new_n343), .A3(new_n608), .A4(new_n832), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n956), .A2(KEYINPUT63), .ZN(new_n959));
  OAI21_X1  g758(.A(KEYINPUT126), .B1(new_n956), .B2(KEYINPUT63), .ZN(new_n960));
  OAI211_X1 g759(.A(new_n957), .B(new_n958), .C1(new_n959), .C2(new_n960), .ZN(G1354gat));
  NOR2_X1   g760(.A1(new_n660), .A2(new_n344), .ZN(new_n962));
  NAND4_X1  g761(.A1(new_n933), .A2(new_n937), .A3(new_n940), .A4(new_n962), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n344), .B1(new_n930), .B2(new_n660), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n965), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


