//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 0 1 0 1 0 1 1 1 0 1 1 0 0 0 0 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0 1 0 1 0 1 1 0 0 1 0 1 1 0 0 0 1 0 1 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:31 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n570,
    new_n572, new_n573, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n592, new_n593, new_n594, new_n597,
    new_n598, new_n599, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n636, new_n639,
    new_n640, new_n642, new_n643, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1167, new_n1168, new_n1169;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT64), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n452), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(new_n453), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  AOI22_X1  g042(.A1(new_n467), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  OR2_X1    g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(G101), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n464), .A2(new_n466), .ZN(new_n472));
  INV_X1    g047(.A(G137), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(new_n469), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  NOR2_X1   g052(.A1(new_n472), .A2(new_n469), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n472), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n469), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  OAI21_X1  g060(.A(G2104), .B1(new_n469), .B2(G114), .ZN(new_n486));
  INV_X1    g061(.A(G102), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n486), .B1(new_n487), .B2(new_n469), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n467), .A2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G126), .ZN(new_n490));
  OAI21_X1  g065(.A(KEYINPUT65), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT65), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n478), .A2(new_n492), .A3(G126), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n488), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n480), .A2(G138), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n480), .A2(new_n497), .A3(G138), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n494), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  XNOR2_X1  g076(.A(KEYINPUT5), .B(G543), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n502), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G543), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  OAI211_X1 g086(.A(new_n507), .B(new_n509), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  OAI21_X1  g088(.A(G543), .B1(new_n510), .B2(new_n511), .ZN(new_n514));
  INV_X1    g089(.A(G50), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n505), .A2(new_n516), .ZN(G166));
  INV_X1    g092(.A(new_n514), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G51), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n502), .A2(G63), .A3(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AND3_X1   g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  OR2_X1    g097(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n523));
  NAND2_X1  g098(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  AND2_X1   g101(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n527));
  NOR2_X1   g102(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n525), .A2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  XNOR2_X1  g106(.A(KEYINPUT67), .B(G89), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  XNOR2_X1  g108(.A(KEYINPUT6), .B(G651), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n533), .A2(new_n502), .A3(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n531), .A2(KEYINPUT68), .A3(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT68), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n512), .A2(new_n532), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n537), .B1(new_n538), .B2(new_n530), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n521), .B1(new_n536), .B2(new_n539), .ZN(G168));
  NAND3_X1  g115(.A1(new_n507), .A2(new_n509), .A3(G64), .ZN(new_n541));
  NAND2_X1  g116(.A1(G77), .A2(G543), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G651), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT70), .ZN(new_n545));
  OAI211_X1 g120(.A(G52), .B(G543), .C1(new_n510), .C2(new_n511), .ZN(new_n546));
  XOR2_X1   g121(.A(KEYINPUT69), .B(G90), .Z(new_n547));
  NAND3_X1  g122(.A1(new_n547), .A2(new_n502), .A3(new_n534), .ZN(new_n548));
  NAND4_X1  g123(.A1(new_n544), .A2(new_n545), .A3(new_n546), .A4(new_n548), .ZN(new_n549));
  XNOR2_X1  g124(.A(KEYINPUT69), .B(G90), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n546), .B1(new_n512), .B2(new_n550), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n504), .B1(new_n541), .B2(new_n542), .ZN(new_n552));
  OAI21_X1  g127(.A(KEYINPUT70), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n549), .A2(new_n553), .ZN(G171));
  NAND2_X1  g129(.A1(new_n507), .A2(new_n509), .ZN(new_n555));
  INV_X1    g130(.A(G56), .ZN(new_n556));
  INV_X1    g131(.A(G68), .ZN(new_n557));
  OAI22_X1  g132(.A1(new_n555), .A2(new_n556), .B1(new_n557), .B2(new_n506), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT71), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI221_X1 g135(.A(KEYINPUT71), .B1(new_n557), .B2(new_n506), .C1(new_n555), .C2(new_n556), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n560), .A2(G651), .A3(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(G81), .ZN(new_n563));
  INV_X1    g138(.A(G43), .ZN(new_n564));
  OAI22_X1  g139(.A1(new_n512), .A2(new_n563), .B1(new_n514), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G860), .ZN(G153));
  AND3_X1   g144(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G36), .ZN(G176));
  NAND2_X1  g146(.A1(G1), .A2(G3), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT8), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n570), .A2(new_n573), .ZN(G188));
  OAI211_X1 g149(.A(G53), .B(G543), .C1(new_n510), .C2(new_n511), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(KEYINPUT9), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT9), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n534), .A2(new_n577), .A3(G53), .A4(G543), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n512), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(G91), .ZN(new_n581));
  AND3_X1   g156(.A1(new_n507), .A2(new_n509), .A3(G65), .ZN(new_n582));
  INV_X1    g157(.A(G78), .ZN(new_n583));
  OAI21_X1  g158(.A(KEYINPUT72), .B1(new_n583), .B2(new_n506), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT72), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n585), .A2(G78), .A3(G543), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n582), .B2(new_n587), .ZN(new_n588));
  AND3_X1   g163(.A1(new_n579), .A2(new_n581), .A3(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G299));
  INV_X1    g165(.A(G171), .ZN(G301));
  INV_X1    g166(.A(new_n521), .ZN(new_n592));
  AOI21_X1  g167(.A(KEYINPUT68), .B1(new_n531), .B2(new_n535), .ZN(new_n593));
  NOR3_X1   g168(.A1(new_n538), .A2(new_n530), .A3(new_n537), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(G286));
  INV_X1    g170(.A(G166), .ZN(G303));
  NAND2_X1  g171(.A1(new_n518), .A2(G49), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n597), .B(KEYINPUT73), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n580), .A2(G87), .ZN(new_n599));
  OAI21_X1  g174(.A(G651), .B1(new_n502), .B2(G74), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(G288));
  AOI22_X1  g176(.A1(new_n502), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(new_n504), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n502), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n510), .A2(new_n511), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OR2_X1    g181(.A1(new_n603), .A2(new_n606), .ZN(G305));
  AOI22_X1  g182(.A1(new_n502), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n608), .A2(new_n504), .ZN(new_n609));
  INV_X1    g184(.A(G85), .ZN(new_n610));
  INV_X1    g185(.A(G47), .ZN(new_n611));
  OAI22_X1  g186(.A1(new_n512), .A2(new_n610), .B1(new_n514), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(G290));
  INV_X1    g189(.A(G868), .ZN(new_n615));
  NOR2_X1   g190(.A1(G171), .A2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT74), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(G92), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n512), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT10), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n514), .A2(KEYINPUT75), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT75), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n623), .B(G543), .C1(new_n510), .C2(new_n511), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n622), .A2(G54), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n507), .A2(new_n509), .A3(G66), .ZN(new_n626));
  NAND2_X1  g201(.A1(G79), .A2(G543), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G651), .ZN(new_n629));
  AND3_X1   g204(.A1(new_n625), .A2(KEYINPUT76), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g205(.A(KEYINPUT76), .B1(new_n625), .B2(new_n629), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n621), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g207(.A(KEYINPUT74), .B1(new_n632), .B2(new_n615), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n618), .B1(new_n633), .B2(new_n616), .ZN(G284));
  OAI21_X1  g209(.A(new_n618), .B1(new_n633), .B2(new_n616), .ZN(G321));
  NAND2_X1  g210(.A1(G299), .A2(new_n615), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n636), .B1(G168), .B2(new_n615), .ZN(G297));
  OAI21_X1  g212(.A(new_n636), .B1(G168), .B2(new_n615), .ZN(G280));
  INV_X1    g213(.A(new_n632), .ZN(new_n639));
  INV_X1    g214(.A(G559), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n639), .B1(new_n640), .B2(G860), .ZN(G148));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(G868), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n643), .B1(G868), .B2(new_n568), .ZN(G323));
  XNOR2_X1  g219(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g220(.A1(new_n480), .A2(G2104), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT77), .B(KEYINPUT12), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2100), .ZN(new_n649));
  XOR2_X1   g224(.A(KEYINPUT78), .B(KEYINPUT13), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n480), .A2(G135), .ZN(new_n652));
  OAI21_X1  g227(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n653), .A2(KEYINPUT79), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(KEYINPUT79), .ZN(new_n655));
  OAI211_X1 g230(.A(new_n654), .B(new_n655), .C1(G111), .C2(new_n469), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n478), .A2(G123), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n652), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(G2096), .Z(new_n659));
  NAND2_X1  g234(.A1(new_n651), .A2(new_n659), .ZN(G156));
  XNOR2_X1  g235(.A(KEYINPUT15), .B(G2435), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT80), .B(G2438), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2427), .B(G2430), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n665), .A2(KEYINPUT14), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT81), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1341), .B(G1348), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT16), .B(G2443), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n667), .B(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2451), .B(G2454), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G2446), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n671), .B(new_n673), .Z(new_n674));
  NAND2_X1  g249(.A1(new_n674), .A2(G14), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(G401));
  XOR2_X1   g251(.A(G2072), .B(G2078), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT17), .ZN(new_n678));
  XOR2_X1   g253(.A(G2067), .B(G2678), .Z(new_n679));
  XOR2_X1   g254(.A(G2084), .B(G2090), .Z(new_n680));
  NAND3_X1  g255(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT82), .Z(new_n682));
  INV_X1    g257(.A(new_n680), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n679), .A2(new_n677), .ZN(new_n684));
  OAI211_X1 g259(.A(new_n683), .B(new_n684), .C1(new_n678), .C2(new_n679), .ZN(new_n685));
  NOR3_X1   g260(.A1(new_n683), .A2(new_n679), .A3(new_n677), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT18), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n682), .A2(new_n685), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G2096), .B(G2100), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(G227));
  XNOR2_X1  g266(.A(G1971), .B(G1976), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT19), .ZN(new_n693));
  XOR2_X1   g268(.A(G1956), .B(G2474), .Z(new_n694));
  XOR2_X1   g269(.A(G1961), .B(G1966), .Z(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT20), .Z(new_n698));
  NOR2_X1   g273(.A1(new_n694), .A2(new_n695), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n700), .A2(new_n693), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT83), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n700), .A2(new_n693), .A3(new_n696), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n698), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT84), .B(G1981), .ZN(new_n705));
  XNOR2_X1  g280(.A(G1986), .B(G1991), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n704), .B(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT85), .ZN(new_n710));
  INV_X1    g285(.A(G1996), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n708), .B(new_n712), .ZN(G229));
  INV_X1    g288(.A(G16), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G23), .ZN(new_n715));
  INV_X1    g290(.A(G288), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(new_n716), .B2(new_n714), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT33), .ZN(new_n718));
  INV_X1    g293(.A(G1976), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n714), .A2(G6), .ZN(new_n721));
  INV_X1    g296(.A(G305), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n721), .B1(new_n722), .B2(new_n714), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT32), .B(G1981), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n718), .A2(new_n719), .ZN(new_n726));
  AND2_X1   g301(.A1(KEYINPUT86), .A2(G16), .ZN(new_n727));
  NOR2_X1   g302(.A1(KEYINPUT86), .A2(G16), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G22), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G166), .B2(new_n730), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(G1971), .Z(new_n733));
  NAND4_X1  g308(.A1(new_n720), .A2(new_n725), .A3(new_n726), .A4(new_n733), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT34), .Z(new_n735));
  INV_X1    g310(.A(G29), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(G25), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n478), .A2(G119), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n480), .A2(G131), .ZN(new_n739));
  OR2_X1    g314(.A1(G95), .A2(G2105), .ZN(new_n740));
  OAI211_X1 g315(.A(new_n740), .B(G2104), .C1(G107), .C2(new_n469), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n738), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n737), .B1(new_n743), .B2(new_n736), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT35), .B(G1991), .Z(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n729), .A2(G24), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n613), .B(KEYINPUT87), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n747), .B1(new_n748), .B2(new_n729), .ZN(new_n749));
  INV_X1    g324(.A(G1986), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n735), .A2(new_n746), .A3(new_n751), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT36), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n736), .A2(G33), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT25), .Z(new_n756));
  NAND2_X1  g331(.A1(new_n480), .A2(G139), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n467), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n756), .B(new_n757), .C1(new_n758), .C2(new_n469), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT90), .Z(new_n760));
  OAI21_X1  g335(.A(new_n754), .B1(new_n760), .B2(new_n736), .ZN(new_n761));
  OR2_X1    g336(.A1(KEYINPUT24), .A2(G34), .ZN(new_n762));
  NAND2_X1  g337(.A1(KEYINPUT24), .A2(G34), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n762), .A2(new_n736), .A3(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G160), .B2(new_n736), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n761), .A2(G2072), .B1(G2084), .B2(new_n765), .ZN(new_n766));
  AOI22_X1  g341(.A1(G129), .A2(new_n478), .B1(new_n480), .B2(G141), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n469), .A2(G105), .A3(G2104), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT92), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT91), .B(KEYINPUT26), .ZN(new_n771));
  NAND3_X1  g346(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  OR3_X1    g348(.A1(new_n769), .A2(new_n770), .A3(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n770), .B1(new_n769), .B2(new_n773), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n777), .A2(G29), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT93), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n778), .B(new_n779), .C1(G29), .C2(G32), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(new_n779), .B2(new_n778), .ZN(new_n781));
  XOR2_X1   g356(.A(KEYINPUT27), .B(G1996), .Z(new_n782));
  OAI221_X1 g357(.A(new_n766), .B1(G2072), .B2(new_n761), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT94), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT31), .B(G11), .ZN(new_n785));
  AND2_X1   g360(.A1(new_n781), .A2(new_n782), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n736), .A2(G27), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G164), .B2(new_n736), .ZN(new_n788));
  XOR2_X1   g363(.A(KEYINPUT96), .B(G2078), .Z(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n714), .A2(G21), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G168), .B2(new_n714), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G1966), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n765), .A2(G2084), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n795), .A2(KEYINPUT95), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(KEYINPUT95), .ZN(new_n797));
  INV_X1    g372(.A(new_n658), .ZN(new_n798));
  INV_X1    g373(.A(G28), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n799), .A2(KEYINPUT30), .ZN(new_n800));
  AOI21_X1  g375(.A(G29), .B1(new_n799), .B2(KEYINPUT30), .ZN(new_n801));
  AOI22_X1  g376(.A1(new_n798), .A2(G29), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(G5), .A2(G16), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G171), .B2(G16), .ZN(new_n804));
  INV_X1    g379(.A(G1961), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n796), .A2(new_n797), .A3(new_n802), .A4(new_n806), .ZN(new_n807));
  NOR4_X1   g382(.A1(new_n786), .A2(new_n790), .A3(new_n793), .A4(new_n807), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n784), .A2(new_n785), .A3(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n810), .A2(KEYINPUT97), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n736), .A2(G35), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G162), .B2(new_n736), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT29), .Z(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n815), .A2(G2090), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n478), .A2(G128), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n480), .A2(G140), .ZN(new_n818));
  NOR2_X1   g393(.A1(G104), .A2(G2105), .ZN(new_n819));
  OAI21_X1  g394(.A(G2104), .B1(new_n469), .B2(G116), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n817), .B(new_n818), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(G29), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n736), .A2(G26), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT89), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT28), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(G2067), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n730), .A2(KEYINPUT23), .A3(G20), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT23), .ZN(new_n829));
  INV_X1    g404(.A(G20), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n829), .B1(new_n729), .B2(new_n830), .ZN(new_n831));
  OAI211_X1 g406(.A(new_n828), .B(new_n831), .C1(new_n589), .C2(new_n714), .ZN(new_n832));
  INV_X1    g407(.A(G1956), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n568), .A2(new_n730), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(G19), .B2(new_n730), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(G2090), .ZN(new_n838));
  OAI221_X1 g413(.A(new_n834), .B1(G1341), .B2(new_n837), .C1(new_n814), .C2(new_n838), .ZN(new_n839));
  AOI211_X1 g414(.A(new_n827), .B(new_n839), .C1(G1341), .C2(new_n837), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n714), .A2(G4), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(new_n639), .B2(new_n714), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT88), .Z(new_n843));
  INV_X1    g418(.A(G1348), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n843), .A2(new_n844), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n840), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n847), .B1(new_n810), .B2(KEYINPUT97), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n753), .A2(new_n811), .A3(new_n816), .A4(new_n848), .ZN(G150));
  INV_X1    g424(.A(G150), .ZN(G311));
  NAND2_X1  g425(.A1(new_n580), .A2(G93), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n518), .A2(G55), .ZN(new_n852));
  AOI22_X1  g427(.A1(new_n502), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n851), .B(new_n852), .C1(new_n504), .C2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(G860), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n855), .B(KEYINPUT37), .Z(new_n856));
  NAND2_X1  g431(.A1(new_n639), .A2(G559), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT38), .ZN(new_n858));
  INV_X1    g433(.A(new_n854), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n567), .B(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT39), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n858), .B(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n856), .B1(new_n862), .B2(G860), .ZN(G145));
  XNOR2_X1  g438(.A(new_n776), .B(new_n821), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(new_n500), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT98), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n760), .A2(new_n866), .ZN(new_n867));
  AND2_X1   g442(.A1(new_n760), .A2(new_n866), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n865), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT99), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n478), .A2(G130), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n480), .A2(G142), .ZN(new_n872));
  NOR2_X1   g447(.A1(G106), .A2(G2105), .ZN(new_n873));
  OAI21_X1  g448(.A(G2104), .B1(new_n469), .B2(G118), .ZN(new_n874));
  OAI211_X1 g449(.A(new_n871), .B(new_n872), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n743), .B(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(new_n648), .ZN(new_n877));
  OAI221_X1 g452(.A(new_n869), .B1(new_n870), .B2(new_n877), .C1(new_n867), .C2(new_n865), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n870), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  OR2_X1    g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n878), .A2(new_n880), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n476), .B(new_n658), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(new_n484), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(G37), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n881), .A2(new_n885), .A3(new_n882), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g466(.A(G166), .B(new_n613), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(new_n722), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(new_n716), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(KEYINPUT42), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n625), .A2(new_n629), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT76), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n625), .A2(KEYINPUT76), .A3(new_n629), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n589), .B1(new_n900), .B2(new_n621), .ZN(new_n901));
  OAI211_X1 g476(.A(new_n589), .B(new_n621), .C1(new_n630), .C2(new_n631), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(KEYINPUT41), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT100), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n632), .A2(G299), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT41), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n906), .A2(new_n907), .A3(new_n902), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n904), .A2(new_n905), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n906), .A2(new_n902), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n910), .A2(KEYINPUT100), .A3(KEYINPUT41), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n910), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n567), .B(new_n854), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n642), .B(new_n914), .ZN(new_n915));
  MUX2_X1   g490(.A(new_n912), .B(new_n913), .S(new_n915), .Z(new_n916));
  XNOR2_X1  g491(.A(new_n895), .B(new_n916), .ZN(new_n917));
  OR3_X1    g492(.A1(new_n917), .A2(KEYINPUT101), .A3(new_n615), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n917), .A2(new_n615), .ZN(new_n919));
  AOI21_X1  g494(.A(KEYINPUT101), .B1(new_n854), .B2(new_n615), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n918), .B1(new_n919), .B2(new_n920), .ZN(G295));
  OAI21_X1  g496(.A(new_n918), .B1(new_n919), .B2(new_n920), .ZN(G331));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n923));
  INV_X1    g498(.A(new_n894), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT102), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n549), .A2(new_n553), .A3(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n925), .B1(new_n549), .B2(new_n553), .ZN(new_n928));
  NOR3_X1   g503(.A1(new_n927), .A2(new_n928), .A3(G286), .ZN(new_n929));
  NAND2_X1  g504(.A1(G171), .A2(KEYINPUT102), .ZN(new_n930));
  AOI21_X1  g505(.A(G168), .B1(new_n930), .B2(new_n926), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n860), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(G286), .B1(new_n927), .B2(new_n928), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n930), .A2(G168), .A3(new_n926), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n914), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  AOI22_X1  g510(.A1(new_n932), .A2(new_n935), .B1(new_n904), .B2(new_n908), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT103), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n932), .A2(new_n937), .A3(new_n935), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n914), .A2(new_n933), .A3(new_n934), .A4(KEYINPUT103), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n910), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n924), .B1(new_n936), .B2(new_n940), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n912), .A2(KEYINPUT104), .A3(new_n939), .A4(new_n938), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n938), .A2(new_n911), .A3(new_n909), .A4(new_n939), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT104), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n932), .A2(new_n913), .A3(new_n935), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n942), .A2(new_n945), .A3(new_n894), .A4(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT105), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n947), .A2(new_n948), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n888), .B(new_n941), .C1(new_n949), .C2(new_n950), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n951), .A2(KEYINPUT43), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT43), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n947), .B(new_n948), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n942), .A2(new_n945), .A3(new_n946), .ZN(new_n955));
  AOI21_X1  g530(.A(G37), .B1(new_n955), .B2(new_n924), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n953), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n923), .B1(new_n952), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT107), .ZN(new_n959));
  OAI211_X1 g534(.A(new_n953), .B(new_n956), .C1(new_n949), .C2(new_n950), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT106), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n954), .A2(KEYINPUT106), .A3(new_n953), .A4(new_n956), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n923), .B1(new_n951), .B2(KEYINPUT43), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n959), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  AND4_X1   g541(.A1(new_n959), .A2(new_n965), .A3(new_n962), .A4(new_n963), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n958), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT108), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI211_X1 g545(.A(KEYINPUT108), .B(new_n958), .C1(new_n966), .C2(new_n967), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(G397));
  XNOR2_X1  g547(.A(KEYINPUT109), .B(G1384), .ZN(new_n973));
  AOI21_X1  g548(.A(KEYINPUT45), .B1(new_n500), .B2(new_n973), .ZN(new_n974));
  XOR2_X1   g549(.A(KEYINPUT110), .B(G40), .Z(new_n975));
  NOR2_X1   g550(.A1(new_n476), .A2(new_n975), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n711), .ZN(new_n978));
  XOR2_X1   g553(.A(new_n978), .B(KEYINPUT111), .Z(new_n979));
  NOR2_X1   g554(.A1(new_n979), .A2(new_n776), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n821), .B(G2067), .ZN(new_n981));
  XOR2_X1   g556(.A(new_n981), .B(KEYINPUT112), .Z(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n777), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(new_n977), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n984), .B1(new_n711), .B2(new_n982), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n980), .A2(new_n985), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n742), .B(new_n745), .ZN(new_n987));
  XOR2_X1   g562(.A(new_n987), .B(KEYINPUT113), .Z(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(new_n977), .ZN(new_n989));
  NOR2_X1   g564(.A1(G290), .A2(G1986), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n977), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n991), .B(KEYINPUT48), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n986), .A2(new_n989), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n743), .A2(new_n745), .ZN(new_n994));
  XOR2_X1   g569(.A(new_n994), .B(KEYINPUT126), .Z(new_n995));
  NOR3_X1   g570(.A1(new_n980), .A2(new_n985), .A3(new_n995), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n821), .A2(G2067), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n977), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  AND2_X1   g573(.A1(new_n979), .A2(KEYINPUT46), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n979), .A2(KEYINPUT46), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n984), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n1001), .B(KEYINPUT127), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT47), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n998), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  AOI211_X1 g579(.A(new_n993), .B(new_n1004), .C1(new_n1003), .C2(new_n1002), .ZN(new_n1005));
  AOI21_X1  g580(.A(G1384), .B1(new_n494), .B2(new_n499), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n976), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(G8), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1008), .B1(G1976), .B2(new_n716), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n1010));
  OR2_X1    g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  OAI211_X1 g586(.A(new_n1009), .B(new_n1010), .C1(G1976), .C2(new_n716), .ZN(new_n1012));
  INV_X1    g587(.A(G1981), .ZN(new_n1013));
  XNOR2_X1  g588(.A(G305), .B(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(KEYINPUT116), .A2(KEYINPUT49), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n1014), .B(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1016), .A2(G8), .A3(new_n1007), .ZN(new_n1017));
  AND3_X1   g592(.A1(new_n1011), .A2(new_n1012), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G8), .ZN(new_n1019));
  INV_X1    g594(.A(G1384), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n500), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT45), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n976), .B1(new_n1006), .B2(KEYINPUT45), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  OR2_X1    g600(.A1(new_n1025), .A2(G1966), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1021), .A2(KEYINPUT50), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT50), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1006), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1027), .A2(new_n976), .A3(new_n1029), .ZN(new_n1030));
  OR2_X1    g605(.A1(new_n1030), .A2(G2084), .ZN(new_n1031));
  AOI211_X1 g606(.A(new_n1019), .B(G286), .C1(new_n1026), .C2(new_n1031), .ZN(new_n1032));
  AND3_X1   g607(.A1(new_n1018), .A2(KEYINPUT63), .A3(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n500), .A2(KEYINPUT45), .A3(new_n973), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1035), .A2(new_n1024), .ZN(new_n1036));
  OAI22_X1  g611(.A1(new_n1036), .A2(G1971), .B1(new_n1030), .B2(G2090), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(G8), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT115), .ZN(new_n1039));
  NAND2_X1  g614(.A1(G303), .A2(G8), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1039), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1040), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1045));
  AND3_X1   g620(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT117), .ZN(new_n1047));
  XNOR2_X1  g622(.A(new_n1038), .B(new_n1047), .ZN(new_n1048));
  OR2_X1    g623(.A1(new_n1038), .A2(new_n1046), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1038), .A2(new_n1046), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1018), .A2(new_n1049), .A3(new_n1050), .A4(new_n1032), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT63), .ZN(new_n1052));
  AOI22_X1  g627(.A1(new_n1033), .A2(new_n1048), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1018), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1054), .A2(new_n1049), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1017), .A2(new_n719), .A3(new_n716), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n722), .A2(new_n1013), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1008), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NOR3_X1   g633(.A1(new_n1053), .A2(new_n1055), .A3(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1026), .A2(new_n1031), .A3(G168), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(G8), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(KEYINPUT51), .ZN(new_n1062));
  AOI21_X1  g637(.A(G168), .B1(new_n1026), .B2(new_n1031), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT51), .ZN(new_n1064));
  OAI211_X1 g639(.A(G8), .B(new_n1060), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1062), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT62), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(KEYINPUT62), .B1(new_n1062), .B2(new_n1065), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1071), .A2(G2078), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1025), .A2(new_n1072), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1034), .B(new_n976), .C1(KEYINPUT45), .C2(new_n1006), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1071), .B1(new_n1074), .B2(G2078), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1030), .A2(new_n805), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1073), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(G171), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT121), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1077), .A2(KEYINPUT121), .A3(G171), .ZN(new_n1081));
  AND2_X1   g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1070), .A2(new_n1082), .ZN(new_n1083));
  AND2_X1   g658(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1035), .A2(new_n476), .ZN(new_n1085));
  INV_X1    g660(.A(new_n974), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1085), .A2(G40), .A3(new_n1072), .A4(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(G301), .B1(new_n1084), .B2(new_n1087), .ZN(new_n1088));
  OR2_X1    g663(.A1(new_n1088), .A2(KEYINPUT124), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1084), .A2(G301), .A3(new_n1073), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1084), .A2(new_n1087), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1091), .A2(KEYINPUT124), .A3(G171), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1089), .A2(KEYINPUT54), .A3(new_n1090), .A4(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n1066), .ZN(new_n1094));
  XNOR2_X1  g669(.A(KEYINPUT56), .B(G2072), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1036), .A2(new_n1095), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n1027), .A2(new_n976), .A3(new_n1029), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1096), .B1(G1956), .B2(new_n1097), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n589), .B(KEYINPUT57), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1007), .A2(G2067), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1103), .B1(new_n1030), .B2(new_n844), .ZN(new_n1104));
  AOI21_X1  g679(.A(KEYINPUT119), .B1(new_n1104), .B2(KEYINPUT60), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  OAI22_X1  g681(.A1(new_n1097), .A2(G1348), .B1(G2067), .B2(new_n1007), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT60), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n632), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1104), .A2(KEYINPUT119), .A3(KEYINPUT60), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1106), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n639), .B1(new_n1104), .B2(KEYINPUT60), .ZN(new_n1112));
  AND3_X1   g687(.A1(new_n1104), .A2(KEYINPUT119), .A3(KEYINPUT60), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1112), .B1(new_n1113), .B2(new_n1105), .ZN(new_n1114));
  AOI22_X1  g689(.A1(new_n1036), .A2(new_n1095), .B1(new_n1030), .B2(new_n833), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(new_n1099), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1101), .A2(KEYINPUT61), .A3(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1111), .A2(new_n1114), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1007), .ZN(new_n1119));
  XNOR2_X1  g694(.A(KEYINPUT58), .B(G1341), .ZN(new_n1120));
  OAI22_X1  g695(.A1(new_n1074), .A2(G1996), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(KEYINPUT118), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT118), .ZN(new_n1123));
  OAI221_X1 g698(.A(new_n1123), .B1(new_n1119), .B2(new_n1120), .C1(new_n1074), .C2(G1996), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1122), .A2(new_n568), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT59), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1122), .A2(KEYINPUT59), .A3(new_n1124), .A4(new_n568), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1118), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT61), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1116), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1131), .B1(new_n1102), .B2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1102), .B1(new_n1130), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1116), .A2(new_n639), .A3(new_n1107), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1094), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1084), .A2(KEYINPUT122), .A3(G301), .A4(new_n1087), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1087), .A2(G301), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT122), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1080), .A2(new_n1137), .A3(new_n1081), .A4(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g716(.A(KEYINPUT120), .B(KEYINPUT54), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1141), .A2(KEYINPUT123), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(KEYINPUT123), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1083), .B1(new_n1136), .B2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1018), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1059), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n613), .A2(new_n750), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n977), .B1(new_n990), .B2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n986), .A2(new_n1150), .A3(new_n989), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n1151), .B(KEYINPUT114), .ZN(new_n1152));
  AOI21_X1  g727(.A(KEYINPUT125), .B1(new_n1148), .B2(new_n1152), .ZN(new_n1153));
  AND2_X1   g728(.A1(new_n1111), .A2(new_n1117), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1129), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1154), .A2(new_n1155), .A3(new_n1133), .A4(new_n1114), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1156), .A2(new_n1135), .A3(new_n1101), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1094), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1157), .A2(new_n1158), .A3(new_n1145), .ZN(new_n1159));
  OR2_X1    g734(.A1(new_n1070), .A2(new_n1082), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1147), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1059), .ZN(new_n1162));
  OAI211_X1 g737(.A(KEYINPUT125), .B(new_n1152), .C1(new_n1161), .C2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1005), .B1(new_n1153), .B2(new_n1164), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g740(.A1(new_n890), .A2(new_n675), .A3(new_n690), .ZN(new_n1167));
  NOR2_X1   g741(.A1(G229), .A2(new_n461), .ZN(new_n1168));
  OAI21_X1  g742(.A(new_n1168), .B1(new_n952), .B2(new_n957), .ZN(new_n1169));
  NOR2_X1   g743(.A1(new_n1167), .A2(new_n1169), .ZN(G308));
  INV_X1    g744(.A(G308), .ZN(G225));
endmodule


