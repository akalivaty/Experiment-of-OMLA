

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U551 ( .A1(n695), .A2(n983), .ZN(n694) );
  AND2_X1 U552 ( .A1(n538), .A2(n537), .ZN(G160) );
  NOR2_X2 U553 ( .A1(n626), .A2(n553), .ZN(n644) );
  NOR2_X1 U554 ( .A1(n711), .A2(n710), .ZN(n712) );
  AND2_X1 U555 ( .A1(n692), .A2(n691), .ZN(n695) );
  AND2_X1 U556 ( .A1(n690), .A2(n689), .ZN(n691) );
  BUF_X1 U557 ( .A(n696), .Z(n718) );
  INV_X1 U558 ( .A(KEYINPUT29), .ZN(n715) );
  AND2_X1 U559 ( .A1(n737), .A2(n743), .ZN(n739) );
  INV_X1 U560 ( .A(n990), .ZN(n756) );
  INV_X1 U561 ( .A(KEYINPUT17), .ZN(n522) );
  NOR2_X1 U562 ( .A1(G2105), .A2(G2104), .ZN(n523) );
  NOR2_X1 U563 ( .A1(G651), .A2(n626), .ZN(n643) );
  XNOR2_X1 U564 ( .A(KEYINPUT23), .B(n534), .ZN(n517) );
  OR2_X1 U565 ( .A1(n809), .A2(n946), .ZN(n518) );
  INV_X1 U566 ( .A(n977), .ZN(n689) );
  INV_X1 U567 ( .A(KEYINPUT95), .ZN(n703) );
  XNOR2_X1 U568 ( .A(n703), .B(KEYINPUT27), .ZN(n704) );
  XNOR2_X1 U569 ( .A(n705), .B(n704), .ZN(n707) );
  INV_X1 U570 ( .A(KEYINPUT99), .ZN(n726) );
  XNOR2_X1 U571 ( .A(n726), .B(KEYINPUT30), .ZN(n727) );
  INV_X1 U572 ( .A(KEYINPUT31), .ZN(n732) );
  XNOR2_X1 U573 ( .A(n732), .B(KEYINPUT100), .ZN(n733) );
  NOR2_X1 U574 ( .A1(G1966), .A2(n769), .ZN(n724) );
  NAND2_X1 U575 ( .A1(n736), .A2(n735), .ZN(n743) );
  INV_X1 U576 ( .A(KEYINPUT101), .ZN(n738) );
  INV_X1 U577 ( .A(KEYINPUT64), .ZN(n678) );
  XNOR2_X1 U578 ( .A(n679), .B(n678), .ZN(n696) );
  AND2_X1 U579 ( .A1(n758), .A2(n757), .ZN(n759) );
  NOR2_X1 U580 ( .A1(G164), .A2(G1384), .ZN(n792) );
  NAND2_X1 U581 ( .A1(n805), .A2(n518), .ZN(n806) );
  INV_X1 U582 ( .A(KEYINPUT71), .ZN(n557) );
  XNOR2_X1 U583 ( .A(n557), .B(KEYINPUT13), .ZN(n558) );
  NAND2_X1 U584 ( .A1(G2104), .A2(G2105), .ZN(n525) );
  XNOR2_X1 U585 ( .A(n559), .B(n558), .ZN(n560) );
  INV_X1 U586 ( .A(KEYINPUT83), .ZN(n526) );
  NOR2_X1 U587 ( .A1(G543), .A2(G651), .ZN(n639) );
  XNOR2_X1 U588 ( .A(n527), .B(n526), .ZN(n528) );
  NAND2_X1 U589 ( .A1(n890), .A2(G137), .ZN(n536) );
  NOR2_X1 U590 ( .A1(n531), .A2(n530), .ZN(G164) );
  INV_X1 U591 ( .A(G2105), .ZN(n519) );
  NOR2_X2 U592 ( .A1(G2104), .A2(n519), .ZN(n894) );
  NAND2_X1 U593 ( .A1(G126), .A2(n894), .ZN(n521) );
  AND2_X2 U594 ( .A1(n519), .A2(G2104), .ZN(n891) );
  NAND2_X1 U595 ( .A1(G102), .A2(n891), .ZN(n520) );
  NAND2_X1 U596 ( .A1(n521), .A2(n520), .ZN(n531) );
  XNOR2_X2 U597 ( .A(n523), .B(n522), .ZN(n890) );
  NAND2_X1 U598 ( .A1(G138), .A2(n890), .ZN(n524) );
  XNOR2_X1 U599 ( .A(n524), .B(KEYINPUT84), .ZN(n529) );
  XNOR2_X2 U600 ( .A(n525), .B(KEYINPUT65), .ZN(n896) );
  NAND2_X1 U601 ( .A1(n896), .A2(G114), .ZN(n527) );
  NAND2_X1 U602 ( .A1(n529), .A2(n528), .ZN(n530) );
  NAND2_X1 U603 ( .A1(G125), .A2(n894), .ZN(n533) );
  NAND2_X1 U604 ( .A1(G113), .A2(n896), .ZN(n532) );
  NAND2_X1 U605 ( .A1(n533), .A2(n532), .ZN(n535) );
  NAND2_X1 U606 ( .A1(G101), .A2(n891), .ZN(n534) );
  NOR2_X1 U607 ( .A1(n535), .A2(n517), .ZN(n538) );
  XNOR2_X1 U608 ( .A(n536), .B(KEYINPUT66), .ZN(n537) );
  AND2_X1 U609 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U610 ( .A1(G135), .A2(n890), .ZN(n540) );
  NAND2_X1 U611 ( .A1(G111), .A2(n896), .ZN(n539) );
  NAND2_X1 U612 ( .A1(n540), .A2(n539), .ZN(n543) );
  NAND2_X1 U613 ( .A1(n894), .A2(G123), .ZN(n541) );
  XOR2_X1 U614 ( .A(KEYINPUT18), .B(n541), .Z(n542) );
  NOR2_X1 U615 ( .A1(n543), .A2(n542), .ZN(n545) );
  NAND2_X1 U616 ( .A1(n891), .A2(G99), .ZN(n544) );
  NAND2_X1 U617 ( .A1(n545), .A2(n544), .ZN(n953) );
  XNOR2_X1 U618 ( .A(G2096), .B(n953), .ZN(n546) );
  OR2_X1 U619 ( .A1(G2100), .A2(n546), .ZN(G156) );
  INV_X1 U620 ( .A(G57), .ZN(G237) );
  NAND2_X1 U621 ( .A1(G7), .A2(G661), .ZN(n547) );
  XOR2_X1 U622 ( .A(n547), .B(KEYINPUT10), .Z(n826) );
  NAND2_X1 U623 ( .A1(n826), .A2(G567), .ZN(n548) );
  XOR2_X1 U624 ( .A(KEYINPUT11), .B(n548), .Z(G234) );
  INV_X1 U625 ( .A(G651), .ZN(n553) );
  NOR2_X1 U626 ( .A1(G543), .A2(n553), .ZN(n549) );
  XOR2_X1 U627 ( .A(KEYINPUT1), .B(n549), .Z(n638) );
  NAND2_X1 U628 ( .A1(n638), .A2(G56), .ZN(n550) );
  XOR2_X1 U629 ( .A(KEYINPUT14), .B(n550), .Z(n561) );
  NAND2_X1 U630 ( .A1(n639), .A2(G81), .ZN(n551) );
  XOR2_X1 U631 ( .A(KEYINPUT12), .B(n551), .Z(n556) );
  XNOR2_X1 U632 ( .A(G543), .B(KEYINPUT0), .ZN(n552) );
  XNOR2_X1 U633 ( .A(n552), .B(KEYINPUT67), .ZN(n626) );
  NAND2_X1 U634 ( .A1(n644), .A2(G68), .ZN(n554) );
  XOR2_X1 U635 ( .A(n554), .B(KEYINPUT70), .Z(n555) );
  NOR2_X1 U636 ( .A1(n556), .A2(n555), .ZN(n559) );
  NOR2_X1 U637 ( .A1(n561), .A2(n560), .ZN(n563) );
  NAND2_X1 U638 ( .A1(n643), .A2(G43), .ZN(n562) );
  NAND2_X1 U639 ( .A1(n563), .A2(n562), .ZN(n977) );
  INV_X1 U640 ( .A(G860), .ZN(n603) );
  OR2_X1 U641 ( .A1(n977), .A2(n603), .ZN(G153) );
  NAND2_X1 U642 ( .A1(G64), .A2(n638), .ZN(n565) );
  NAND2_X1 U643 ( .A1(G52), .A2(n643), .ZN(n564) );
  AND2_X1 U644 ( .A1(n565), .A2(n564), .ZN(n571) );
  XNOR2_X1 U645 ( .A(KEYINPUT68), .B(KEYINPUT9), .ZN(n569) );
  NAND2_X1 U646 ( .A1(G77), .A2(n644), .ZN(n567) );
  NAND2_X1 U647 ( .A1(G90), .A2(n639), .ZN(n566) );
  NAND2_X1 U648 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U649 ( .A(n569), .B(n568), .ZN(n570) );
  NAND2_X1 U650 ( .A1(n571), .A2(n570), .ZN(G301) );
  NAND2_X1 U651 ( .A1(G868), .A2(G301), .ZN(n582) );
  NAND2_X1 U652 ( .A1(G54), .A2(n643), .ZN(n573) );
  NAND2_X1 U653 ( .A1(G79), .A2(n644), .ZN(n572) );
  NAND2_X1 U654 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U655 ( .A(KEYINPUT72), .B(n574), .ZN(n578) );
  NAND2_X1 U656 ( .A1(G66), .A2(n638), .ZN(n576) );
  NAND2_X1 U657 ( .A1(G92), .A2(n639), .ZN(n575) );
  NAND2_X1 U658 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U659 ( .A1(n578), .A2(n577), .ZN(n580) );
  XNOR2_X1 U660 ( .A(KEYINPUT73), .B(KEYINPUT15), .ZN(n579) );
  XNOR2_X1 U661 ( .A(n580), .B(n579), .ZN(n983) );
  OR2_X1 U662 ( .A1(n983), .A2(G868), .ZN(n581) );
  NAND2_X1 U663 ( .A1(n582), .A2(n581), .ZN(G284) );
  NAND2_X1 U664 ( .A1(n639), .A2(G89), .ZN(n583) );
  XNOR2_X1 U665 ( .A(n583), .B(KEYINPUT4), .ZN(n585) );
  NAND2_X1 U666 ( .A1(G76), .A2(n644), .ZN(n584) );
  NAND2_X1 U667 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U668 ( .A(KEYINPUT5), .B(n586), .ZN(n592) );
  NAND2_X1 U669 ( .A1(G63), .A2(n638), .ZN(n588) );
  NAND2_X1 U670 ( .A1(G51), .A2(n643), .ZN(n587) );
  NAND2_X1 U671 ( .A1(n588), .A2(n587), .ZN(n590) );
  XOR2_X1 U672 ( .A(KEYINPUT6), .B(KEYINPUT74), .Z(n589) );
  XNOR2_X1 U673 ( .A(n590), .B(n589), .ZN(n591) );
  NAND2_X1 U674 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U675 ( .A(KEYINPUT7), .B(n593), .ZN(G168) );
  XOR2_X1 U676 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U677 ( .A1(G78), .A2(n644), .ZN(n595) );
  NAND2_X1 U678 ( .A1(G91), .A2(n639), .ZN(n594) );
  NAND2_X1 U679 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U680 ( .A(KEYINPUT69), .B(n596), .ZN(n600) );
  NAND2_X1 U681 ( .A1(G65), .A2(n638), .ZN(n598) );
  NAND2_X1 U682 ( .A1(G53), .A2(n643), .ZN(n597) );
  AND2_X1 U683 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U684 ( .A1(n600), .A2(n599), .ZN(G299) );
  INV_X1 U685 ( .A(G868), .ZN(n658) );
  NOR2_X1 U686 ( .A1(G286), .A2(n658), .ZN(n602) );
  NOR2_X1 U687 ( .A1(G868), .A2(G299), .ZN(n601) );
  NOR2_X1 U688 ( .A1(n602), .A2(n601), .ZN(G297) );
  NAND2_X1 U689 ( .A1(n603), .A2(G559), .ZN(n604) );
  NAND2_X1 U690 ( .A1(n604), .A2(n983), .ZN(n605) );
  XNOR2_X1 U691 ( .A(n605), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U692 ( .A1(G868), .A2(n977), .ZN(n608) );
  NAND2_X1 U693 ( .A1(G868), .A2(n983), .ZN(n606) );
  NOR2_X1 U694 ( .A1(G559), .A2(n606), .ZN(n607) );
  NOR2_X1 U695 ( .A1(n608), .A2(n607), .ZN(G282) );
  NAND2_X1 U696 ( .A1(G67), .A2(n638), .ZN(n610) );
  NAND2_X1 U697 ( .A1(G55), .A2(n643), .ZN(n609) );
  NAND2_X1 U698 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U699 ( .A(KEYINPUT76), .B(n611), .ZN(n615) );
  NAND2_X1 U700 ( .A1(G80), .A2(n644), .ZN(n613) );
  NAND2_X1 U701 ( .A1(G93), .A2(n639), .ZN(n612) );
  NAND2_X1 U702 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U703 ( .A1(n615), .A2(n614), .ZN(n657) );
  NAND2_X1 U704 ( .A1(G559), .A2(n983), .ZN(n616) );
  XOR2_X1 U705 ( .A(n977), .B(n616), .Z(n655) );
  XNOR2_X1 U706 ( .A(KEYINPUT75), .B(n655), .ZN(n617) );
  NOR2_X1 U707 ( .A1(G860), .A2(n617), .ZN(n618) );
  XNOR2_X1 U708 ( .A(n657), .B(n618), .ZN(G145) );
  NAND2_X1 U709 ( .A1(G61), .A2(n638), .ZN(n620) );
  NAND2_X1 U710 ( .A1(G48), .A2(n643), .ZN(n619) );
  NAND2_X1 U711 ( .A1(n620), .A2(n619), .ZN(n623) );
  NAND2_X1 U712 ( .A1(n644), .A2(G73), .ZN(n621) );
  XOR2_X1 U713 ( .A(KEYINPUT2), .B(n621), .Z(n622) );
  NOR2_X1 U714 ( .A1(n623), .A2(n622), .ZN(n625) );
  NAND2_X1 U715 ( .A1(n639), .A2(G86), .ZN(n624) );
  NAND2_X1 U716 ( .A1(n625), .A2(n624), .ZN(G305) );
  NAND2_X1 U717 ( .A1(G49), .A2(n643), .ZN(n628) );
  NAND2_X1 U718 ( .A1(G87), .A2(n626), .ZN(n627) );
  NAND2_X1 U719 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U720 ( .A1(n638), .A2(n629), .ZN(n631) );
  NAND2_X1 U721 ( .A1(G651), .A2(G74), .ZN(n630) );
  NAND2_X1 U722 ( .A1(n631), .A2(n630), .ZN(G288) );
  AND2_X1 U723 ( .A1(n638), .A2(G60), .ZN(n635) );
  NAND2_X1 U724 ( .A1(G47), .A2(n643), .ZN(n633) );
  NAND2_X1 U725 ( .A1(G72), .A2(n644), .ZN(n632) );
  NAND2_X1 U726 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U727 ( .A1(n635), .A2(n634), .ZN(n637) );
  NAND2_X1 U728 ( .A1(n639), .A2(G85), .ZN(n636) );
  NAND2_X1 U729 ( .A1(n637), .A2(n636), .ZN(G290) );
  NAND2_X1 U730 ( .A1(n638), .A2(G62), .ZN(n642) );
  NAND2_X1 U731 ( .A1(G88), .A2(n639), .ZN(n640) );
  XOR2_X1 U732 ( .A(KEYINPUT77), .B(n640), .Z(n641) );
  NAND2_X1 U733 ( .A1(n642), .A2(n641), .ZN(n648) );
  NAND2_X1 U734 ( .A1(G50), .A2(n643), .ZN(n646) );
  NAND2_X1 U735 ( .A1(G75), .A2(n644), .ZN(n645) );
  NAND2_X1 U736 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U737 ( .A1(n648), .A2(n647), .ZN(G166) );
  INV_X1 U738 ( .A(G166), .ZN(G303) );
  XOR2_X1 U739 ( .A(G299), .B(n657), .Z(n654) );
  XNOR2_X1 U740 ( .A(KEYINPUT19), .B(G305), .ZN(n649) );
  XNOR2_X1 U741 ( .A(n649), .B(G288), .ZN(n650) );
  XNOR2_X1 U742 ( .A(KEYINPUT78), .B(n650), .ZN(n652) );
  XOR2_X1 U743 ( .A(G290), .B(G303), .Z(n651) );
  XNOR2_X1 U744 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U745 ( .A(n654), .B(n653), .ZN(n863) );
  XNOR2_X1 U746 ( .A(n655), .B(n863), .ZN(n656) );
  NAND2_X1 U747 ( .A1(n656), .A2(G868), .ZN(n660) );
  NAND2_X1 U748 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U749 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U750 ( .A(KEYINPUT79), .B(n661), .ZN(G295) );
  NAND2_X1 U751 ( .A1(G2084), .A2(G2078), .ZN(n662) );
  XOR2_X1 U752 ( .A(KEYINPUT20), .B(n662), .Z(n663) );
  NAND2_X1 U753 ( .A1(G2090), .A2(n663), .ZN(n664) );
  XNOR2_X1 U754 ( .A(KEYINPUT21), .B(n664), .ZN(n665) );
  NAND2_X1 U755 ( .A1(n665), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U756 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U757 ( .A1(G132), .A2(G82), .ZN(n666) );
  XNOR2_X1 U758 ( .A(n666), .B(KEYINPUT80), .ZN(n667) );
  XNOR2_X1 U759 ( .A(n667), .B(KEYINPUT22), .ZN(n668) );
  NOR2_X1 U760 ( .A1(G218), .A2(n668), .ZN(n669) );
  XOR2_X1 U761 ( .A(KEYINPUT81), .B(n669), .Z(n670) );
  NAND2_X1 U762 ( .A1(G96), .A2(n670), .ZN(n830) );
  NAND2_X1 U763 ( .A1(G2106), .A2(n830), .ZN(n671) );
  XNOR2_X1 U764 ( .A(KEYINPUT82), .B(n671), .ZN(n675) );
  NAND2_X1 U765 ( .A1(G69), .A2(G120), .ZN(n672) );
  NOR2_X1 U766 ( .A1(G237), .A2(n672), .ZN(n673) );
  NAND2_X1 U767 ( .A1(G108), .A2(n673), .ZN(n831) );
  NAND2_X1 U768 ( .A1(G567), .A2(n831), .ZN(n674) );
  NAND2_X1 U769 ( .A1(n675), .A2(n674), .ZN(n832) );
  NAND2_X1 U770 ( .A1(G483), .A2(G661), .ZN(n676) );
  NOR2_X1 U771 ( .A1(n832), .A2(n676), .ZN(n829) );
  NAND2_X1 U772 ( .A1(n829), .A2(G36), .ZN(G176) );
  INV_X1 U773 ( .A(G301), .ZN(G171) );
  XOR2_X1 U774 ( .A(G1981), .B(G305), .Z(n978) );
  NAND2_X1 U775 ( .A1(G160), .A2(G40), .ZN(n791) );
  XNOR2_X1 U776 ( .A(n791), .B(KEYINPUT91), .ZN(n677) );
  NAND2_X1 U777 ( .A1(n677), .A2(n792), .ZN(n679) );
  INV_X1 U778 ( .A(n696), .ZN(n744) );
  NAND2_X1 U779 ( .A1(G8), .A2(n744), .ZN(n769) );
  NOR2_X1 U780 ( .A1(G1976), .A2(G288), .ZN(n680) );
  XNOR2_X1 U781 ( .A(KEYINPUT102), .B(n680), .ZN(n754) );
  INV_X1 U782 ( .A(n754), .ZN(n987) );
  NOR2_X1 U783 ( .A1(n769), .A2(n987), .ZN(n681) );
  NAND2_X1 U784 ( .A1(KEYINPUT33), .A2(n681), .ZN(n682) );
  NAND2_X1 U785 ( .A1(n978), .A2(n682), .ZN(n761) );
  INV_X1 U786 ( .A(n724), .ZN(n737) );
  NAND2_X1 U787 ( .A1(G1996), .A2(n696), .ZN(n683) );
  XNOR2_X1 U788 ( .A(n683), .B(KEYINPUT26), .ZN(n685) );
  INV_X1 U789 ( .A(G1341), .ZN(n920) );
  NOR2_X1 U790 ( .A1(n696), .A2(n920), .ZN(n684) );
  NAND2_X1 U791 ( .A1(KEYINPUT26), .A2(n684), .ZN(n688) );
  NAND2_X1 U792 ( .A1(n685), .A2(n688), .ZN(n687) );
  INV_X1 U793 ( .A(KEYINPUT97), .ZN(n686) );
  NAND2_X1 U794 ( .A1(n687), .A2(n686), .ZN(n692) );
  NAND2_X1 U795 ( .A1(n688), .A2(KEYINPUT97), .ZN(n690) );
  INV_X1 U796 ( .A(KEYINPUT98), .ZN(n693) );
  XNOR2_X1 U797 ( .A(n694), .B(n693), .ZN(n702) );
  NAND2_X1 U798 ( .A1(n695), .A2(n983), .ZN(n700) );
  NOR2_X1 U799 ( .A1(G1348), .A2(n718), .ZN(n698) );
  NOR2_X1 U800 ( .A1(n744), .A2(G2067), .ZN(n697) );
  NOR2_X1 U801 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U802 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U803 ( .A1(n702), .A2(n701), .ZN(n709) );
  INV_X1 U804 ( .A(G299), .ZN(n711) );
  NAND2_X1 U805 ( .A1(n718), .A2(G2072), .ZN(n705) );
  XOR2_X1 U806 ( .A(G1956), .B(KEYINPUT96), .Z(n925) );
  NOR2_X1 U807 ( .A1(n925), .A2(n718), .ZN(n706) );
  NOR2_X1 U808 ( .A1(n707), .A2(n706), .ZN(n710) );
  NAND2_X1 U809 ( .A1(n711), .A2(n710), .ZN(n708) );
  NAND2_X1 U810 ( .A1(n709), .A2(n708), .ZN(n714) );
  XOR2_X1 U811 ( .A(n712), .B(KEYINPUT28), .Z(n713) );
  NAND2_X1 U812 ( .A1(n714), .A2(n713), .ZN(n716) );
  XNOR2_X1 U813 ( .A(n716), .B(n715), .ZN(n722) );
  XNOR2_X1 U814 ( .A(KEYINPUT25), .B(G2078), .ZN(n1005) );
  NAND2_X1 U815 ( .A1(n718), .A2(n1005), .ZN(n717) );
  XNOR2_X1 U816 ( .A(n717), .B(KEYINPUT94), .ZN(n720) );
  OR2_X1 U817 ( .A1(n718), .A2(G1961), .ZN(n719) );
  NAND2_X1 U818 ( .A1(n720), .A2(n719), .ZN(n723) );
  NAND2_X1 U819 ( .A1(n723), .A2(G171), .ZN(n721) );
  NAND2_X1 U820 ( .A1(n722), .A2(n721), .ZN(n736) );
  NOR2_X1 U821 ( .A1(G171), .A2(n723), .ZN(n731) );
  NOR2_X1 U822 ( .A1(n744), .A2(G2084), .ZN(n740) );
  NOR2_X1 U823 ( .A1(n740), .A2(n724), .ZN(n725) );
  NAND2_X1 U824 ( .A1(n725), .A2(G8), .ZN(n728) );
  XNOR2_X1 U825 ( .A(n728), .B(n727), .ZN(n729) );
  NOR2_X1 U826 ( .A1(G168), .A2(n729), .ZN(n730) );
  NOR2_X1 U827 ( .A1(n731), .A2(n730), .ZN(n734) );
  XNOR2_X1 U828 ( .A(n734), .B(n733), .ZN(n735) );
  XNOR2_X1 U829 ( .A(n739), .B(n738), .ZN(n742) );
  NAND2_X1 U830 ( .A1(G8), .A2(n740), .ZN(n741) );
  NAND2_X1 U831 ( .A1(n742), .A2(n741), .ZN(n753) );
  NAND2_X1 U832 ( .A1(G286), .A2(n743), .ZN(n749) );
  NOR2_X1 U833 ( .A1(G1971), .A2(n769), .ZN(n746) );
  NOR2_X1 U834 ( .A1(n744), .A2(G2090), .ZN(n745) );
  NOR2_X1 U835 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U836 ( .A1(n747), .A2(G303), .ZN(n748) );
  NAND2_X1 U837 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U838 ( .A1(n750), .A2(G8), .ZN(n751) );
  XNOR2_X1 U839 ( .A(n751), .B(KEYINPUT32), .ZN(n752) );
  NAND2_X1 U840 ( .A1(n753), .A2(n752), .ZN(n768) );
  NOR2_X1 U841 ( .A1(G1971), .A2(G303), .ZN(n989) );
  NOR2_X1 U842 ( .A1(n989), .A2(n754), .ZN(n755) );
  NAND2_X1 U843 ( .A1(n768), .A2(n755), .ZN(n758) );
  NAND2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n990) );
  NOR2_X1 U845 ( .A1(n769), .A2(n756), .ZN(n757) );
  NOR2_X1 U846 ( .A1(KEYINPUT33), .A2(n759), .ZN(n760) );
  NOR2_X1 U847 ( .A1(n761), .A2(n760), .ZN(n774) );
  NOR2_X1 U848 ( .A1(G1981), .A2(G305), .ZN(n762) );
  XOR2_X1 U849 ( .A(KEYINPUT92), .B(n762), .Z(n763) );
  XNOR2_X1 U850 ( .A(KEYINPUT24), .B(n763), .ZN(n764) );
  NOR2_X1 U851 ( .A1(n769), .A2(n764), .ZN(n765) );
  XNOR2_X1 U852 ( .A(n765), .B(KEYINPUT93), .ZN(n772) );
  NOR2_X1 U853 ( .A1(G2090), .A2(G303), .ZN(n766) );
  NAND2_X1 U854 ( .A1(G8), .A2(n766), .ZN(n767) );
  NAND2_X1 U855 ( .A1(n768), .A2(n767), .ZN(n770) );
  NAND2_X1 U856 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U857 ( .A1(n772), .A2(n771), .ZN(n773) );
  NOR2_X1 U858 ( .A1(n774), .A2(n773), .ZN(n807) );
  NAND2_X1 U859 ( .A1(G95), .A2(n891), .ZN(n776) );
  NAND2_X1 U860 ( .A1(G107), .A2(n896), .ZN(n775) );
  NAND2_X1 U861 ( .A1(n776), .A2(n775), .ZN(n779) );
  NAND2_X1 U862 ( .A1(n890), .A2(G131), .ZN(n777) );
  XOR2_X1 U863 ( .A(KEYINPUT88), .B(n777), .Z(n778) );
  NOR2_X1 U864 ( .A1(n779), .A2(n778), .ZN(n781) );
  NAND2_X1 U865 ( .A1(n894), .A2(G119), .ZN(n780) );
  AND2_X1 U866 ( .A1(n781), .A2(n780), .ZN(n903) );
  XNOR2_X1 U867 ( .A(KEYINPUT89), .B(G1991), .ZN(n1010) );
  NOR2_X1 U868 ( .A1(n903), .A2(n1010), .ZN(n790) );
  NAND2_X1 U869 ( .A1(G141), .A2(n890), .ZN(n783) );
  NAND2_X1 U870 ( .A1(G117), .A2(n896), .ZN(n782) );
  NAND2_X1 U871 ( .A1(n783), .A2(n782), .ZN(n786) );
  NAND2_X1 U872 ( .A1(n891), .A2(G105), .ZN(n784) );
  XOR2_X1 U873 ( .A(KEYINPUT38), .B(n784), .Z(n785) );
  NOR2_X1 U874 ( .A1(n786), .A2(n785), .ZN(n788) );
  NAND2_X1 U875 ( .A1(n894), .A2(G129), .ZN(n787) );
  NAND2_X1 U876 ( .A1(n788), .A2(n787), .ZN(n883) );
  AND2_X1 U877 ( .A1(n883), .A2(G1996), .ZN(n789) );
  NOR2_X1 U878 ( .A1(n790), .A2(n789), .ZN(n957) );
  NOR2_X1 U879 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U880 ( .A(KEYINPUT85), .B(n793), .ZN(n809) );
  NOR2_X1 U881 ( .A1(n957), .A2(n809), .ZN(n814) );
  XOR2_X1 U882 ( .A(KEYINPUT90), .B(n814), .Z(n805) );
  XNOR2_X1 U883 ( .A(G2067), .B(KEYINPUT37), .ZN(n818) );
  XNOR2_X1 U884 ( .A(KEYINPUT86), .B(KEYINPUT34), .ZN(n797) );
  NAND2_X1 U885 ( .A1(G140), .A2(n890), .ZN(n795) );
  NAND2_X1 U886 ( .A1(G104), .A2(n891), .ZN(n794) );
  NAND2_X1 U887 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U888 ( .A(n797), .B(n796), .ZN(n803) );
  XNOR2_X1 U889 ( .A(KEYINPUT35), .B(KEYINPUT87), .ZN(n801) );
  NAND2_X1 U890 ( .A1(G128), .A2(n894), .ZN(n799) );
  NAND2_X1 U891 ( .A1(G116), .A2(n896), .ZN(n798) );
  NAND2_X1 U892 ( .A1(n799), .A2(n798), .ZN(n800) );
  XNOR2_X1 U893 ( .A(n801), .B(n800), .ZN(n802) );
  NOR2_X1 U894 ( .A1(n803), .A2(n802), .ZN(n804) );
  XNOR2_X1 U895 ( .A(n804), .B(KEYINPUT36), .ZN(n909) );
  OR2_X1 U896 ( .A1(n818), .A2(n909), .ZN(n946) );
  OR2_X1 U897 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U898 ( .A(n808), .B(KEYINPUT103), .ZN(n811) );
  XNOR2_X1 U899 ( .A(G1986), .B(G290), .ZN(n988) );
  INV_X1 U900 ( .A(n809), .ZN(n820) );
  NAND2_X1 U901 ( .A1(n988), .A2(n820), .ZN(n810) );
  NAND2_X1 U902 ( .A1(n811), .A2(n810), .ZN(n823) );
  NOR2_X1 U903 ( .A1(G1996), .A2(n883), .ZN(n948) );
  NOR2_X1 U904 ( .A1(G1986), .A2(G290), .ZN(n812) );
  AND2_X1 U905 ( .A1(n1010), .A2(n903), .ZN(n955) );
  NOR2_X1 U906 ( .A1(n812), .A2(n955), .ZN(n813) );
  NOR2_X1 U907 ( .A1(n814), .A2(n813), .ZN(n815) );
  NOR2_X1 U908 ( .A1(n948), .A2(n815), .ZN(n816) );
  XNOR2_X1 U909 ( .A(n816), .B(KEYINPUT39), .ZN(n817) );
  NAND2_X1 U910 ( .A1(n817), .A2(n518), .ZN(n819) );
  NAND2_X1 U911 ( .A1(n818), .A2(n909), .ZN(n945) );
  NAND2_X1 U912 ( .A1(n819), .A2(n945), .ZN(n821) );
  NAND2_X1 U913 ( .A1(n821), .A2(n820), .ZN(n822) );
  NAND2_X1 U914 ( .A1(n823), .A2(n822), .ZN(n825) );
  XNOR2_X1 U915 ( .A(KEYINPUT104), .B(KEYINPUT40), .ZN(n824) );
  XNOR2_X1 U916 ( .A(n825), .B(n824), .ZN(G329) );
  NAND2_X1 U917 ( .A1(G2106), .A2(n826), .ZN(G217) );
  INV_X1 U918 ( .A(n826), .ZN(G223) );
  AND2_X1 U919 ( .A1(G15), .A2(G2), .ZN(n827) );
  NAND2_X1 U920 ( .A1(G661), .A2(n827), .ZN(G259) );
  NAND2_X1 U921 ( .A1(G3), .A2(G1), .ZN(n828) );
  NAND2_X1 U922 ( .A1(n829), .A2(n828), .ZN(G188) );
  INV_X1 U924 ( .A(G132), .ZN(G219) );
  INV_X1 U925 ( .A(G120), .ZN(G236) );
  INV_X1 U926 ( .A(G96), .ZN(G221) );
  INV_X1 U927 ( .A(G82), .ZN(G220) );
  INV_X1 U928 ( .A(G69), .ZN(G235) );
  NOR2_X1 U929 ( .A1(n831), .A2(n830), .ZN(G325) );
  INV_X1 U930 ( .A(G325), .ZN(G261) );
  INV_X1 U931 ( .A(n832), .ZN(G319) );
  XOR2_X1 U932 ( .A(G2430), .B(G2451), .Z(n834) );
  XNOR2_X1 U933 ( .A(G2446), .B(G2427), .ZN(n833) );
  XNOR2_X1 U934 ( .A(n834), .B(n833), .ZN(n841) );
  XOR2_X1 U935 ( .A(G2438), .B(G2435), .Z(n836) );
  XNOR2_X1 U936 ( .A(G2443), .B(KEYINPUT105), .ZN(n835) );
  XNOR2_X1 U937 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U938 ( .A(n837), .B(G2454), .Z(n839) );
  XOR2_X1 U939 ( .A(G1348), .B(n920), .Z(n838) );
  XNOR2_X1 U940 ( .A(n839), .B(n838), .ZN(n840) );
  XNOR2_X1 U941 ( .A(n841), .B(n840), .ZN(n842) );
  NAND2_X1 U942 ( .A1(n842), .A2(G14), .ZN(n843) );
  XOR2_X1 U943 ( .A(KEYINPUT106), .B(n843), .Z(G401) );
  XOR2_X1 U944 ( .A(G1956), .B(G1971), .Z(n845) );
  XNOR2_X1 U945 ( .A(G1986), .B(G1976), .ZN(n844) );
  XNOR2_X1 U946 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U947 ( .A(n846), .B(KEYINPUT41), .Z(n848) );
  XNOR2_X1 U948 ( .A(G1981), .B(G1966), .ZN(n847) );
  XNOR2_X1 U949 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U950 ( .A(G2474), .B(G1991), .Z(n850) );
  XNOR2_X1 U951 ( .A(G1961), .B(G1996), .ZN(n849) );
  XNOR2_X1 U952 ( .A(n850), .B(n849), .ZN(n851) );
  XNOR2_X1 U953 ( .A(n852), .B(n851), .ZN(G229) );
  XOR2_X1 U954 ( .A(KEYINPUT108), .B(KEYINPUT107), .Z(n854) );
  XNOR2_X1 U955 ( .A(G2678), .B(KEYINPUT43), .ZN(n853) );
  XNOR2_X1 U956 ( .A(n854), .B(n853), .ZN(n858) );
  XOR2_X1 U957 ( .A(KEYINPUT42), .B(G2090), .Z(n856) );
  XNOR2_X1 U958 ( .A(G2067), .B(G2072), .ZN(n855) );
  XNOR2_X1 U959 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U960 ( .A(n858), .B(n857), .Z(n860) );
  XNOR2_X1 U961 ( .A(G2096), .B(G2100), .ZN(n859) );
  XNOR2_X1 U962 ( .A(n860), .B(n859), .ZN(n862) );
  XOR2_X1 U963 ( .A(G2084), .B(G2078), .Z(n861) );
  XNOR2_X1 U964 ( .A(n862), .B(n861), .ZN(G227) );
  XOR2_X1 U965 ( .A(n863), .B(G286), .Z(n865) );
  XOR2_X1 U966 ( .A(G301), .B(n983), .Z(n864) );
  XNOR2_X1 U967 ( .A(n865), .B(n864), .ZN(n866) );
  XNOR2_X1 U968 ( .A(n866), .B(n977), .ZN(n867) );
  NOR2_X1 U969 ( .A1(G37), .A2(n867), .ZN(G397) );
  NAND2_X1 U970 ( .A1(n894), .A2(G124), .ZN(n868) );
  XNOR2_X1 U971 ( .A(n868), .B(KEYINPUT44), .ZN(n870) );
  NAND2_X1 U972 ( .A1(G112), .A2(n896), .ZN(n869) );
  NAND2_X1 U973 ( .A1(n870), .A2(n869), .ZN(n874) );
  NAND2_X1 U974 ( .A1(G136), .A2(n890), .ZN(n872) );
  NAND2_X1 U975 ( .A1(G100), .A2(n891), .ZN(n871) );
  NAND2_X1 U976 ( .A1(n872), .A2(n871), .ZN(n873) );
  NOR2_X1 U977 ( .A1(n874), .A2(n873), .ZN(G162) );
  NAND2_X1 U978 ( .A1(G142), .A2(n890), .ZN(n876) );
  NAND2_X1 U979 ( .A1(G106), .A2(n891), .ZN(n875) );
  NAND2_X1 U980 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U981 ( .A(n877), .B(KEYINPUT45), .ZN(n882) );
  NAND2_X1 U982 ( .A1(G130), .A2(n894), .ZN(n879) );
  NAND2_X1 U983 ( .A1(G118), .A2(n896), .ZN(n878) );
  NAND2_X1 U984 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U985 ( .A(KEYINPUT109), .B(n880), .ZN(n881) );
  NAND2_X1 U986 ( .A1(n882), .A2(n881), .ZN(n884) );
  XNOR2_X1 U987 ( .A(n884), .B(n883), .ZN(n908) );
  XNOR2_X1 U988 ( .A(KEYINPUT113), .B(KEYINPUT48), .ZN(n886) );
  XNOR2_X1 U989 ( .A(n953), .B(KEYINPUT46), .ZN(n885) );
  XNOR2_X1 U990 ( .A(n886), .B(n885), .ZN(n887) );
  XOR2_X1 U991 ( .A(n887), .B(KEYINPUT112), .Z(n889) );
  XNOR2_X1 U992 ( .A(G164), .B(KEYINPUT110), .ZN(n888) );
  XNOR2_X1 U993 ( .A(n889), .B(n888), .ZN(n902) );
  NAND2_X1 U994 ( .A1(G139), .A2(n890), .ZN(n893) );
  NAND2_X1 U995 ( .A1(G103), .A2(n891), .ZN(n892) );
  NAND2_X1 U996 ( .A1(n893), .A2(n892), .ZN(n901) );
  NAND2_X1 U997 ( .A1(n894), .A2(G127), .ZN(n895) );
  XOR2_X1 U998 ( .A(KEYINPUT111), .B(n895), .Z(n898) );
  NAND2_X1 U999 ( .A1(n896), .A2(G115), .ZN(n897) );
  NAND2_X1 U1000 ( .A1(n898), .A2(n897), .ZN(n899) );
  XOR2_X1 U1001 ( .A(KEYINPUT47), .B(n899), .Z(n900) );
  NOR2_X1 U1002 ( .A1(n901), .A2(n900), .ZN(n958) );
  XOR2_X1 U1003 ( .A(n902), .B(n958), .Z(n905) );
  XNOR2_X1 U1004 ( .A(G160), .B(n903), .ZN(n904) );
  XNOR2_X1 U1005 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U1006 ( .A(G162), .B(n906), .Z(n907) );
  XNOR2_X1 U1007 ( .A(n908), .B(n907), .ZN(n910) );
  XOR2_X1 U1008 ( .A(n910), .B(n909), .Z(n911) );
  NOR2_X1 U1009 ( .A1(G37), .A2(n911), .ZN(n912) );
  XNOR2_X1 U1010 ( .A(KEYINPUT114), .B(n912), .ZN(G395) );
  NOR2_X1 U1011 ( .A1(G229), .A2(G227), .ZN(n913) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(n913), .ZN(n914) );
  NOR2_X1 U1013 ( .A1(G401), .A2(n914), .ZN(n915) );
  AND2_X1 U1014 ( .A1(G319), .A2(n915), .ZN(n917) );
  NOR2_X1 U1015 ( .A1(G397), .A2(G395), .ZN(n916) );
  NAND2_X1 U1016 ( .A1(n917), .A2(n916), .ZN(G225) );
  INV_X1 U1017 ( .A(G225), .ZN(G308) );
  INV_X1 U1018 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1019 ( .A(G16), .B(KEYINPUT124), .Z(n943) );
  XNOR2_X1 U1020 ( .A(KEYINPUT125), .B(G1961), .ZN(n918) );
  XNOR2_X1 U1021 ( .A(n918), .B(G5), .ZN(n933) );
  XNOR2_X1 U1022 ( .A(G1348), .B(KEYINPUT59), .ZN(n919) );
  XNOR2_X1 U1023 ( .A(n919), .B(G4), .ZN(n924) );
  XNOR2_X1 U1024 ( .A(G1981), .B(G6), .ZN(n922) );
  XOR2_X1 U1025 ( .A(n920), .B(G19), .Z(n921) );
  NOR2_X1 U1026 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1027 ( .A1(n924), .A2(n923), .ZN(n928) );
  XOR2_X1 U1028 ( .A(G20), .B(n925), .Z(n926) );
  XNOR2_X1 U1029 ( .A(KEYINPUT126), .B(n926), .ZN(n927) );
  NOR2_X1 U1030 ( .A1(n928), .A2(n927), .ZN(n929) );
  XOR2_X1 U1031 ( .A(KEYINPUT60), .B(n929), .Z(n931) );
  XNOR2_X1 U1032 ( .A(G1966), .B(G21), .ZN(n930) );
  NOR2_X1 U1033 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1034 ( .A1(n933), .A2(n932), .ZN(n940) );
  XNOR2_X1 U1035 ( .A(G1976), .B(G23), .ZN(n935) );
  XNOR2_X1 U1036 ( .A(G1971), .B(G22), .ZN(n934) );
  NOR2_X1 U1037 ( .A1(n935), .A2(n934), .ZN(n937) );
  XOR2_X1 U1038 ( .A(G1986), .B(G24), .Z(n936) );
  NAND2_X1 U1039 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1040 ( .A(KEYINPUT58), .B(n938), .ZN(n939) );
  NOR2_X1 U1041 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1042 ( .A(n941), .B(KEYINPUT61), .ZN(n942) );
  NAND2_X1 U1043 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1044 ( .A1(G11), .A2(n944), .ZN(n975) );
  NAND2_X1 U1045 ( .A1(n946), .A2(n945), .ZN(n968) );
  XOR2_X1 U1046 ( .A(G2090), .B(G162), .Z(n947) );
  NOR2_X1 U1047 ( .A1(n948), .A2(n947), .ZN(n949) );
  XOR2_X1 U1048 ( .A(KEYINPUT51), .B(n949), .Z(n950) );
  XNOR2_X1 U1049 ( .A(KEYINPUT116), .B(n950), .ZN(n966) );
  XOR2_X1 U1050 ( .A(G160), .B(G2084), .Z(n951) );
  XNOR2_X1 U1051 ( .A(KEYINPUT115), .B(n951), .ZN(n952) );
  NAND2_X1 U1052 ( .A1(n953), .A2(n952), .ZN(n954) );
  NOR2_X1 U1053 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1054 ( .A1(n957), .A2(n956), .ZN(n964) );
  XNOR2_X1 U1055 ( .A(G2072), .B(n958), .ZN(n960) );
  XNOR2_X1 U1056 ( .A(G164), .B(G2078), .ZN(n959) );
  NAND2_X1 U1057 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1058 ( .A(KEYINPUT50), .B(n961), .Z(n962) );
  XNOR2_X1 U1059 ( .A(KEYINPUT117), .B(n962), .ZN(n963) );
  NOR2_X1 U1060 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n967) );
  NOR2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n969) );
  XOR2_X1 U1063 ( .A(KEYINPUT52), .B(n969), .Z(n970) );
  NOR2_X1 U1064 ( .A1(KEYINPUT55), .A2(n970), .ZN(n971) );
  XOR2_X1 U1065 ( .A(KEYINPUT118), .B(n971), .Z(n972) );
  NAND2_X1 U1066 ( .A1(n972), .A2(G29), .ZN(n973) );
  XNOR2_X1 U1067 ( .A(KEYINPUT119), .B(n973), .ZN(n974) );
  NOR2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n1003) );
  XOR2_X1 U1069 ( .A(G16), .B(KEYINPUT56), .Z(n976) );
  XNOR2_X1 U1070 ( .A(KEYINPUT123), .B(n976), .ZN(n1001) );
  XOR2_X1 U1071 ( .A(n977), .B(G1341), .Z(n982) );
  XNOR2_X1 U1072 ( .A(G1966), .B(G168), .ZN(n979) );
  NAND2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1074 ( .A(n980), .B(KEYINPUT57), .ZN(n981) );
  NAND2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n985) );
  XOR2_X1 U1076 ( .A(G1348), .B(n983), .Z(n984) );
  NOR2_X1 U1077 ( .A1(n985), .A2(n984), .ZN(n999) );
  NAND2_X1 U1078 ( .A1(G1971), .A2(G303), .ZN(n986) );
  NAND2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n997) );
  XOR2_X1 U1080 ( .A(G299), .B(G1956), .Z(n995) );
  NOR2_X1 U1081 ( .A1(n989), .A2(n988), .ZN(n991) );
  NAND2_X1 U1082 ( .A1(n991), .A2(n990), .ZN(n993) );
  XOR2_X1 U1083 ( .A(G1961), .B(G171), .Z(n992) );
  NOR2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n996) );
  NOR2_X1 U1086 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1087 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1088 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1089 ( .A1(n1003), .A2(n1002), .ZN(n1027) );
  XOR2_X1 U1090 ( .A(G2084), .B(KEYINPUT54), .Z(n1004) );
  XNOR2_X1 U1091 ( .A(G34), .B(n1004), .ZN(n1022) );
  XNOR2_X1 U1092 ( .A(G2090), .B(G35), .ZN(n1020) );
  XOR2_X1 U1093 ( .A(G1996), .B(G32), .Z(n1007) );
  XNOR2_X1 U1094 ( .A(n1005), .B(G27), .ZN(n1006) );
  NAND2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1096 ( .A(KEYINPUT121), .B(n1008), .ZN(n1015) );
  XOR2_X1 U1097 ( .A(G2072), .B(G33), .Z(n1009) );
  NAND2_X1 U1098 ( .A1(n1009), .A2(G28), .ZN(n1013) );
  XOR2_X1 U1099 ( .A(KEYINPUT120), .B(n1010), .Z(n1011) );
  XNOR2_X1 U1100 ( .A(G25), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1017) );
  XNOR2_X1 U1103 ( .A(G26), .B(G2067), .ZN(n1016) );
  NOR2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1105 ( .A(KEYINPUT53), .B(n1018), .ZN(n1019) );
  NOR2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1107 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1108 ( .A(n1023), .B(KEYINPUT55), .ZN(n1024) );
  XNOR2_X1 U1109 ( .A(n1024), .B(KEYINPUT122), .ZN(n1025) );
  NOR2_X1 U1110 ( .A1(G29), .A2(n1025), .ZN(n1026) );
  NOR2_X1 U1111 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XOR2_X1 U1112 ( .A(n1028), .B(KEYINPUT62), .Z(G150) );
  INV_X1 U1113 ( .A(G150), .ZN(G311) );
endmodule

