//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 0 1 1 1 1 0 0 0 0 1 0 0 0 1 1 0 0 1 0 1 0 0 1 0 1 1 1 1 1 1 1 1 1 1 1 0 1 0 1 1 0 1 1 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n630,
    new_n631, new_n633, new_n634, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n788, new_n789, new_n790, new_n791, new_n792, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n853, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887;
  INV_X1    g000(.A(G218gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G43gat), .B(G50gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT15), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT95), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n203), .A2(KEYINPUT15), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  NOR3_X1   g006(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n210));
  AOI22_X1  g009(.A1(new_n209), .A2(new_n210), .B1(G29gat), .B2(G36gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n207), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT96), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT96), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n207), .A2(new_n214), .A3(new_n211), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  XOR2_X1   g015(.A(new_n208), .B(KEYINPUT94), .Z(new_n217));
  INV_X1    g016(.A(new_n210), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n218), .A2(KEYINPUT93), .ZN(new_n219));
  AOI22_X1  g018(.A1(new_n217), .A2(new_n219), .B1(G29gat), .B2(G36gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n220), .B1(new_n219), .B2(new_n217), .ZN(new_n221));
  INV_X1    g020(.A(new_n204), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AOI21_X1  g022(.A(KEYINPUT17), .B1(new_n216), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(G85gat), .A2(G92gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n226), .B(KEYINPUT7), .ZN(new_n227));
  INV_X1    g026(.A(G99gat), .ZN(new_n228));
  INV_X1    g027(.A(G106gat), .ZN(new_n229));
  OAI21_X1  g028(.A(KEYINPUT8), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n227), .B(new_n230), .C1(G85gat), .C2(G92gat), .ZN(new_n231));
  XOR2_X1   g030(.A(G99gat), .B(G106gat), .Z(new_n232));
  XOR2_X1   g031(.A(new_n231), .B(new_n232), .Z(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  AOI22_X1  g033(.A1(new_n213), .A2(new_n215), .B1(new_n222), .B2(new_n221), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT97), .ZN(new_n236));
  AND3_X1   g035(.A1(new_n235), .A2(new_n236), .A3(KEYINPUT17), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n236), .B1(new_n235), .B2(KEYINPUT17), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n225), .B(new_n234), .C1(new_n237), .C2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(G190gat), .ZN(new_n240));
  INV_X1    g039(.A(new_n235), .ZN(new_n241));
  AND2_X1   g040(.A1(G232gat), .A2(G233gat), .ZN(new_n242));
  AOI22_X1  g041(.A1(new_n241), .A2(new_n233), .B1(KEYINPUT41), .B2(new_n242), .ZN(new_n243));
  AND3_X1   g042(.A1(new_n239), .A2(new_n240), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n240), .B1(new_n239), .B2(new_n243), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n202), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n216), .A2(KEYINPUT17), .A3(new_n223), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(KEYINPUT97), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n235), .A2(new_n236), .A3(KEYINPUT17), .ZN(new_n249));
  AOI211_X1 g048(.A(new_n224), .B(new_n233), .C1(new_n248), .C2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n243), .ZN(new_n251));
  OAI21_X1  g050(.A(G190gat), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n239), .A2(new_n240), .A3(new_n243), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n252), .A2(G218gat), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n246), .A2(new_n254), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n255), .A2(KEYINPUT102), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n246), .A2(new_n254), .A3(KEYINPUT101), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n242), .A2(KEYINPUT41), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(G134gat), .ZN(new_n260));
  INV_X1    g059(.A(new_n258), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n246), .A2(new_n254), .A3(KEYINPUT101), .A4(new_n261), .ZN(new_n262));
  AND3_X1   g061(.A1(new_n259), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n260), .B1(new_n259), .B2(new_n262), .ZN(new_n264));
  NOR3_X1   g063(.A1(new_n263), .A2(new_n264), .A3(G162gat), .ZN(new_n265));
  INV_X1    g064(.A(G162gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n259), .A2(new_n262), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(G134gat), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n259), .A2(new_n260), .A3(new_n262), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n266), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n256), .B1(new_n265), .B2(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(G162gat), .B1(new_n263), .B2(new_n264), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n268), .A2(new_n266), .A3(new_n269), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n272), .A2(new_n273), .A3(KEYINPUT102), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G15gat), .B(G22gat), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT16), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n276), .B1(new_n277), .B2(G1gat), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n278), .B1(G1gat), .B2(new_n276), .ZN(new_n279));
  INV_X1    g078(.A(G8gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G57gat), .B(G64gat), .ZN(new_n283));
  XOR2_X1   g082(.A(new_n283), .B(KEYINPUT99), .Z(new_n284));
  NAND2_X1  g083(.A1(G71gat), .A2(G78gat), .ZN(new_n285));
  OR2_X1    g084(.A1(G71gat), .A2(G78gat), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT9), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n284), .A2(new_n288), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n285), .B(new_n286), .C1(new_n283), .C2(new_n287), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n282), .B1(new_n292), .B2(KEYINPUT21), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n293), .B(G183gat), .ZN(new_n294));
  XOR2_X1   g093(.A(G127gat), .B(G155gat), .Z(new_n295));
  XNOR2_X1  g094(.A(new_n294), .B(new_n295), .ZN(new_n296));
  XOR2_X1   g095(.A(KEYINPUT100), .B(G211gat), .Z(new_n297));
  NAND2_X1  g096(.A1(G231gat), .A2(G233gat), .ZN(new_n298));
  XOR2_X1   g097(.A(new_n297), .B(new_n298), .Z(new_n299));
  XNOR2_X1  g098(.A(new_n296), .B(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n292), .A2(KEYINPUT21), .ZN(new_n301));
  XNOR2_X1  g100(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n301), .B(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n300), .B(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n275), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n233), .B(new_n291), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n234), .A2(new_n291), .ZN(new_n307));
  MUX2_X1   g106(.A(new_n306), .B(new_n307), .S(KEYINPUT10), .Z(new_n308));
  NAND2_X1  g107(.A1(G230gat), .A2(G233gat), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n309), .B(KEYINPUT103), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n306), .A2(new_n310), .ZN(new_n313));
  OAI21_X1  g112(.A(KEYINPUT104), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n314), .B1(KEYINPUT104), .B2(new_n313), .ZN(new_n315));
  XNOR2_X1  g114(.A(G176gat), .B(G204gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n316), .B(G148gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n317), .B(KEYINPUT105), .ZN(new_n318));
  INV_X1    g117(.A(G120gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n318), .B(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n315), .B(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n305), .A2(new_n323), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n281), .B(new_n225), .C1(new_n237), .C2(new_n238), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n241), .A2(new_n282), .ZN(new_n326));
  AND2_X1   g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(G229gat), .A2(G233gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n329), .B(KEYINPUT18), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n235), .A2(new_n281), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n331), .B(KEYINPUT98), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(new_n326), .ZN(new_n333));
  XOR2_X1   g132(.A(new_n328), .B(KEYINPUT13), .Z(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AND2_X1   g134(.A1(new_n330), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G113gat), .B(G141gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n337), .B(new_n338), .ZN(new_n339));
  XOR2_X1   g138(.A(G169gat), .B(G197gat), .Z(new_n340));
  XNOR2_X1  g139(.A(new_n339), .B(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n341), .B(KEYINPUT12), .ZN(new_n342));
  OR2_X1    g141(.A1(new_n336), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n336), .A2(new_n342), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT89), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT38), .ZN(new_n347));
  XNOR2_X1  g146(.A(G197gat), .B(G204gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(KEYINPUT69), .B(G211gat), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n350), .A2(new_n202), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n348), .B1(new_n351), .B2(KEYINPUT22), .ZN(new_n352));
  XOR2_X1   g151(.A(new_n352), .B(G211gat), .Z(new_n353));
  XNOR2_X1  g152(.A(new_n353), .B(G218gat), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT29), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT65), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n240), .A2(KEYINPUT64), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT64), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(G190gat), .ZN(new_n359));
  AOI21_X1  g158(.A(G183gat), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(G183gat), .A2(G190gat), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT24), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n356), .B1(new_n360), .B2(new_n365), .ZN(new_n366));
  AND3_X1   g165(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(KEYINPUT64), .B(G190gat), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n369), .B(KEYINPUT65), .C1(G183gat), .C2(new_n370), .ZN(new_n371));
  NOR3_X1   g170(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n374));
  AOI22_X1  g173(.A1(new_n373), .A2(new_n374), .B1(G169gat), .B2(G176gat), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n366), .A2(new_n371), .A3(KEYINPUT25), .A4(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT66), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n374), .ZN(new_n379));
  INV_X1    g178(.A(G169gat), .ZN(new_n380));
  INV_X1    g179(.A(G176gat), .ZN(new_n381));
  OAI22_X1  g180(.A1(new_n379), .A2(new_n372), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n360), .A2(new_n365), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n382), .B1(new_n383), .B2(KEYINPUT65), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT25), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n363), .B(new_n364), .C1(new_n370), .C2(G183gat), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n385), .B1(new_n386), .B2(new_n356), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n384), .A2(new_n387), .A3(KEYINPUT66), .ZN(new_n388));
  INV_X1    g187(.A(G183gat), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n365), .B1(new_n389), .B2(new_n240), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n385), .B1(new_n390), .B2(new_n382), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n378), .A2(new_n388), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n357), .A2(new_n359), .ZN(new_n393));
  XNOR2_X1  g192(.A(KEYINPUT27), .B(G183gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  XOR2_X1   g194(.A(new_n395), .B(KEYINPUT28), .Z(new_n396));
  AOI21_X1  g195(.A(KEYINPUT26), .B1(new_n380), .B2(new_n381), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n397), .B1(new_n380), .B2(new_n381), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n380), .A2(new_n381), .A3(KEYINPUT26), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n396), .A2(new_n398), .A3(new_n399), .A4(new_n361), .ZN(new_n400));
  AND3_X1   g199(.A1(new_n392), .A2(KEYINPUT70), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(KEYINPUT70), .B1(new_n392), .B2(new_n400), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n355), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT71), .ZN(new_n404));
  NAND2_X1  g203(.A1(G226gat), .A2(G233gat), .ZN(new_n405));
  AND3_X1   g204(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n392), .A2(new_n400), .ZN(new_n407));
  INV_X1    g206(.A(new_n405), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT71), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n410), .B1(new_n403), .B2(new_n405), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n354), .B1(new_n406), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(KEYINPUT86), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n407), .A2(new_n355), .A3(new_n405), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT70), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n407), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n392), .A2(KEYINPUT70), .A3(new_n400), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n414), .B1(new_n418), .B2(new_n405), .ZN(new_n419));
  OR2_X1    g218(.A1(new_n419), .A2(new_n354), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT86), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n421), .B(new_n354), .C1(new_n406), .C2(new_n411), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n413), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT37), .ZN(new_n424));
  XOR2_X1   g223(.A(G8gat), .B(G36gat), .Z(new_n425));
  XNOR2_X1  g224(.A(new_n425), .B(G64gat), .ZN(new_n426));
  INV_X1    g225(.A(G92gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n426), .B(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n429));
  INV_X1    g228(.A(new_n354), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n408), .B1(new_n418), .B2(new_n355), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n429), .B(new_n430), .C1(new_n431), .C2(new_n410), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT72), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n433), .B1(new_n419), .B2(new_n354), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n411), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n436), .A2(new_n433), .A3(new_n430), .A4(new_n429), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT37), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  AND4_X1   g239(.A1(new_n347), .A2(new_n424), .A3(new_n428), .A4(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n428), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT73), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  XOR2_X1   g244(.A(G1gat), .B(G29gat), .Z(new_n446));
  XNOR2_X1  g245(.A(G57gat), .B(G85gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n446), .B(new_n447), .ZN(new_n448));
  XNOR2_X1  g247(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n449));
  XOR2_X1   g248(.A(new_n448), .B(new_n449), .Z(new_n450));
  INV_X1    g249(.A(KEYINPUT5), .ZN(new_n451));
  XNOR2_X1  g250(.A(G127gat), .B(G134gat), .ZN(new_n452));
  XOR2_X1   g251(.A(KEYINPUT68), .B(KEYINPUT1), .Z(new_n453));
  XNOR2_X1  g252(.A(KEYINPUT67), .B(G120gat), .ZN(new_n454));
  INV_X1    g253(.A(G113gat), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n319), .A2(G113gat), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n452), .B(new_n453), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  XNOR2_X1  g257(.A(G113gat), .B(G120gat), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n459), .A2(KEYINPUT1), .ZN(new_n460));
  OR2_X1    g259(.A1(new_n460), .A2(new_n452), .ZN(new_n461));
  AND2_X1   g260(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  XOR2_X1   g261(.A(new_n462), .B(KEYINPUT81), .Z(new_n463));
  XNOR2_X1  g262(.A(G155gat), .B(G162gat), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(G141gat), .B(G148gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n466), .B(KEYINPUT74), .ZN(new_n467));
  INV_X1    g266(.A(G155gat), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT2), .B1(new_n468), .B2(new_n266), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n469), .B(KEYINPUT75), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n465), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n469), .ZN(new_n472));
  XNOR2_X1  g271(.A(KEYINPUT77), .B(G148gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(G141gat), .ZN(new_n474));
  INV_X1    g273(.A(G148gat), .ZN(new_n475));
  OR3_X1    g274(.A1(new_n475), .A2(KEYINPUT76), .A3(G141gat), .ZN(new_n476));
  OAI21_X1  g275(.A(KEYINPUT76), .B1(new_n475), .B2(G141gat), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n474), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT78), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n474), .A2(KEYINPUT78), .A3(new_n476), .A4(new_n477), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n472), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n464), .B(KEYINPUT79), .ZN(new_n483));
  AND3_X1   g282(.A1(new_n482), .A2(KEYINPUT80), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(KEYINPUT80), .B1(new_n482), .B2(new_n483), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n471), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n463), .B1(new_n486), .B2(KEYINPUT3), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n482), .A2(new_n483), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT80), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n482), .A2(KEYINPUT80), .A3(new_n483), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT3), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n492), .A2(new_n493), .A3(new_n471), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n487), .A2(new_n494), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n471), .B(new_n462), .C1(new_n484), .C2(new_n485), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT4), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n492), .A2(new_n498), .A3(new_n471), .A4(new_n462), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(G225gat), .A2(G233gat), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n495), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n463), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(new_n486), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(new_n496), .ZN(new_n505));
  INV_X1    g304(.A(new_n501), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n451), .B1(new_n502), .B2(new_n507), .ZN(new_n508));
  AOI22_X1  g307(.A1(new_n494), .A2(new_n487), .B1(new_n497), .B2(new_n499), .ZN(new_n509));
  AOI21_X1  g308(.A(KEYINPUT5), .B1(new_n509), .B2(new_n501), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n450), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n450), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n502), .A2(new_n451), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n501), .B1(new_n504), .B2(new_n496), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n514), .B1(new_n509), .B2(new_n501), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n512), .B(new_n513), .C1(new_n515), .C2(new_n451), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT6), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n511), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n508), .A2(new_n510), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n519), .A2(KEYINPUT6), .A3(new_n512), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n428), .B1(new_n435), .B2(new_n437), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(KEYINPUT73), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n445), .A2(new_n518), .A3(new_n520), .A4(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(KEYINPUT87), .B1(new_n441), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n428), .B1(new_n438), .B2(new_n439), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT88), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(new_n440), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n525), .A2(new_n526), .ZN(new_n529));
  OAI21_X1  g328(.A(KEYINPUT38), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  AND2_X1   g329(.A1(new_n518), .A2(new_n520), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n424), .A2(new_n347), .A3(new_n428), .A4(new_n440), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n521), .B(new_n444), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT87), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n531), .A2(new_n532), .A3(new_n533), .A4(new_n534), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n524), .A2(new_n530), .A3(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT30), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n445), .A2(new_n537), .A3(new_n522), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n435), .A2(new_n437), .A3(new_n428), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n521), .A2(KEYINPUT30), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  OR2_X1    g340(.A1(new_n509), .A2(new_n501), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n542), .B(KEYINPUT39), .C1(new_n506), .C2(new_n505), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n543), .B(new_n450), .C1(KEYINPUT39), .C2(new_n542), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT40), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI22_X1  g345(.A1(new_n544), .A2(new_n545), .B1(new_n512), .B2(new_n519), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n541), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n493), .B1(new_n430), .B2(KEYINPUT29), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(new_n486), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n354), .B1(new_n355), .B2(new_n494), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(G228gat), .A2(G233gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(G22gat), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n550), .A2(G228gat), .A3(G233gat), .A4(new_n552), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT85), .ZN(new_n559));
  XNOR2_X1  g358(.A(G50gat), .B(G78gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(G106gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(KEYINPUT84), .B(KEYINPUT31), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n555), .A2(new_n557), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(G22gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(new_n558), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n559), .A2(new_n566), .A3(new_n558), .A4(new_n563), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n548), .A2(new_n570), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n346), .B1(new_n536), .B2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n407), .B(new_n462), .ZN(new_n573));
  INV_X1    g372(.A(G227gat), .ZN(new_n574));
  INV_X1    g373(.A(G233gat), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(KEYINPUT34), .ZN(new_n577));
  OR3_X1    g376(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(KEYINPUT32), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n577), .B(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(G15gat), .B(G43gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(G71gat), .B(G99gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT33), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n583), .B1(new_n578), .B2(new_n584), .ZN(new_n585));
  OR2_X1    g384(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n580), .A2(new_n585), .ZN(new_n587));
  AND3_X1   g386(.A1(new_n586), .A2(KEYINPUT36), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(KEYINPUT36), .B1(new_n586), .B2(new_n587), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n570), .ZN(new_n591));
  INV_X1    g390(.A(new_n541), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n511), .A2(new_n517), .ZN(new_n593));
  AND2_X1   g392(.A1(new_n593), .A2(KEYINPUT83), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n516), .B1(new_n593), .B2(KEYINPUT83), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n520), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n590), .B1(new_n591), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n524), .A2(new_n530), .A3(new_n535), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n599), .A2(KEYINPUT89), .A3(new_n570), .A4(new_n548), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n572), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n587), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n580), .A2(new_n585), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n570), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT90), .ZN(new_n607));
  OR3_X1    g406(.A1(new_n541), .A2(new_n607), .A3(new_n531), .ZN(new_n608));
  XNOR2_X1  g407(.A(KEYINPUT91), .B(KEYINPUT35), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n607), .B1(new_n541), .B2(new_n531), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n606), .A2(new_n608), .A3(new_n609), .A4(new_n610), .ZN(new_n611));
  OAI21_X1  g410(.A(KEYINPUT35), .B1(new_n605), .B2(new_n597), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n601), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n324), .A2(new_n345), .A3(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT106), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n596), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g419(.A1(new_n616), .A2(new_n592), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n277), .A2(new_n280), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n277), .A2(new_n280), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n621), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT42), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n621), .A2(KEYINPUT42), .A3(new_n623), .A4(new_n624), .ZN(new_n628));
  OAI211_X1 g427(.A(new_n627), .B(new_n628), .C1(new_n280), .C2(new_n621), .ZN(G1325gat));
  AND3_X1   g428(.A1(new_n617), .A2(G15gat), .A3(new_n590), .ZN(new_n630));
  AOI21_X1  g429(.A(G15gat), .B1(new_n617), .B2(new_n604), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n630), .A2(new_n631), .ZN(G1326gat));
  NOR2_X1   g431(.A1(new_n616), .A2(new_n570), .ZN(new_n633));
  XOR2_X1   g432(.A(KEYINPUT43), .B(G22gat), .Z(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(G1327gat));
  INV_X1    g434(.A(new_n304), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n345), .A2(new_n636), .A3(new_n322), .ZN(new_n637));
  AOI211_X1 g436(.A(new_n637), .B(new_n275), .C1(new_n601), .C2(new_n613), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NOR3_X1   g438(.A1(new_n639), .A2(G29gat), .A3(new_n596), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n640), .B(KEYINPUT45), .Z(new_n641));
  INV_X1    g440(.A(KEYINPUT44), .ZN(new_n642));
  INV_X1    g441(.A(new_n275), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT108), .ZN(new_n644));
  AND3_X1   g443(.A1(new_n601), .A2(new_n644), .A3(new_n613), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n644), .B1(new_n601), .B2(new_n613), .ZN(new_n646));
  OAI211_X1 g445(.A(new_n642), .B(new_n643), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n614), .A2(new_n643), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(KEYINPUT44), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n637), .B(KEYINPUT107), .Z(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(G29gat), .B1(new_n653), .B2(new_n596), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n641), .A2(new_n654), .ZN(G1328gat));
  NOR3_X1   g454(.A1(new_n639), .A2(G36gat), .A3(new_n592), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(KEYINPUT46), .ZN(new_n657));
  OAI21_X1  g456(.A(G36gat), .B1(new_n653), .B2(new_n592), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(G1329gat));
  NAND3_X1  g458(.A1(new_n650), .A2(new_n590), .A3(new_n652), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(G43gat), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n275), .B1(new_n601), .B2(new_n613), .ZN(new_n662));
  INV_X1    g461(.A(G43gat), .ZN(new_n663));
  INV_X1    g462(.A(new_n637), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n662), .A2(new_n663), .A3(new_n604), .A4(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(KEYINPUT109), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT109), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n638), .A2(new_n667), .A3(new_n663), .A4(new_n604), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n661), .A2(KEYINPUT47), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT110), .ZN(new_n671));
  AND3_X1   g470(.A1(new_n666), .A2(new_n668), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n671), .B1(new_n666), .B2(new_n668), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AOI211_X1 g473(.A(KEYINPUT111), .B(KEYINPUT47), .C1(new_n674), .C2(new_n661), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT111), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n669), .A2(KEYINPUT110), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n666), .A2(new_n668), .A3(new_n671), .ZN(new_n678));
  INV_X1    g477(.A(new_n590), .ZN(new_n679));
  AOI211_X1 g478(.A(new_n679), .B(new_n651), .C1(new_n647), .C2(new_n649), .ZN(new_n680));
  OAI211_X1 g479(.A(new_n677), .B(new_n678), .C1(new_n680), .C2(new_n663), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT47), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n676), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n670), .B1(new_n675), .B2(new_n683), .ZN(G1330gat));
  NAND4_X1  g483(.A1(new_n650), .A2(G50gat), .A3(new_n591), .A4(new_n652), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n639), .A2(new_n570), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n685), .B1(G50gat), .B2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g487(.A1(new_n645), .A2(new_n646), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n689), .A2(new_n305), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n345), .A2(new_n322), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n692), .A2(new_n596), .ZN(new_n693));
  XOR2_X1   g492(.A(KEYINPUT112), .B(G57gat), .Z(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(G1332gat));
  NOR2_X1   g494(.A1(new_n692), .A2(new_n592), .ZN(new_n696));
  NOR2_X1   g495(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n697));
  AND2_X1   g496(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n696), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n699), .B1(new_n696), .B2(new_n697), .ZN(G1333gat));
  NAND4_X1  g499(.A1(new_n690), .A2(G71gat), .A3(new_n590), .A4(new_n691), .ZN(new_n701));
  AND3_X1   g500(.A1(new_n690), .A2(new_n604), .A3(new_n691), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n701), .B1(new_n702), .B2(G71gat), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g503(.A1(new_n692), .A2(new_n570), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n705), .B(G78gat), .Z(G1335gat));
  INV_X1    g505(.A(new_n345), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(new_n636), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT113), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(new_n323), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(KEYINPUT114), .B1(new_n650), .B2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT114), .ZN(new_n714));
  AOI211_X1 g513(.A(new_n714), .B(new_n710), .C1(new_n647), .C2(new_n649), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n596), .B1(new_n713), .B2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(G85gat), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n662), .A2(new_n709), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT51), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n662), .A2(new_n709), .A3(KEYINPUT51), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n596), .A2(G85gat), .A3(new_n322), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT115), .ZN(new_n726));
  OAI22_X1  g525(.A1(new_n717), .A2(new_n718), .B1(new_n724), .B2(new_n726), .ZN(G1336gat));
  NAND2_X1  g526(.A1(new_n650), .A2(new_n711), .ZN(new_n728));
  OAI21_X1  g527(.A(G92gat), .B1(new_n728), .B2(new_n592), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT52), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n723), .A2(new_n427), .A3(new_n323), .ZN(new_n731));
  OAI211_X1 g530(.A(new_n729), .B(new_n730), .C1(new_n592), .C2(new_n731), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n731), .A2(new_n592), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n541), .B1(new_n712), .B2(new_n715), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n733), .B1(new_n734), .B2(G92gat), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n732), .B1(new_n735), .B2(new_n730), .ZN(G1337gat));
  NOR2_X1   g535(.A1(new_n724), .A2(new_n322), .ZN(new_n737));
  AOI21_X1  g536(.A(G99gat), .B1(new_n737), .B2(new_n604), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n228), .B1(new_n713), .B2(new_n716), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n738), .B1(new_n739), .B2(new_n590), .ZN(G1338gat));
  NAND4_X1  g539(.A1(new_n723), .A2(new_n229), .A3(new_n323), .A4(new_n591), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT53), .ZN(new_n742));
  AOI211_X1 g541(.A(new_n570), .B(new_n710), .C1(new_n647), .C2(new_n649), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n741), .B(new_n742), .C1(new_n743), .C2(new_n229), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT116), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(G106gat), .B1(new_n728), .B2(new_n570), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n747), .A2(KEYINPUT116), .A3(new_n742), .A4(new_n741), .ZN(new_n748));
  INV_X1    g547(.A(new_n741), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n591), .B1(new_n712), .B2(new_n715), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n749), .B1(new_n750), .B2(G106gat), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n746), .B(new_n748), .C1(new_n751), .C2(new_n742), .ZN(G1339gat));
  NOR2_X1   g551(.A1(new_n308), .A2(new_n310), .ZN(new_n753));
  XOR2_X1   g552(.A(new_n753), .B(KEYINPUT117), .Z(new_n754));
  NAND3_X1  g553(.A1(new_n754), .A2(KEYINPUT54), .A3(new_n311), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT54), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n321), .B1(new_n312), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT55), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n315), .A2(new_n320), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n345), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n333), .A2(new_n334), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT118), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n327), .A2(new_n328), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n341), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n344), .A2(new_n323), .A3(new_n767), .ZN(new_n768));
  AND3_X1   g567(.A1(new_n272), .A2(new_n273), .A3(KEYINPUT102), .ZN(new_n769));
  INV_X1    g568(.A(new_n256), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n770), .B1(new_n272), .B2(new_n273), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n763), .B(new_n768), .C1(new_n769), .C2(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n762), .A2(new_n344), .A3(new_n767), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n271), .A2(new_n773), .A3(new_n274), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n772), .A2(new_n636), .A3(new_n774), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n275), .A2(new_n707), .A3(new_n304), .A4(new_n322), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n596), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n777), .A2(new_n606), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n592), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n779), .A2(new_n707), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(new_n455), .ZN(G1340gat));
  OR3_X1    g580(.A1(new_n779), .A2(new_n454), .A3(new_n322), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT119), .ZN(new_n783));
  OAI21_X1  g582(.A(G120gat), .B1(new_n779), .B2(new_n322), .ZN(new_n784));
  AND3_X1   g583(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n783), .B1(new_n782), .B2(new_n784), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n785), .A2(new_n786), .ZN(G1341gat));
  NAND3_X1  g586(.A1(new_n778), .A2(new_n304), .A3(new_n592), .ZN(new_n788));
  INV_X1    g587(.A(G127gat), .ZN(new_n789));
  OR3_X1    g588(.A1(new_n788), .A2(KEYINPUT120), .A3(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(KEYINPUT120), .B1(new_n788), .B2(new_n789), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n792), .B1(new_n789), .B2(new_n788), .ZN(G1342gat));
  NAND3_X1  g592(.A1(new_n778), .A2(new_n643), .A3(new_n592), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(KEYINPUT56), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n260), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(KEYINPUT121), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n794), .A2(KEYINPUT56), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT121), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n795), .A2(new_n799), .A3(new_n260), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n797), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n798), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n799), .B1(new_n795), .B2(new_n260), .ZN(new_n803));
  AOI211_X1 g602(.A(KEYINPUT121), .B(G134gat), .C1(new_n794), .C2(KEYINPUT56), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n801), .A2(new_n805), .ZN(G1343gat));
  NAND2_X1  g605(.A1(new_n775), .A2(new_n776), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n591), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT57), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT123), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n570), .B1(new_n775), .B2(new_n776), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n811), .B1(new_n812), .B2(KEYINPUT57), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n590), .A2(new_n596), .A3(new_n541), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n815), .B(KEYINPUT122), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n808), .A2(new_n811), .A3(new_n809), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n814), .A2(new_n345), .A3(new_n816), .A4(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(G141gat), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n679), .A2(new_n591), .ZN(new_n820));
  AOI211_X1 g619(.A(new_n541), .B(new_n820), .C1(new_n777), .C2(KEYINPUT124), .ZN(new_n821));
  INV_X1    g620(.A(G141gat), .ZN(new_n822));
  OR2_X1    g621(.A1(new_n777), .A2(KEYINPUT124), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n821), .A2(new_n822), .A3(new_n345), .A4(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n819), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(KEYINPUT58), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT58), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n819), .A2(new_n824), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n828), .ZN(G1344gat));
  OAI21_X1  g628(.A(new_n809), .B1(new_n570), .B2(KEYINPUT125), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n812), .B(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n831), .A2(new_n323), .A3(new_n816), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n832), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n821), .A2(new_n823), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n323), .A2(new_n473), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n814), .A2(new_n323), .A3(new_n816), .A4(new_n817), .ZN(new_n836));
  INV_X1    g635(.A(new_n473), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI221_X1 g637(.A(new_n833), .B1(new_n834), .B2(new_n835), .C1(new_n838), .C2(KEYINPUT59), .ZN(G1345gat));
  OAI21_X1  g638(.A(new_n468), .B1(new_n834), .B2(new_n636), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n814), .A2(new_n817), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n841), .A2(new_n304), .A3(new_n816), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n840), .B1(new_n842), .B2(new_n468), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(G1346gat));
  OAI21_X1  g643(.A(new_n266), .B1(new_n834), .B2(new_n275), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n841), .A2(G162gat), .A3(new_n816), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n845), .B1(new_n846), .B2(new_n275), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(G1347gat));
  AOI21_X1  g647(.A(new_n618), .B1(new_n775), .B2(new_n776), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n849), .A2(new_n541), .A3(new_n606), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n345), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g651(.A1(new_n850), .A2(new_n323), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n853), .B(G176gat), .ZN(G1349gat));
  NAND3_X1  g653(.A1(new_n850), .A2(new_n304), .A3(new_n394), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n850), .A2(new_n304), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n855), .B1(new_n856), .B2(new_n389), .ZN(new_n857));
  XNOR2_X1  g656(.A(new_n857), .B(KEYINPUT60), .ZN(G1350gat));
  AOI21_X1  g657(.A(new_n240), .B1(new_n850), .B2(new_n643), .ZN(new_n859));
  OR2_X1    g658(.A1(new_n859), .A2(KEYINPUT61), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n850), .A2(new_n643), .A3(new_n393), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(KEYINPUT61), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(G1351gat));
  NOR3_X1   g662(.A1(new_n590), .A2(new_n592), .A3(new_n570), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n864), .B(KEYINPUT126), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n849), .A2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(G197gat), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n866), .A2(new_n867), .A3(new_n345), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n590), .A2(new_n618), .A3(new_n592), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n831), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n345), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n868), .B1(new_n872), .B2(new_n867), .ZN(G1352gat));
  XNOR2_X1  g672(.A(KEYINPUT127), .B(G204gat), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n866), .A2(new_n323), .A3(new_n875), .ZN(new_n876));
  XOR2_X1   g675(.A(new_n876), .B(KEYINPUT62), .Z(new_n877));
  NAND3_X1  g676(.A1(new_n831), .A2(new_n323), .A3(new_n869), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n877), .B1(new_n875), .B2(new_n879), .ZN(G1353gat));
  NAND3_X1  g679(.A1(new_n866), .A2(new_n304), .A3(new_n350), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n831), .A2(new_n304), .A3(new_n869), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n882), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n883));
  AOI21_X1  g682(.A(KEYINPUT63), .B1(new_n882), .B2(G211gat), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n881), .B1(new_n883), .B2(new_n884), .ZN(G1354gat));
  AOI21_X1  g684(.A(G218gat), .B1(new_n866), .B2(new_n643), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n275), .A2(new_n202), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n886), .B1(new_n870), .B2(new_n887), .ZN(G1355gat));
endmodule


