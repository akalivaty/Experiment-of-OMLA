//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 1 1 1 0 0 0 1 0 1 0 1 0 0 1 0 0 1 0 0 0 1 0 1 0 1 1 1 1 1 0 1 1 1 0 1 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:16 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1275, new_n1276, new_n1278, new_n1279,
    new_n1280, new_n1281, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XOR2_X1   g0003(.A(new_n203), .B(KEYINPUT64), .Z(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT0), .Z(new_n213));
  INV_X1    g0013(.A(KEYINPUT65), .ZN(new_n214));
  INV_X1    g0014(.A(G13), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n214), .B1(new_n207), .B2(new_n215), .ZN(new_n216));
  NAND3_X1  g0016(.A1(KEYINPUT65), .A2(G1), .A3(G13), .ZN(new_n217));
  AND2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n208), .ZN(new_n219));
  OAI21_X1  g0019(.A(G50), .B1(G58), .B2(G68), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT66), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n213), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G68), .ZN(new_n223));
  XNOR2_X1  g0023(.A(KEYINPUT67), .B(G238), .ZN(new_n224));
  XNOR2_X1  g0024(.A(KEYINPUT68), .B(G244), .ZN(new_n225));
  INV_X1    g0025(.A(G77), .ZN(new_n226));
  OAI22_X1  g0026(.A1(new_n223), .A2(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n210), .B1(new_n227), .B2(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n222), .B1(KEYINPUT1), .B2(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  INV_X1    g0035(.A(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT2), .B(G226), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G264), .B(G270), .Z(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT69), .ZN(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G68), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n248), .B(new_n249), .Z(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G351));
  NAND2_X1  g0051(.A1(new_n209), .A2(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n218), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n204), .A2(G20), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n208), .A2(G33), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n208), .A2(new_n260), .A3(KEYINPUT71), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT71), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n262), .B1(G20), .B2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  AOI22_X1  g0064(.A1(new_n257), .A2(new_n259), .B1(new_n264), .B2(G150), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n254), .B1(new_n255), .B2(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n215), .A2(G1), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G20), .ZN(new_n268));
  AND4_X1   g0068(.A1(new_n216), .A2(new_n252), .A3(new_n217), .A4(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n208), .A2(G1), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n269), .A2(G50), .A3(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n272), .B1(G50), .B2(new_n268), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n266), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT9), .ZN(new_n276));
  NAND2_X1  g0076(.A1(G33), .A2(G41), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n277), .A2(G1), .A3(G13), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G274), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G41), .ZN(new_n281));
  INV_X1    g0081(.A(G45), .ZN(new_n282));
  AOI21_X1  g0082(.A(G1), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n280), .A2(KEYINPUT70), .A3(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT70), .ZN(new_n285));
  INV_X1    g0085(.A(new_n283), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n285), .B1(new_n279), .B2(new_n286), .ZN(new_n287));
  AND2_X1   g0087(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  AND2_X1   g0088(.A1(new_n286), .A2(new_n278), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n288), .B1(G226), .B2(new_n289), .ZN(new_n290));
  AND2_X1   g0090(.A1(KEYINPUT3), .A2(G33), .ZN(new_n291));
  NOR2_X1   g0091(.A1(KEYINPUT3), .A2(G33), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n293), .A2(G1698), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G222), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT3), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n260), .ZN(new_n297));
  NAND2_X1  g0097(.A1(KEYINPUT3), .A2(G33), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G223), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(G1698), .ZN(new_n301));
  OAI221_X1 g0101(.A(new_n295), .B1(new_n226), .B2(new_n299), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n216), .A2(new_n217), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n277), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n290), .A2(new_n306), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n275), .A2(new_n276), .B1(new_n307), .B2(G200), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n274), .A2(KEYINPUT9), .ZN(new_n309));
  INV_X1    g0109(.A(G190), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n308), .B(new_n309), .C1(new_n310), .C2(new_n307), .ZN(new_n311));
  XNOR2_X1  g0111(.A(new_n311), .B(KEYINPUT10), .ZN(new_n312));
  INV_X1    g0112(.A(G169), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n274), .B1(new_n307), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G179), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n290), .A2(new_n315), .A3(new_n306), .ZN(new_n316));
  AND2_X1   g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n312), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n202), .B1(new_n261), .B2(new_n263), .ZN(new_n320));
  OAI22_X1  g0120(.A1(new_n258), .A2(new_n226), .B1(new_n208), .B2(G68), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n253), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT11), .ZN(new_n323));
  OR2_X1    g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n322), .A2(new_n323), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n270), .A2(new_n223), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n208), .A2(G68), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT74), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT12), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n267), .B(new_n327), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n330), .B1(KEYINPUT74), .B2(KEYINPUT12), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n267), .A2(new_n327), .A3(new_n328), .A4(new_n329), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n269), .A2(new_n326), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n324), .A2(new_n325), .A3(new_n333), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n284), .A2(new_n287), .B1(G238), .B2(new_n289), .ZN(new_n335));
  INV_X1    g0135(.A(G1698), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n299), .A2(G226), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(G33), .A2(G97), .ZN(new_n338));
  XNOR2_X1  g0138(.A(new_n338), .B(KEYINPUT73), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n337), .B(new_n339), .C1(new_n301), .C2(new_n236), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n305), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n335), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(KEYINPUT13), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT13), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n335), .A2(new_n341), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT14), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n346), .A2(new_n347), .A3(G169), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n343), .A2(G179), .A3(new_n345), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n347), .B1(new_n346), .B2(G169), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n334), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n346), .A2(G200), .ZN(new_n353));
  INV_X1    g0153(.A(new_n334), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n343), .A2(G190), .A3(new_n345), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n352), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(G200), .ZN(new_n358));
  INV_X1    g0158(.A(new_n225), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n288), .B1(new_n359), .B2(new_n289), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n294), .A2(G232), .ZN(new_n361));
  XNOR2_X1  g0161(.A(KEYINPUT72), .B(G107), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  OAI221_X1 g0163(.A(new_n361), .B1(new_n224), .B2(new_n301), .C1(new_n299), .C2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(new_n305), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n358), .B1(new_n360), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n257), .A2(new_n264), .ZN(new_n368));
  XOR2_X1   g0168(.A(KEYINPUT15), .B(G87), .Z(new_n369));
  AOI22_X1  g0169(.A1(new_n369), .A2(new_n259), .B1(G20), .B2(G77), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n254), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n268), .ZN(new_n372));
  NOR4_X1   g0172(.A1(new_n253), .A2(new_n226), .A3(new_n372), .A4(new_n270), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n268), .A2(G77), .ZN(new_n374));
  NOR3_X1   g0174(.A1(new_n371), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n360), .A2(new_n365), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n367), .B(new_n375), .C1(new_n310), .C2(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n375), .B1(new_n376), .B2(new_n313), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(G179), .B2(new_n376), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NOR3_X1   g0180(.A1(new_n319), .A2(new_n357), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n260), .A2(KEYINPUT75), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT75), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(G33), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n292), .B1(new_n385), .B2(KEYINPUT3), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n300), .A2(G1698), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(KEYINPUT78), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(G33), .A2(G87), .ZN(new_n390));
  XNOR2_X1  g0190(.A(KEYINPUT75), .B(G33), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n297), .B1(new_n391), .B2(new_n296), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n392), .A2(G226), .A3(G1698), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT78), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n296), .B1(new_n382), .B2(new_n384), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n394), .B(new_n387), .C1(new_n395), .C2(new_n292), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n389), .A2(new_n390), .A3(new_n393), .A4(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n305), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n284), .A2(new_n287), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n289), .A2(G232), .ZN(new_n400));
  AND2_X1   g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n398), .A2(G179), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n399), .A2(new_n400), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n403), .B1(new_n397), .B2(new_n305), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n402), .B1(new_n313), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT18), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n256), .A2(new_n270), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n269), .A2(new_n407), .B1(new_n372), .B2(new_n256), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n208), .B(new_n297), .C1(new_n391), .C2(new_n296), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT7), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n410), .A2(KEYINPUT76), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n385), .A2(KEYINPUT3), .ZN(new_n413));
  XNOR2_X1  g0213(.A(KEYINPUT76), .B(KEYINPUT7), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n413), .A2(new_n208), .A3(new_n297), .A4(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n412), .A2(new_n415), .A3(G68), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n264), .A2(G159), .ZN(new_n417));
  INV_X1    g0217(.A(G58), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n418), .A2(new_n223), .ZN(new_n419));
  OAI21_X1  g0219(.A(G20), .B1(new_n419), .B2(new_n201), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n416), .A2(KEYINPUT16), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n253), .ZN(new_n424));
  AOI21_X1  g0224(.A(G20), .B1(KEYINPUT3), .B2(G33), .ZN(new_n425));
  OAI211_X1 g0225(.A(KEYINPUT7), .B(new_n425), .C1(new_n385), .C2(KEYINPUT3), .ZN(new_n426));
  AOI21_X1  g0226(.A(KEYINPUT7), .B1(new_n297), .B2(new_n425), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT77), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  AOI211_X1 g0229(.A(KEYINPUT77), .B(KEYINPUT7), .C1(new_n297), .C2(new_n425), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n426), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(G68), .ZN(new_n432));
  AOI21_X1  g0232(.A(KEYINPUT16), .B1(new_n432), .B2(new_n422), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n408), .B1(new_n424), .B2(new_n433), .ZN(new_n434));
  AND3_X1   g0234(.A1(new_n405), .A2(new_n406), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n406), .B1(new_n405), .B2(new_n434), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT17), .ZN(new_n438));
  AND4_X1   g0238(.A1(KEYINPUT79), .A2(new_n398), .A3(new_n310), .A4(new_n401), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n404), .A2(new_n310), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT79), .B1(new_n404), .B2(G200), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n438), .B1(new_n442), .B2(new_n434), .ZN(new_n443));
  INV_X1    g0243(.A(new_n434), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n398), .A2(new_n401), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(new_n358), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n446), .A2(KEYINPUT79), .B1(new_n310), .B2(new_n404), .ZN(new_n447));
  OAI211_X1 g0247(.A(KEYINPUT17), .B(new_n444), .C1(new_n447), .C2(new_n439), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n437), .A2(new_n443), .A3(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n381), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n268), .A2(G97), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n207), .A2(G33), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n218), .A2(new_n252), .A3(new_n268), .A4(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n453), .B1(new_n456), .B2(G97), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n226), .B1(new_n261), .B2(new_n263), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(G107), .ZN(new_n460));
  AND3_X1   g0260(.A1(new_n460), .A2(KEYINPUT6), .A3(G97), .ZN(new_n461));
  XNOR2_X1  g0261(.A(G97), .B(G107), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT6), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n459), .B1(new_n464), .B2(new_n208), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n465), .B1(new_n431), .B2(new_n362), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT80), .ZN(new_n467));
  NOR3_X1   g0267(.A1(new_n466), .A2(new_n467), .A3(new_n254), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n462), .A2(new_n463), .ZN(new_n469));
  INV_X1    g0269(.A(new_n461), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n458), .B1(new_n471), .B2(G20), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n298), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n473), .B1(new_n391), .B2(new_n296), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n298), .A2(new_n208), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n410), .B1(new_n475), .B2(new_n292), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT77), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n427), .A2(new_n428), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n474), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n472), .B1(new_n479), .B2(new_n363), .ZN(new_n480));
  AOI21_X1  g0280(.A(KEYINPUT80), .B1(new_n480), .B2(new_n253), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n457), .B1(new_n468), .B2(new_n481), .ZN(new_n482));
  XNOR2_X1  g0282(.A(KEYINPUT5), .B(G41), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n282), .A2(G1), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n485), .A2(new_n279), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n278), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n486), .B1(new_n488), .B2(G257), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n299), .A2(G250), .A3(G1698), .ZN(new_n490));
  AND2_X1   g0290(.A1(KEYINPUT4), .A2(G244), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n299), .A2(new_n336), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(G33), .A2(G283), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT82), .ZN(new_n494));
  XNOR2_X1  g0294(.A(new_n493), .B(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n490), .A2(new_n492), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT4), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n392), .A2(G244), .A3(new_n336), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n489), .B1(new_n499), .B2(new_n304), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(G169), .ZN(new_n501));
  OAI211_X1 g0301(.A(G179), .B(new_n489), .C1(new_n499), .C2(new_n304), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n482), .A2(new_n503), .ZN(new_n504));
  AND3_X1   g0304(.A1(new_n485), .A2(G264), .A3(new_n278), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n392), .A2(G257), .A3(G1698), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n392), .A2(G250), .A3(new_n336), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n385), .A2(G294), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n505), .B1(new_n509), .B2(new_n305), .ZN(new_n510));
  INV_X1    g0310(.A(new_n486), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(KEYINPUT89), .B1(new_n512), .B2(G190), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n358), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT89), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n510), .A2(new_n515), .A3(new_n310), .A4(new_n511), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n513), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n208), .B(G87), .C1(new_n395), .C2(new_n292), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT22), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT22), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n520), .A2(new_n208), .A3(G87), .ZN(new_n521));
  OAI21_X1  g0321(.A(KEYINPUT86), .B1(new_n293), .B2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT86), .ZN(new_n523));
  INV_X1    g0323(.A(G87), .ZN(new_n524));
  NOR3_X1   g0324(.A1(new_n524), .A2(KEYINPUT22), .A3(G20), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n299), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n519), .A2(new_n522), .A3(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT87), .ZN(new_n528));
  AOI21_X1  g0328(.A(KEYINPUT23), .B1(new_n385), .B2(G116), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n529), .A2(G20), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT23), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n531), .A2(new_n460), .A3(G20), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n532), .B1(new_n363), .B2(new_n531), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n527), .A2(new_n528), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n522), .A2(new_n526), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n536), .B1(KEYINPUT22), .B2(new_n518), .ZN(new_n537));
  OAI221_X1 g0337(.A(new_n532), .B1(new_n531), .B2(new_n363), .C1(new_n529), .C2(G20), .ZN(new_n538));
  OAI21_X1  g0338(.A(KEYINPUT87), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT24), .ZN(new_n540));
  AND3_X1   g0340(.A1(new_n535), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n540), .B1(new_n535), .B2(new_n539), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n253), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT25), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(new_n268), .B2(G107), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n372), .A2(KEYINPUT25), .A3(new_n460), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n456), .A2(G107), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n517), .A2(new_n543), .A3(new_n547), .ZN(new_n548));
  MUX2_X1   g0348(.A(new_n310), .B(new_n358), .S(new_n500), .Z(new_n549));
  NAND2_X1  g0349(.A1(new_n482), .A2(KEYINPUT81), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n467), .B1(new_n466), .B2(new_n254), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n480), .A2(KEYINPUT80), .A3(new_n253), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT81), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n553), .A2(new_n554), .A3(new_n457), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n549), .A2(new_n550), .A3(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n392), .A2(new_n208), .A3(G68), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT19), .ZN(new_n558));
  INV_X1    g0358(.A(G97), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n558), .B1(new_n258), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT73), .ZN(new_n561));
  XNOR2_X1  g0361(.A(new_n338), .B(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(G20), .B1(new_n562), .B2(KEYINPUT19), .ZN(new_n563));
  NOR3_X1   g0363(.A1(new_n362), .A2(G87), .A3(G97), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n557), .B(new_n560), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n253), .ZN(new_n566));
  INV_X1    g0366(.A(new_n369), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n372), .ZN(new_n568));
  OAI21_X1  g0368(.A(KEYINPUT84), .B1(new_n455), .B2(new_n524), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT84), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n269), .A2(new_n570), .A3(G87), .A4(new_n454), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n566), .A2(new_n568), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n392), .A2(G244), .A3(G1698), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n392), .A2(G238), .A3(new_n336), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n385), .A2(G116), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n305), .ZN(new_n578));
  INV_X1    g0378(.A(new_n484), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n579), .A2(G250), .A3(new_n278), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(new_n279), .B2(new_n579), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(KEYINPUT83), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT83), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n580), .B(new_n583), .C1(new_n279), .C2(new_n579), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n578), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(G200), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n577), .A2(new_n305), .B1(new_n582), .B2(new_n584), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(G190), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n573), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n586), .A2(new_n313), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n566), .B(new_n568), .C1(new_n567), .C2(new_n455), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n588), .A2(new_n315), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  AND4_X1   g0396(.A1(new_n504), .A2(new_n548), .A3(new_n556), .A4(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT88), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n543), .A2(new_n547), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n512), .A2(new_n313), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n510), .A2(new_n315), .A3(new_n511), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n598), .B1(new_n599), .B2(new_n603), .ZN(new_n604));
  AOI211_X1 g0404(.A(KEYINPUT88), .B(new_n602), .C1(new_n543), .C2(new_n547), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n392), .A2(G257), .A3(new_n336), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n392), .A2(G264), .A3(G1698), .ZN(new_n608));
  INV_X1    g0408(.A(G303), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n607), .B(new_n608), .C1(new_n609), .C2(new_n299), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n305), .ZN(new_n611));
  INV_X1    g0411(.A(G270), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n511), .B1(new_n612), .B2(new_n487), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(G116), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n268), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n617), .B1(new_n456), .B2(new_n616), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n495), .B(new_n208), .C1(G33), .C2(new_n559), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT20), .ZN(new_n620));
  AOI22_X1  g0420(.A1(KEYINPUT85), .A2(new_n620), .B1(new_n616), .B2(G20), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n619), .A2(new_n253), .A3(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n620), .A2(KEYINPUT85), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n623), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n619), .A2(new_n253), .A3(new_n621), .A4(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n618), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n615), .A2(new_n627), .A3(G169), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT21), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n613), .B1(new_n610), .B2(new_n305), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n627), .A2(new_n631), .A3(G179), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n615), .A2(new_n627), .A3(KEYINPUT21), .A4(G169), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n630), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n615), .A2(new_n310), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n631), .A2(new_n358), .ZN(new_n636));
  NOR3_X1   g0436(.A1(new_n635), .A2(new_n627), .A3(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  AND4_X1   g0438(.A1(new_n452), .A2(new_n597), .A3(new_n606), .A4(new_n638), .ZN(G372));
  INV_X1    g0439(.A(KEYINPUT26), .ZN(new_n640));
  NOR3_X1   g0440(.A1(new_n595), .A2(new_n504), .A3(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n503), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n643), .B1(new_n550), .B2(new_n555), .ZN(new_n644));
  AOI21_X1  g0444(.A(KEYINPUT26), .B1(new_n644), .B2(new_n596), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT90), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n642), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n554), .B1(new_n553), .B2(new_n457), .ZN(new_n648));
  INV_X1    g0448(.A(new_n457), .ZN(new_n649));
  AOI211_X1 g0449(.A(KEYINPUT81), .B(new_n649), .C1(new_n551), .C2(new_n552), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n503), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n640), .B1(new_n651), .B2(new_n595), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n652), .A2(KEYINPUT90), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n594), .B1(new_n647), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(KEYINPUT91), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT91), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n656), .B(new_n594), .C1(new_n647), .C2(new_n653), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n528), .B1(new_n527), .B2(new_n534), .ZN(new_n658));
  NOR3_X1   g0458(.A1(new_n537), .A2(new_n538), .A3(KEYINPUT87), .ZN(new_n659));
  OAI21_X1  g0459(.A(KEYINPUT24), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n535), .A2(new_n539), .A3(new_n540), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n254), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n547), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n603), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n597), .B1(new_n665), .B2(new_n634), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n655), .A2(new_n657), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n452), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g0468(.A(new_n668), .B(KEYINPUT92), .Z(new_n669));
  INV_X1    g0469(.A(new_n356), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n352), .B1(new_n670), .B2(new_n379), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n671), .A2(new_n443), .A3(new_n448), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n437), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT93), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n675), .A2(new_n312), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n672), .A2(KEYINPUT93), .A3(new_n437), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n317), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n669), .A2(new_n678), .ZN(G369));
  INV_X1    g0479(.A(KEYINPUT95), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n267), .A2(new_n208), .ZN(new_n681));
  OR2_X1    g0481(.A1(new_n681), .A2(KEYINPUT27), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(KEYINPUT27), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(G213), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g0484(.A(KEYINPUT94), .B(G343), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n599), .A2(new_n686), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n687), .A2(new_n548), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n606), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n665), .A2(new_n686), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n634), .ZN(new_n692));
  INV_X1    g0492(.A(new_n627), .ZN(new_n693));
  INV_X1    g0493(.A(new_n686), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n634), .A2(new_n637), .A3(new_n695), .ZN(new_n698));
  OAI21_X1  g0498(.A(G330), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n680), .B1(new_n691), .B2(new_n700), .ZN(new_n701));
  AOI211_X1 g0501(.A(KEYINPUT95), .B(new_n699), .C1(new_n689), .C2(new_n690), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n665), .A2(new_n694), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n692), .A2(new_n686), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n606), .A2(new_n688), .A3(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n704), .A2(new_n705), .A3(new_n707), .ZN(G399));
  INV_X1    g0508(.A(new_n211), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(G41), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n564), .A2(new_n616), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n711), .A2(G1), .A3(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n221), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n714), .B1(new_n715), .B2(new_n711), .ZN(new_n716));
  XNOR2_X1  g0516(.A(new_n716), .B(KEYINPUT96), .ZN(new_n717));
  XNOR2_X1  g0517(.A(new_n717), .B(KEYINPUT28), .ZN(new_n718));
  AND2_X1   g0518(.A1(new_n631), .A2(new_n510), .ZN(new_n719));
  INV_X1    g0519(.A(new_n502), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n719), .A2(new_n720), .A3(KEYINPUT30), .A4(new_n588), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT30), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n631), .A2(new_n588), .A3(new_n510), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n722), .B1(new_n723), .B2(new_n502), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n631), .A2(G179), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n725), .A2(new_n512), .A3(new_n500), .A4(new_n586), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n721), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n727), .A2(KEYINPUT31), .A3(new_n686), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT97), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n727), .A2(KEYINPUT97), .A3(KEYINPUT31), .A4(new_n686), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n727), .A2(new_n686), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT31), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n730), .A2(new_n731), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(KEYINPUT98), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n606), .A2(new_n597), .A3(new_n638), .A4(new_n694), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT98), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n730), .A2(new_n734), .A3(new_n738), .A4(new_n731), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n736), .A2(new_n737), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G330), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n667), .A2(new_n694), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT29), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n664), .A2(KEYINPUT88), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n599), .A2(new_n598), .A3(new_n603), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n746), .A2(new_n747), .A3(new_n692), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(new_n597), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n640), .B1(new_n644), .B2(new_n596), .ZN(new_n750));
  XOR2_X1   g0550(.A(new_n594), .B(KEYINPUT99), .Z(new_n751));
  NOR3_X1   g0551(.A1(new_n595), .A2(new_n504), .A3(KEYINPUT26), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n686), .B1(new_n749), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(KEYINPUT29), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n742), .B1(new_n745), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n718), .B1(new_n756), .B2(G1), .ZN(G364));
  INV_X1    g0557(.A(new_n697), .ZN(new_n758));
  INV_X1    g0558(.A(G330), .ZN(new_n759));
  INV_X1    g0559(.A(new_n698), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n215), .A2(G20), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n207), .B1(new_n762), .B2(G45), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n710), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n761), .A2(new_n699), .A3(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G13), .A2(G33), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(G20), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n758), .A2(new_n760), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n211), .A2(new_n299), .ZN(new_n772));
  INV_X1    g0572(.A(G355), .ZN(new_n773));
  OAI22_X1  g0573(.A1(new_n772), .A2(new_n773), .B1(G116), .B2(new_n211), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n774), .B(KEYINPUT100), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n709), .A2(new_n392), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n221), .A2(new_n282), .ZN(new_n777));
  OAI211_X1 g0577(.A(new_n776), .B(new_n777), .C1(new_n250), .C2(new_n282), .ZN(new_n778));
  AND2_X1   g0578(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n779), .A2(KEYINPUT101), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(KEYINPUT101), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n218), .B1(G20), .B2(new_n313), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n770), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n780), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n208), .A2(new_n315), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G200), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(G190), .ZN(new_n787));
  AND2_X1   g0587(.A1(new_n787), .A2(KEYINPUT103), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n787), .A2(KEYINPUT103), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  XNOR2_X1  g0591(.A(KEYINPUT33), .B(G317), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n785), .A2(G190), .A3(new_n358), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n208), .A2(G179), .ZN(new_n796));
  NOR2_X1   g0596(.A1(G190), .A2(G200), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n795), .A2(G322), .B1(new_n799), .B2(G329), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n785), .A2(new_n797), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n299), .B1(new_n802), .B2(G311), .ZN(new_n803));
  AND2_X1   g0603(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  NOR3_X1   g0604(.A1(new_n310), .A2(G179), .A3(G200), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(new_n208), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n796), .A2(G190), .A3(G200), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n807), .A2(G294), .B1(new_n809), .B2(G303), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n786), .A2(new_n310), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n796), .A2(new_n310), .A3(G200), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n811), .A2(G326), .B1(new_n813), .B2(G283), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n793), .A2(new_n804), .A3(new_n810), .A4(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n812), .A2(new_n460), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n293), .B(new_n816), .C1(G87), .C2(new_n809), .ZN(new_n817));
  XOR2_X1   g0617(.A(new_n817), .B(KEYINPUT102), .Z(new_n818));
  NAND2_X1  g0618(.A1(new_n791), .A2(G68), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n794), .A2(new_n418), .B1(new_n801), .B2(new_n226), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT32), .ZN(new_n821));
  INV_X1    g0621(.A(G159), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n798), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n820), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n807), .A2(G97), .ZN(new_n825));
  INV_X1    g0625(.A(new_n823), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n826), .A2(KEYINPUT32), .B1(new_n811), .B2(G50), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n819), .A2(new_n824), .A3(new_n825), .A4(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n815), .B1(new_n818), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n766), .B1(new_n829), .B2(new_n782), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n771), .A2(new_n784), .A3(new_n830), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n767), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(G396));
  NOR2_X1   g0633(.A1(new_n379), .A2(new_n686), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n377), .B1(new_n375), .B2(new_n694), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n834), .B1(new_n835), .B2(new_n379), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n836), .A2(new_n769), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n791), .A2(G283), .ZN(new_n838));
  INV_X1    g0638(.A(G294), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n794), .A2(new_n839), .B1(new_n801), .B2(new_n616), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n299), .B(new_n840), .C1(G311), .C2(new_n799), .ZN(new_n841));
  AOI22_X1  g0641(.A1(G97), .A2(new_n807), .B1(new_n811), .B2(G303), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n812), .A2(new_n524), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(G107), .B2(new_n809), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n838), .A2(new_n841), .A3(new_n842), .A4(new_n844), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n807), .A2(G58), .B1(new_n813), .B2(G68), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(new_n202), .B2(new_n808), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n386), .B(new_n847), .C1(G132), .C2(new_n799), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n795), .A2(G143), .B1(new_n802), .B2(G159), .ZN(new_n849));
  INV_X1    g0649(.A(G137), .ZN(new_n850));
  INV_X1    g0650(.A(new_n811), .ZN(new_n851));
  INV_X1    g0651(.A(G150), .ZN(new_n852));
  OAI221_X1 g0652(.A(new_n849), .B1(new_n850), .B2(new_n851), .C1(new_n790), .C2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT34), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n848), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n853), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n856), .A2(KEYINPUT34), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n845), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n782), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n782), .A2(new_n768), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n859), .B(new_n765), .C1(G77), .C2(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n837), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n836), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n743), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n380), .A2(new_n686), .ZN(new_n866));
  INV_X1    g0666(.A(new_n594), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n641), .B1(new_n652), .B2(KEYINPUT90), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n645), .A2(new_n646), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n666), .B1(new_n870), .B2(new_n656), .ZN(new_n871));
  INV_X1    g0671(.A(new_n657), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n866), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n865), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n874), .A2(new_n741), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n765), .B1(new_n874), .B2(new_n741), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n863), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(G384));
  NOR2_X1   g0679(.A1(new_n762), .A2(new_n207), .ZN(new_n880));
  AOI21_X1  g0680(.A(KEYINPUT16), .B1(new_n416), .B2(new_n422), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n408), .B1(new_n424), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(KEYINPUT104), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT104), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n884), .B(new_n408), .C1(new_n424), .C2(new_n881), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n684), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n405), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n442), .A2(new_n434), .ZN(new_n890));
  OAI21_X1  g0690(.A(KEYINPUT37), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT106), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n892), .B1(new_n434), .B2(new_n887), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n434), .A2(new_n892), .A3(new_n887), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n444), .B1(new_n447), .B2(new_n439), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT37), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n405), .A2(new_n434), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n896), .A2(new_n897), .A3(new_n898), .A4(new_n899), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n891), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n886), .A2(new_n684), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n449), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(KEYINPUT105), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT105), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n449), .A2(new_n905), .A3(new_n902), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n901), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n907), .A2(KEYINPUT38), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n891), .A2(new_n900), .ZN(new_n909));
  AND3_X1   g0709(.A1(new_n449), .A2(new_n905), .A3(new_n902), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n905), .B1(new_n449), .B2(new_n902), .ZN(new_n911));
  OAI211_X1 g0711(.A(KEYINPUT38), .B(new_n909), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(KEYINPUT39), .B1(new_n908), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(KEYINPUT107), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT39), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n899), .B1(new_n442), .B2(new_n434), .ZN(new_n917));
  AND3_X1   g0717(.A1(new_n434), .A2(new_n892), .A3(new_n887), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n918), .A2(new_n893), .ZN(new_n919));
  OAI21_X1  g0719(.A(KEYINPUT37), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n900), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n921), .A2(KEYINPUT108), .B1(new_n449), .B2(new_n919), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT108), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n920), .A2(new_n900), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(KEYINPUT38), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT109), .B1(new_n907), .B2(KEYINPUT38), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT109), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n912), .A2(new_n928), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n916), .B(new_n926), .C1(new_n927), .C2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT107), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n931), .B(KEYINPUT39), .C1(new_n908), .C2(new_n913), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n915), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n346), .A2(G169), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(KEYINPUT14), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n935), .A2(new_n349), .A3(new_n348), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n936), .A2(new_n334), .A3(new_n694), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n933), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n834), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n873), .A2(new_n940), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n334), .B(new_n686), .C1(new_n936), .C2(new_n670), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n334), .A2(new_n686), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n352), .A2(new_n356), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n941), .B(new_n945), .C1(new_n913), .C2(new_n908), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n437), .A2(new_n887), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n939), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n676), .A2(new_n677), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n318), .ZN(new_n951));
  INV_X1    g0751(.A(new_n755), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n952), .A2(new_n451), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n951), .B1(new_n745), .B2(new_n953), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n949), .B(new_n954), .Z(new_n955));
  NAND2_X1  g0755(.A1(new_n912), .A2(new_n928), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n904), .A2(new_n906), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n957), .A2(KEYINPUT109), .A3(KEYINPUT38), .A4(new_n909), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n925), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n945), .A2(new_n836), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n734), .A2(new_n728), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n960), .B1(new_n737), .B2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(KEYINPUT40), .B1(new_n959), .B2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT40), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n965), .B(new_n962), .C1(new_n908), .C2(new_n913), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n451), .B1(new_n737), .B2(new_n961), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n967), .A2(new_n968), .ZN(new_n971));
  NOR3_X1   g0771(.A1(new_n970), .A2(new_n971), .A3(new_n759), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n880), .B1(new_n955), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n955), .B2(new_n973), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n471), .A2(KEYINPUT35), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n471), .A2(KEYINPUT35), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n976), .A2(G116), .A3(new_n219), .A4(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT36), .ZN(new_n979));
  NOR3_X1   g0779(.A1(new_n715), .A2(new_n226), .A3(new_n419), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n223), .A2(G50), .ZN(new_n981));
  OAI211_X1 g0781(.A(G1), .B(new_n215), .C1(new_n980), .C2(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n975), .A2(new_n979), .A3(new_n982), .ZN(G367));
  OAI21_X1  g0783(.A(new_n783), .B1(new_n211), .B2(new_n567), .ZN(new_n984));
  INV_X1    g0784(.A(new_n776), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n985), .A2(new_n242), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n765), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n791), .A2(G159), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n794), .A2(new_n852), .B1(new_n798), .B2(new_n850), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n293), .B(new_n989), .C1(G50), .C2(new_n802), .ZN(new_n990));
  AOI22_X1  g0790(.A1(G68), .A2(new_n807), .B1(new_n811), .B2(G143), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n809), .A2(G58), .B1(new_n813), .B2(G77), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n988), .A2(new_n990), .A3(new_n991), .A4(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n791), .A2(G294), .ZN(new_n994));
  INV_X1    g0794(.A(G283), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n794), .A2(new_n609), .B1(new_n801), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(KEYINPUT46), .B1(new_n809), .B2(G116), .ZN(new_n997));
  AOI211_X1 g0797(.A(new_n996), .B(new_n997), .C1(G317), .C2(new_n799), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n392), .B1(G97), .B2(new_n813), .ZN(new_n999));
  XNOR2_X1  g0799(.A(KEYINPUT111), .B(G311), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n362), .A2(new_n807), .B1(new_n811), .B2(new_n1001), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n994), .A2(new_n998), .A3(new_n999), .A4(new_n1002), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n809), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT112), .Z(new_n1005));
  OAI21_X1  g0805(.A(new_n993), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT47), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n987), .B1(new_n1007), .B2(new_n782), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n770), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n573), .A2(new_n694), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n596), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n594), .B2(new_n1010), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1008), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n686), .B1(new_n648), .B2(new_n650), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n556), .A2(new_n1014), .A3(new_n504), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n644), .A2(new_n686), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n707), .A2(new_n705), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT45), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n707), .A2(KEYINPUT45), .A3(new_n705), .A4(new_n1017), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1017), .B1(new_n707), .B2(new_n705), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1023), .A2(KEYINPUT44), .ZN(new_n1024));
  AND2_X1   g0824(.A1(new_n1023), .A2(KEYINPUT44), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n703), .B(new_n1022), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1023), .B(KEYINPUT44), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n703), .B1(new_n1028), .B2(new_n1022), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n707), .B1(new_n691), .B2(new_n706), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(new_n699), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n756), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n710), .B(KEYINPUT41), .Z(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1033), .A2(KEYINPUT110), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT110), .ZN(new_n1037));
  AOI21_X1  g0837(.A(KEYINPUT29), .B1(new_n667), .B2(new_n694), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n741), .B1(new_n1038), .B2(new_n952), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1025), .A2(new_n1024), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1022), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n704), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n1026), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1032), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1039), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1037), .B1(new_n1045), .B2(new_n1034), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n764), .B1(new_n1036), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1012), .A2(KEYINPUT43), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1017), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n707), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1050), .A2(KEYINPUT42), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n504), .B1(new_n1049), .B2(new_n606), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n694), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1050), .A2(KEYINPUT42), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1048), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1012), .A2(KEYINPUT43), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1056), .B(new_n1057), .Z(new_n1058));
  NOR2_X1   g0858(.A1(new_n704), .A2(new_n1049), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1058), .B(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1013), .B1(new_n1047), .B2(new_n1060), .ZN(G387));
  NOR2_X1   g0861(.A1(new_n1039), .A2(new_n1032), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1062), .A2(new_n711), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1039), .A2(new_n1032), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  OR3_X1    g0865(.A1(new_n1032), .A2(KEYINPUT113), .A3(new_n763), .ZN(new_n1066));
  OAI21_X1  g0866(.A(KEYINPUT113), .B1(new_n1032), .B2(new_n763), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n689), .A2(new_n690), .A3(new_n770), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n713), .A2(new_n772), .B1(G107), .B2(new_n211), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n239), .A2(new_n282), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT114), .Z(new_n1071));
  AOI211_X1 g0871(.A(G45), .B(new_n712), .C1(G68), .C2(G77), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n256), .A2(G50), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT50), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n985), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1069), .B1(new_n1071), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n783), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n765), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n791), .A2(new_n257), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n808), .A2(new_n226), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n567), .A2(new_n806), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n1080), .B(new_n1081), .C1(G159), .C2(new_n811), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n801), .A2(new_n223), .B1(new_n798), .B2(new_n852), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(G50), .B2(new_n795), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n386), .B1(G97), .B2(new_n813), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1079), .A2(new_n1082), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n811), .A2(G322), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n795), .A2(G317), .B1(new_n802), .B2(G303), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1087), .B(new_n1088), .C1(new_n790), .C2(new_n1000), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT48), .ZN(new_n1090));
  OR2_X1    g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n806), .A2(new_n995), .B1(new_n808), .B2(new_n839), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1091), .A2(KEYINPUT49), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n813), .A2(G116), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n799), .A2(G326), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1094), .A2(new_n386), .A3(new_n1095), .A4(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(KEYINPUT49), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1086), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT115), .ZN(new_n1100));
  OR2_X1    g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n782), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1078), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n1066), .A2(new_n1067), .B1(new_n1068), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1065), .A2(new_n1105), .ZN(G393));
  AOI21_X1  g0906(.A(new_n711), .B1(new_n1062), .B2(new_n1043), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1030), .B1(new_n1039), .B2(new_n1032), .ZN(new_n1108));
  AND2_X1   g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  AND2_X1   g0909(.A1(new_n247), .A2(new_n776), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n783), .B1(new_n559), .B2(new_n211), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n765), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(G150), .A2(new_n811), .B1(new_n795), .B2(G159), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT51), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n808), .A2(new_n223), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n843), .B(new_n1115), .C1(G77), .C2(new_n807), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n801), .A2(new_n256), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n386), .B(new_n1117), .C1(G143), .C2(new_n799), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1116), .B(new_n1118), .C1(new_n790), .C2(new_n202), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n808), .A2(new_n995), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n816), .B(new_n1120), .C1(G116), .C2(new_n807), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n293), .B1(new_n801), .B2(new_n839), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(G322), .B2(new_n799), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1121), .B(new_n1123), .C1(new_n790), .C2(new_n609), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(G317), .A2(new_n811), .B1(new_n795), .B2(G311), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT52), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n1114), .A2(new_n1119), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1112), .B1(new_n1127), .B2(new_n782), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n1017), .B2(new_n1009), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1129), .B1(new_n1030), .B2(new_n763), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1109), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(G390));
  INV_X1    g0932(.A(KEYINPUT116), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n740), .A2(G330), .A3(new_n836), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n945), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n759), .B(new_n960), .C1(new_n737), .C2(new_n961), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n759), .B1(new_n737), .B2(new_n961), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n945), .B1(new_n1140), .B2(new_n836), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n835), .A2(new_n379), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n754), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n940), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1141), .A2(new_n1144), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n740), .A2(G330), .A3(new_n836), .A4(new_n945), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n1139), .A2(new_n941), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n452), .A2(new_n1140), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n452), .A2(new_n755), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n678), .B(new_n1148), .C1(new_n1038), .C2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1133), .B1(new_n1147), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n834), .B1(new_n754), .B2(new_n1142), .ZN(new_n1152));
  AND2_X1   g0952(.A1(new_n1140), .A2(new_n836), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1152), .B(new_n1146), .C1(new_n1153), .C2(new_n945), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1137), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n834), .B1(new_n667), .B2(new_n866), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1154), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n954), .A2(new_n1157), .A3(KEYINPUT116), .A4(new_n1148), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n926), .B1(new_n927), .B2(new_n929), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1159), .B(new_n937), .C1(new_n1135), .C2(new_n1152), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n938), .B1(new_n941), .B2(new_n945), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1160), .B(new_n1146), .C1(new_n933), .C2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n937), .B1(new_n1156), .B2(new_n1135), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1164), .A2(new_n930), .A3(new_n932), .A4(new_n915), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1138), .B1(new_n1165), .B2(new_n1160), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1151), .B(new_n1158), .C1(new_n1163), .C2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1151), .A2(new_n1158), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1160), .B1(new_n933), .B2(new_n1161), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n1137), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1168), .A2(new_n1170), .A3(new_n1162), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1167), .A2(new_n710), .A3(new_n1171), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1163), .A2(new_n1166), .ZN(new_n1173));
  OR2_X1    g0973(.A1(new_n933), .A2(new_n769), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n765), .B1(new_n861), .B2(new_n257), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n808), .A2(new_n852), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT53), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n790), .B2(new_n850), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(G159), .A2(new_n807), .B1(new_n811), .B2(G128), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n293), .B1(new_n795), .B2(G132), .ZN(new_n1180));
  XOR2_X1   g0980(.A(KEYINPUT54), .B(G143), .Z(new_n1181));
  AOI22_X1  g0981(.A1(new_n802), .A2(new_n1181), .B1(new_n799), .B2(G125), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n813), .A2(G50), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1179), .A2(new_n1180), .A3(new_n1182), .A4(new_n1183), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n790), .A2(new_n363), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(G77), .A2(new_n807), .B1(new_n811), .B2(G283), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n299), .B1(new_n799), .B2(G294), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n795), .A2(G116), .B1(new_n802), .B2(G97), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n809), .A2(G87), .B1(new_n813), .B2(G68), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .A4(new_n1189), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n1178), .A2(new_n1184), .B1(new_n1185), .B2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1175), .B1(new_n1191), .B2(new_n782), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n1173), .A2(new_n764), .B1(new_n1174), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1172), .A2(new_n1193), .ZN(G378));
  INV_X1    g0994(.A(new_n1150), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1171), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n275), .A2(new_n887), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n319), .B(new_n1197), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1198), .B(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(new_n967), .B2(G330), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n759), .B(new_n1201), .C1(new_n964), .C2(new_n966), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n949), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n966), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1159), .A2(new_n962), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1206), .B1(new_n1207), .B2(KEYINPUT40), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1201), .B1(new_n1208), .B2(new_n759), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n947), .B1(new_n933), .B2(new_n938), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n967), .A2(G330), .A3(new_n1202), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1209), .A2(new_n946), .A3(new_n1210), .A4(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1205), .A2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1196), .A2(new_n1213), .A3(KEYINPUT57), .ZN(new_n1214));
  OAI21_X1  g1014(.A(KEYINPUT120), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n949), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n949), .B(KEYINPUT120), .C1(new_n1203), .C2(new_n1204), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  AND2_X1   g1019(.A1(new_n1219), .A2(new_n1196), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n710), .B(new_n1214), .C1(new_n1220), .C2(KEYINPUT57), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n765), .B1(new_n861), .B2(G50), .ZN(new_n1222));
  AOI211_X1 g1022(.A(G33), .B(G41), .C1(new_n799), .C2(G124), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n811), .A2(G125), .B1(new_n809), .B2(new_n1181), .ZN(new_n1224));
  INV_X1    g1024(.A(G128), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1224), .B1(new_n1225), .B2(new_n794), .C1(new_n852), .C2(new_n806), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n791), .A2(G132), .B1(G137), .B2(new_n802), .ZN(new_n1227));
  OR2_X1    g1027(.A1(new_n1227), .A2(KEYINPUT118), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(KEYINPUT118), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1226), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT59), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1223), .B1(new_n822), .B2(new_n812), .C1(new_n1230), .C2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(new_n1231), .B2(new_n1230), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n386), .A2(new_n281), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1234), .A2(new_n1080), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(new_n1235), .B(KEYINPUT117), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n790), .A2(new_n559), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n795), .A2(G107), .B1(new_n802), .B2(new_n369), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1238), .B1(new_n995), .B2(new_n798), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n813), .A2(G58), .ZN(new_n1240));
  OAI221_X1 g1040(.A(new_n1240), .B1(new_n223), .B2(new_n806), .C1(new_n851), .C2(new_n616), .ZN(new_n1241));
  NOR4_X1   g1041(.A1(new_n1236), .A2(new_n1237), .A3(new_n1239), .A4(new_n1241), .ZN(new_n1242));
  OR2_X1    g1042(.A1(new_n1242), .A2(KEYINPUT58), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(KEYINPUT58), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1234), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n782), .B1(new_n1233), .B2(new_n1246), .ZN(new_n1247));
  XOR2_X1   g1047(.A(new_n1247), .B(KEYINPUT119), .Z(new_n1248));
  AOI211_X1 g1048(.A(new_n1222), .B(new_n1248), .C1(new_n1201), .C2(new_n768), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(new_n1219), .B2(new_n764), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1221), .A2(new_n1250), .ZN(G375));
  NAND2_X1  g1051(.A1(new_n1135), .A2(new_n768), .ZN(new_n1252));
  XNOR2_X1  g1052(.A(new_n1252), .B(KEYINPUT121), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n765), .B1(new_n861), .B2(G68), .ZN(new_n1254));
  OAI221_X1 g1054(.A(new_n1240), .B1(new_n822), .B2(new_n808), .C1(new_n202), .C2(new_n806), .ZN(new_n1255));
  OAI22_X1  g1055(.A1(new_n801), .A2(new_n852), .B1(new_n798), .B2(new_n1225), .ZN(new_n1256));
  NOR3_X1   g1056(.A1(new_n1255), .A2(new_n386), .A3(new_n1256), .ZN(new_n1257));
  XOR2_X1   g1057(.A(new_n1257), .B(KEYINPUT123), .Z(new_n1258));
  NAND2_X1  g1058(.A1(new_n791), .A2(new_n1181), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(G132), .A2(new_n811), .B1(new_n795), .B2(G137), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n293), .B1(new_n812), .B2(new_n226), .ZN(new_n1262));
  XOR2_X1   g1062(.A(new_n1262), .B(KEYINPUT122), .Z(new_n1263));
  NOR2_X1   g1063(.A1(new_n808), .A2(new_n559), .ZN(new_n1264));
  AOI211_X1 g1064(.A(new_n1264), .B(new_n1081), .C1(G294), .C2(new_n811), .ZN(new_n1265));
  OAI22_X1  g1065(.A1(new_n363), .A2(new_n801), .B1(new_n794), .B2(new_n995), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1266), .B1(G303), .B2(new_n799), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1265), .B(new_n1267), .C1(new_n616), .C2(new_n790), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n1258), .A2(new_n1261), .B1(new_n1263), .B2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1254), .B1(new_n1269), .B2(new_n782), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(new_n1157), .A2(new_n764), .B1(new_n1253), .B2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1151), .A2(new_n1158), .A3(new_n1272), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1271), .B1(new_n1273), .B2(new_n1034), .ZN(G381));
  NAND3_X1  g1074(.A1(new_n1065), .A2(new_n832), .A3(new_n1105), .ZN(new_n1275));
  OR4_X1    g1075(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1275), .ZN(new_n1276));
  OR4_X1    g1076(.A1(G387), .A2(G375), .A3(G378), .A4(new_n1276), .ZN(G407));
  INV_X1    g1077(.A(G378), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n685), .A2(G213), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1278), .A2(new_n1280), .ZN(new_n1281));
  OAI211_X1 g1081(.A(G407), .B(G213), .C1(G375), .C2(new_n1281), .ZN(G409));
  NOR3_X1   g1082(.A1(new_n949), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1283));
  AOI22_X1  g1083(.A1(new_n1209), .A2(new_n1211), .B1(new_n1210), .B2(new_n946), .ZN(new_n1284));
  OAI21_X1  g1084(.A(KEYINPUT57), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1150), .B1(new_n1173), .B2(new_n1168), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n710), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(KEYINPUT57), .B1(new_n1219), .B2(new_n1196), .ZN(new_n1288));
  OAI211_X1 g1088(.A(G378), .B(new_n1250), .C1(new_n1287), .C2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1219), .A2(new_n1035), .A3(new_n1196), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1249), .B1(new_n1213), .B2(new_n764), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(new_n1278), .ZN(new_n1293));
  AND2_X1   g1093(.A1(new_n1289), .A2(new_n1293), .ZN(new_n1294));
  OAI21_X1  g1094(.A(KEYINPUT124), .B1(new_n1294), .B2(new_n1280), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1273), .A2(KEYINPUT60), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT60), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n711), .B1(new_n1272), .B2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1296), .A2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n1271), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n878), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1299), .A2(G384), .A3(new_n1271), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1280), .A2(G2897), .ZN(new_n1303));
  XOR2_X1   g1103(.A(new_n1303), .B(KEYINPUT125), .Z(new_n1304));
  AND3_X1   g1104(.A1(new_n1301), .A2(new_n1302), .A3(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1304), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1280), .B1(new_n1289), .B2(new_n1293), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT124), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1307), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1295), .A2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1308), .A2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT63), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT126), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(G393), .A2(G396), .ZN(new_n1318));
  AND2_X1   g1118(.A1(new_n1318), .A2(new_n1275), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1036), .A2(new_n1046), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(new_n763), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1060), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1131), .B1(new_n1323), .B2(new_n1013), .ZN(new_n1324));
  OAI211_X1 g1124(.A(new_n1131), .B(new_n1013), .C1(new_n1047), .C2(new_n1060), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1325), .ZN(new_n1326));
  OAI211_X1 g1126(.A(new_n1317), .B(new_n1319), .C1(new_n1324), .C2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT61), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1317), .B1(new_n1318), .B2(new_n1275), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1329), .B1(G387), .B2(G390), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1319), .A2(new_n1317), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1330), .A2(new_n1331), .A3(new_n1325), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1327), .A2(new_n1328), .A3(new_n1332), .ZN(new_n1333));
  AOI211_X1 g1133(.A(new_n1280), .B(new_n1312), .C1(new_n1289), .C2(new_n1293), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1333), .B1(new_n1334), .B2(KEYINPUT63), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1311), .A2(new_n1316), .A3(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT62), .ZN(new_n1337));
  AND3_X1   g1137(.A1(new_n1308), .A2(new_n1337), .A3(new_n1313), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1328), .B1(new_n1308), .B2(new_n1307), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1337), .B1(new_n1308), .B2(new_n1313), .ZN(new_n1340));
  NOR3_X1   g1140(.A1(new_n1338), .A2(new_n1339), .A3(new_n1340), .ZN(new_n1341));
  AND3_X1   g1141(.A1(new_n1330), .A2(new_n1331), .A3(new_n1325), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1331), .B1(new_n1330), .B2(new_n1325), .ZN(new_n1343));
  NOR2_X1   g1143(.A1(new_n1342), .A2(new_n1343), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1336), .B1(new_n1341), .B2(new_n1344), .ZN(G405));
  NAND2_X1  g1145(.A1(G375), .A2(new_n1278), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1346), .A2(new_n1289), .A3(new_n1312), .ZN(new_n1347));
  AOI21_X1  g1147(.A(G378), .B1(new_n1221), .B2(new_n1250), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1289), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1313), .B1(new_n1348), .B2(new_n1349), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1347), .A2(new_n1350), .ZN(new_n1351));
  INV_X1    g1151(.A(KEYINPUT127), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1352), .B1(new_n1342), .B2(new_n1343), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1327), .A2(KEYINPUT127), .A3(new_n1332), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1353), .A2(new_n1354), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1351), .A2(new_n1355), .ZN(new_n1356));
  NAND4_X1  g1156(.A1(new_n1347), .A2(new_n1350), .A3(new_n1353), .A4(new_n1354), .ZN(new_n1357));
  AND2_X1   g1157(.A1(new_n1356), .A2(new_n1357), .ZN(G402));
endmodule


