

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X2 U548 ( .A1(n520), .A2(G2105), .ZN(n871) );
  INV_X1 U549 ( .A(G2104), .ZN(n520) );
  XNOR2_X1 U550 ( .A(n586), .B(KEYINPUT15), .ZN(n976) );
  XNOR2_X2 U551 ( .A(n685), .B(n684), .ZN(n687) );
  NAND2_X1 U552 ( .A1(n680), .A2(G40), .ZN(n771) );
  AND2_X2 U553 ( .A1(G2104), .A2(G2105), .ZN(n872) );
  NOR2_X2 U554 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X2 U555 ( .A(n689), .B(n688), .ZN(n703) );
  AND2_X2 U556 ( .A1(n533), .A2(G137), .ZN(n516) );
  XNOR2_X1 U557 ( .A(n771), .B(n681), .ZN(n682) );
  AND2_X1 U558 ( .A1(n769), .A2(n768), .ZN(n514) );
  AND2_X1 U559 ( .A1(n517), .A2(n804), .ZN(n515) );
  AND2_X1 U560 ( .A1(n785), .A2(n811), .ZN(n517) );
  INV_X1 U561 ( .A(KEYINPUT27), .ZN(n684) );
  XNOR2_X1 U562 ( .A(n727), .B(KEYINPUT94), .ZN(n741) );
  XNOR2_X1 U563 ( .A(n737), .B(KEYINPUT32), .ZN(n747) );
  NOR2_X1 U564 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U565 ( .A1(n682), .A2(n772), .ZN(n716) );
  NOR2_X1 U566 ( .A1(G164), .A2(G1384), .ZN(n772) );
  INV_X1 U567 ( .A(KEYINPUT17), .ZN(n526) );
  INV_X1 U568 ( .A(KEYINPUT64), .ZN(n523) );
  NOR2_X1 U569 ( .A1(G651), .A2(n633), .ZN(n639) );
  XNOR2_X1 U570 ( .A(n524), .B(n523), .ZN(n530) );
  BUF_X1 U571 ( .A(n680), .Z(G160) );
  NOR2_X2 U572 ( .A1(G2105), .A2(n520), .ZN(n531) );
  NAND2_X1 U573 ( .A1(n531), .A2(G101), .ZN(n519) );
  INV_X1 U574 ( .A(KEYINPUT23), .ZN(n518) );
  XNOR2_X1 U575 ( .A(n519), .B(n518), .ZN(n522) );
  NAND2_X1 U576 ( .A1(n871), .A2(G125), .ZN(n521) );
  NAND2_X1 U577 ( .A1(n522), .A2(n521), .ZN(n524) );
  NAND2_X1 U578 ( .A1(G113), .A2(n872), .ZN(n525) );
  XNOR2_X1 U579 ( .A(KEYINPUT65), .B(n525), .ZN(n528) );
  NOR2_X2 U580 ( .A1(G2104), .A2(G2105), .ZN(n527) );
  XNOR2_X2 U581 ( .A(n527), .B(n526), .ZN(n533) );
  NOR2_X1 U582 ( .A1(n528), .A2(n516), .ZN(n529) );
  AND2_X2 U583 ( .A1(n530), .A2(n529), .ZN(n680) );
  INV_X1 U584 ( .A(n531), .ZN(n532) );
  INV_X1 U585 ( .A(n532), .ZN(n868) );
  NAND2_X1 U586 ( .A1(G102), .A2(n868), .ZN(n535) );
  NAND2_X1 U587 ( .A1(G138), .A2(n533), .ZN(n534) );
  NAND2_X1 U588 ( .A1(n535), .A2(n534), .ZN(n539) );
  NAND2_X1 U589 ( .A1(G126), .A2(n871), .ZN(n537) );
  NAND2_X1 U590 ( .A1(G114), .A2(n872), .ZN(n536) );
  NAND2_X1 U591 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U592 ( .A1(n539), .A2(n538), .ZN(G164) );
  XOR2_X1 U593 ( .A(KEYINPUT0), .B(G543), .Z(n633) );
  NAND2_X1 U594 ( .A1(n639), .A2(G47), .ZN(n543) );
  XOR2_X1 U595 ( .A(KEYINPUT66), .B(G651), .Z(n544) );
  NOR2_X1 U596 ( .A1(G543), .A2(n544), .ZN(n540) );
  XNOR2_X1 U597 ( .A(n540), .B(KEYINPUT67), .ZN(n541) );
  XNOR2_X2 U598 ( .A(KEYINPUT1), .B(n541), .ZN(n642) );
  NAND2_X1 U599 ( .A1(G60), .A2(n642), .ZN(n542) );
  NAND2_X1 U600 ( .A1(n543), .A2(n542), .ZN(n548) );
  NOR2_X1 U601 ( .A1(G651), .A2(G543), .ZN(n645) );
  NAND2_X1 U602 ( .A1(n645), .A2(G85), .ZN(n546) );
  NOR2_X1 U603 ( .A1(n633), .A2(n544), .ZN(n641) );
  NAND2_X1 U604 ( .A1(G72), .A2(n641), .ZN(n545) );
  NAND2_X1 U605 ( .A1(n546), .A2(n545), .ZN(n547) );
  OR2_X1 U606 ( .A1(n548), .A2(n547), .ZN(G290) );
  NAND2_X1 U607 ( .A1(n639), .A2(G52), .ZN(n550) );
  NAND2_X1 U608 ( .A1(G64), .A2(n642), .ZN(n549) );
  NAND2_X1 U609 ( .A1(n550), .A2(n549), .ZN(n556) );
  NAND2_X1 U610 ( .A1(G77), .A2(n641), .ZN(n551) );
  XNOR2_X1 U611 ( .A(n551), .B(KEYINPUT68), .ZN(n553) );
  NAND2_X1 U612 ( .A1(G90), .A2(n645), .ZN(n552) );
  NAND2_X1 U613 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U614 ( .A(KEYINPUT9), .B(n554), .Z(n555) );
  NOR2_X1 U615 ( .A1(n556), .A2(n555), .ZN(G171) );
  INV_X1 U616 ( .A(G171), .ZN(G301) );
  AND2_X1 U617 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U618 ( .A(G57), .ZN(G237) );
  NAND2_X1 U619 ( .A1(n645), .A2(G89), .ZN(n557) );
  XNOR2_X1 U620 ( .A(n557), .B(KEYINPUT4), .ZN(n559) );
  NAND2_X1 U621 ( .A1(G76), .A2(n641), .ZN(n558) );
  NAND2_X1 U622 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U623 ( .A(n560), .B(KEYINPUT5), .ZN(n565) );
  NAND2_X1 U624 ( .A1(n639), .A2(G51), .ZN(n562) );
  NAND2_X1 U625 ( .A1(G63), .A2(n642), .ZN(n561) );
  NAND2_X1 U626 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U627 ( .A(KEYINPUT6), .B(n563), .Z(n564) );
  NAND2_X1 U628 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U629 ( .A(n566), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U630 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U631 ( .A1(G7), .A2(G661), .ZN(n567) );
  XNOR2_X1 U632 ( .A(n567), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U633 ( .A(G223), .ZN(n821) );
  NAND2_X1 U634 ( .A1(n821), .A2(G567), .ZN(n568) );
  XOR2_X1 U635 ( .A(KEYINPUT11), .B(n568), .Z(G234) );
  XOR2_X1 U636 ( .A(KEYINPUT69), .B(KEYINPUT14), .Z(n570) );
  NAND2_X1 U637 ( .A1(G56), .A2(n642), .ZN(n569) );
  XNOR2_X1 U638 ( .A(n570), .B(n569), .ZN(n579) );
  NAND2_X1 U639 ( .A1(G43), .A2(n639), .ZN(n571) );
  XOR2_X1 U640 ( .A(KEYINPUT70), .B(n571), .Z(n577) );
  NAND2_X1 U641 ( .A1(n645), .A2(G81), .ZN(n572) );
  XNOR2_X1 U642 ( .A(n572), .B(KEYINPUT12), .ZN(n574) );
  NAND2_X1 U643 ( .A1(G68), .A2(n641), .ZN(n573) );
  NAND2_X1 U644 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U645 ( .A(KEYINPUT13), .B(n575), .Z(n576) );
  NOR2_X1 U646 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U647 ( .A1(n579), .A2(n578), .ZN(n981) );
  INV_X1 U648 ( .A(G860), .ZN(n598) );
  OR2_X1 U649 ( .A1(n981), .A2(n598), .ZN(G153) );
  NAND2_X1 U650 ( .A1(G868), .A2(G301), .ZN(n588) );
  NAND2_X1 U651 ( .A1(n645), .A2(G92), .ZN(n581) );
  NAND2_X1 U652 ( .A1(G79), .A2(n641), .ZN(n580) );
  NAND2_X1 U653 ( .A1(n581), .A2(n580), .ZN(n585) );
  NAND2_X1 U654 ( .A1(n639), .A2(G54), .ZN(n583) );
  NAND2_X1 U655 ( .A1(G66), .A2(n642), .ZN(n582) );
  NAND2_X1 U656 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U657 ( .A1(n585), .A2(n584), .ZN(n586) );
  INV_X1 U658 ( .A(G868), .ZN(n661) );
  NAND2_X1 U659 ( .A1(n976), .A2(n661), .ZN(n587) );
  NAND2_X1 U660 ( .A1(n588), .A2(n587), .ZN(G284) );
  NAND2_X1 U661 ( .A1(n639), .A2(G53), .ZN(n590) );
  NAND2_X1 U662 ( .A1(G65), .A2(n642), .ZN(n589) );
  NAND2_X1 U663 ( .A1(n590), .A2(n589), .ZN(n594) );
  NAND2_X1 U664 ( .A1(n645), .A2(G91), .ZN(n592) );
  NAND2_X1 U665 ( .A1(G78), .A2(n641), .ZN(n591) );
  NAND2_X1 U666 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U667 ( .A1(n594), .A2(n593), .ZN(n704) );
  INV_X1 U668 ( .A(n704), .ZN(G299) );
  NOR2_X1 U669 ( .A1(G286), .A2(n661), .ZN(n596) );
  NOR2_X1 U670 ( .A1(G868), .A2(G299), .ZN(n595) );
  NOR2_X1 U671 ( .A1(n596), .A2(n595), .ZN(n597) );
  XOR2_X1 U672 ( .A(KEYINPUT71), .B(n597), .Z(G297) );
  NAND2_X1 U673 ( .A1(n598), .A2(G559), .ZN(n599) );
  INV_X1 U674 ( .A(n976), .ZN(n621) );
  NAND2_X1 U675 ( .A1(n599), .A2(n621), .ZN(n600) );
  XNOR2_X1 U676 ( .A(n600), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U677 ( .A1(G868), .A2(n981), .ZN(n603) );
  NAND2_X1 U678 ( .A1(G868), .A2(n621), .ZN(n601) );
  NOR2_X1 U679 ( .A1(G559), .A2(n601), .ZN(n602) );
  NOR2_X1 U680 ( .A1(n603), .A2(n602), .ZN(G282) );
  NAND2_X1 U681 ( .A1(G123), .A2(n871), .ZN(n604) );
  XNOR2_X1 U682 ( .A(n604), .B(KEYINPUT18), .ZN(n607) );
  NAND2_X1 U683 ( .A1(G99), .A2(n868), .ZN(n605) );
  XNOR2_X1 U684 ( .A(n605), .B(KEYINPUT72), .ZN(n606) );
  NAND2_X1 U685 ( .A1(n607), .A2(n606), .ZN(n611) );
  NAND2_X1 U686 ( .A1(G111), .A2(n872), .ZN(n609) );
  NAND2_X1 U687 ( .A1(G135), .A2(n533), .ZN(n608) );
  NAND2_X1 U688 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U689 ( .A1(n611), .A2(n610), .ZN(n938) );
  XNOR2_X1 U690 ( .A(n938), .B(G2096), .ZN(n613) );
  INV_X1 U691 ( .A(G2100), .ZN(n612) );
  NAND2_X1 U692 ( .A1(n613), .A2(n612), .ZN(G156) );
  NAND2_X1 U693 ( .A1(n645), .A2(G93), .ZN(n615) );
  NAND2_X1 U694 ( .A1(G67), .A2(n642), .ZN(n614) );
  NAND2_X1 U695 ( .A1(n615), .A2(n614), .ZN(n618) );
  NAND2_X1 U696 ( .A1(G55), .A2(n639), .ZN(n616) );
  XNOR2_X1 U697 ( .A(KEYINPUT73), .B(n616), .ZN(n617) );
  NOR2_X1 U698 ( .A1(n618), .A2(n617), .ZN(n620) );
  NAND2_X1 U699 ( .A1(G80), .A2(n641), .ZN(n619) );
  NAND2_X1 U700 ( .A1(n620), .A2(n619), .ZN(n662) );
  NAND2_X1 U701 ( .A1(n621), .A2(G559), .ZN(n659) );
  XNOR2_X1 U702 ( .A(n981), .B(n659), .ZN(n622) );
  NOR2_X1 U703 ( .A1(G860), .A2(n622), .ZN(n623) );
  XOR2_X1 U704 ( .A(n662), .B(n623), .Z(G145) );
  NAND2_X1 U705 ( .A1(n641), .A2(G73), .ZN(n624) );
  XNOR2_X1 U706 ( .A(n624), .B(KEYINPUT2), .ZN(n631) );
  NAND2_X1 U707 ( .A1(n645), .A2(G86), .ZN(n626) );
  NAND2_X1 U708 ( .A1(G61), .A2(n642), .ZN(n625) );
  NAND2_X1 U709 ( .A1(n626), .A2(n625), .ZN(n629) );
  NAND2_X1 U710 ( .A1(n639), .A2(G48), .ZN(n627) );
  XOR2_X1 U711 ( .A(KEYINPUT74), .B(n627), .Z(n628) );
  NOR2_X1 U712 ( .A1(n629), .A2(n628), .ZN(n630) );
  NAND2_X1 U713 ( .A1(n631), .A2(n630), .ZN(n632) );
  XOR2_X1 U714 ( .A(KEYINPUT75), .B(n632), .Z(G305) );
  NAND2_X1 U715 ( .A1(G87), .A2(n633), .ZN(n635) );
  NAND2_X1 U716 ( .A1(G74), .A2(G651), .ZN(n634) );
  NAND2_X1 U717 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U718 ( .A1(n642), .A2(n636), .ZN(n638) );
  NAND2_X1 U719 ( .A1(n639), .A2(G49), .ZN(n637) );
  NAND2_X1 U720 ( .A1(n638), .A2(n637), .ZN(G288) );
  NAND2_X1 U721 ( .A1(G50), .A2(n639), .ZN(n640) );
  XNOR2_X1 U722 ( .A(n640), .B(KEYINPUT76), .ZN(n650) );
  NAND2_X1 U723 ( .A1(G75), .A2(n641), .ZN(n644) );
  NAND2_X1 U724 ( .A1(G62), .A2(n642), .ZN(n643) );
  NAND2_X1 U725 ( .A1(n644), .A2(n643), .ZN(n648) );
  NAND2_X1 U726 ( .A1(G88), .A2(n645), .ZN(n646) );
  XNOR2_X1 U727 ( .A(KEYINPUT77), .B(n646), .ZN(n647) );
  NOR2_X1 U728 ( .A1(n648), .A2(n647), .ZN(n649) );
  NAND2_X1 U729 ( .A1(n650), .A2(n649), .ZN(G303) );
  XNOR2_X1 U730 ( .A(n981), .B(G305), .ZN(n658) );
  XNOR2_X1 U731 ( .A(KEYINPUT19), .B(KEYINPUT79), .ZN(n652) );
  XNOR2_X1 U732 ( .A(G288), .B(KEYINPUT78), .ZN(n651) );
  XNOR2_X1 U733 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U734 ( .A(n653), .B(G303), .ZN(n654) );
  XNOR2_X1 U735 ( .A(n654), .B(n662), .ZN(n655) );
  XNOR2_X1 U736 ( .A(n704), .B(n655), .ZN(n656) );
  XNOR2_X1 U737 ( .A(n656), .B(G290), .ZN(n657) );
  XNOR2_X1 U738 ( .A(n658), .B(n657), .ZN(n892) );
  XOR2_X1 U739 ( .A(n892), .B(n659), .Z(n660) );
  NOR2_X1 U740 ( .A1(n661), .A2(n660), .ZN(n664) );
  NOR2_X1 U741 ( .A1(G868), .A2(n662), .ZN(n663) );
  NOR2_X1 U742 ( .A1(n664), .A2(n663), .ZN(G295) );
  NAND2_X1 U743 ( .A1(G2078), .A2(G2084), .ZN(n665) );
  XOR2_X1 U744 ( .A(KEYINPUT20), .B(n665), .Z(n666) );
  NAND2_X1 U745 ( .A1(G2090), .A2(n666), .ZN(n667) );
  XNOR2_X1 U746 ( .A(KEYINPUT21), .B(n667), .ZN(n668) );
  NAND2_X1 U747 ( .A1(n668), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U748 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U749 ( .A1(G132), .A2(G82), .ZN(n669) );
  XNOR2_X1 U750 ( .A(n669), .B(KEYINPUT80), .ZN(n670) );
  XNOR2_X1 U751 ( .A(n670), .B(KEYINPUT22), .ZN(n671) );
  NOR2_X1 U752 ( .A1(G218), .A2(n671), .ZN(n672) );
  NAND2_X1 U753 ( .A1(G96), .A2(n672), .ZN(n826) );
  NAND2_X1 U754 ( .A1(G2106), .A2(n826), .ZN(n676) );
  NAND2_X1 U755 ( .A1(G108), .A2(G120), .ZN(n673) );
  NOR2_X1 U756 ( .A1(G237), .A2(n673), .ZN(n674) );
  NAND2_X1 U757 ( .A1(G69), .A2(n674), .ZN(n827) );
  NAND2_X1 U758 ( .A1(G567), .A2(n827), .ZN(n675) );
  NAND2_X1 U759 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U760 ( .A(KEYINPUT81), .B(n677), .ZN(G319) );
  INV_X1 U761 ( .A(G319), .ZN(n679) );
  NAND2_X1 U762 ( .A1(G661), .A2(G483), .ZN(n678) );
  NOR2_X1 U763 ( .A1(n679), .A2(n678), .ZN(n825) );
  NAND2_X1 U764 ( .A1(n825), .A2(G36), .ZN(G176) );
  INV_X1 U765 ( .A(G303), .ZN(G166) );
  INV_X1 U766 ( .A(KEYINPUT88), .ZN(n681) );
  BUF_X2 U767 ( .A(n716), .Z(n729) );
  NAND2_X1 U768 ( .A1(G8), .A2(n729), .ZN(n766) );
  INV_X1 U769 ( .A(G2072), .ZN(n683) );
  OR2_X2 U770 ( .A1(n716), .A2(n683), .ZN(n685) );
  NAND2_X1 U771 ( .A1(G1956), .A2(n729), .ZN(n686) );
  NAND2_X1 U772 ( .A1(n687), .A2(n686), .ZN(n689) );
  INV_X1 U773 ( .A(KEYINPUT92), .ZN(n688) );
  NOR2_X2 U774 ( .A1(n704), .A2(n703), .ZN(n691) );
  INV_X1 U775 ( .A(KEYINPUT28), .ZN(n690) );
  XNOR2_X1 U776 ( .A(n691), .B(n690), .ZN(n708) );
  INV_X1 U777 ( .A(G1996), .ZN(n993) );
  NOR2_X1 U778 ( .A1(n716), .A2(n993), .ZN(n692) );
  XOR2_X1 U779 ( .A(n692), .B(KEYINPUT26), .Z(n694) );
  NAND2_X1 U780 ( .A1(n729), .A2(G1341), .ZN(n693) );
  NAND2_X1 U781 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U782 ( .A1(n981), .A2(n695), .ZN(n699) );
  NAND2_X1 U783 ( .A1(G1348), .A2(n729), .ZN(n697) );
  INV_X1 U784 ( .A(n729), .ZN(n710) );
  NAND2_X1 U785 ( .A1(G2067), .A2(n710), .ZN(n696) );
  NAND2_X1 U786 ( .A1(n697), .A2(n696), .ZN(n700) );
  NOR2_X1 U787 ( .A1(n976), .A2(n700), .ZN(n698) );
  OR2_X1 U788 ( .A1(n699), .A2(n698), .ZN(n702) );
  NAND2_X1 U789 ( .A1(n976), .A2(n700), .ZN(n701) );
  NAND2_X1 U790 ( .A1(n702), .A2(n701), .ZN(n706) );
  NAND2_X1 U791 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U792 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U793 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U794 ( .A(n709), .B(KEYINPUT29), .ZN(n714) );
  XNOR2_X1 U795 ( .A(G2078), .B(KEYINPUT25), .ZN(n992) );
  NOR2_X1 U796 ( .A1(n729), .A2(n992), .ZN(n712) );
  INV_X1 U797 ( .A(G1961), .ZN(n912) );
  NOR2_X1 U798 ( .A1(n710), .A2(n912), .ZN(n711) );
  NOR2_X1 U799 ( .A1(n712), .A2(n711), .ZN(n721) );
  AND2_X1 U800 ( .A1(G171), .A2(n721), .ZN(n713) );
  XNOR2_X1 U801 ( .A(n715), .B(KEYINPUT93), .ZN(n726) );
  NOR2_X1 U802 ( .A1(G1966), .A2(n766), .ZN(n745) );
  NOR2_X1 U803 ( .A1(G2084), .A2(n716), .ZN(n717) );
  XOR2_X1 U804 ( .A(KEYINPUT90), .B(n717), .Z(n738) );
  NAND2_X1 U805 ( .A1(G8), .A2(n738), .ZN(n718) );
  NOR2_X1 U806 ( .A1(n745), .A2(n718), .ZN(n719) );
  XOR2_X1 U807 ( .A(KEYINPUT30), .B(n719), .Z(n720) );
  NOR2_X1 U808 ( .A1(G168), .A2(n720), .ZN(n723) );
  NOR2_X1 U809 ( .A1(G171), .A2(n721), .ZN(n722) );
  NOR2_X1 U810 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U811 ( .A(KEYINPUT31), .B(n724), .Z(n725) );
  NAND2_X1 U812 ( .A1(n726), .A2(n725), .ZN(n727) );
  AND2_X1 U813 ( .A1(G286), .A2(G8), .ZN(n728) );
  NAND2_X1 U814 ( .A1(n741), .A2(n728), .ZN(n736) );
  INV_X1 U815 ( .A(G8), .ZN(n734) );
  NOR2_X1 U816 ( .A1(G1971), .A2(n766), .ZN(n731) );
  NOR2_X1 U817 ( .A1(G2090), .A2(n729), .ZN(n730) );
  NOR2_X1 U818 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U819 ( .A1(n732), .A2(G303), .ZN(n733) );
  OR2_X1 U820 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U821 ( .A1(n736), .A2(n735), .ZN(n737) );
  INV_X1 U822 ( .A(n738), .ZN(n739) );
  NAND2_X1 U823 ( .A1(G8), .A2(n739), .ZN(n740) );
  XOR2_X1 U824 ( .A(KEYINPUT91), .B(n740), .Z(n743) );
  BUF_X1 U825 ( .A(n741), .Z(n742) );
  NAND2_X1 U826 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U827 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U828 ( .A(n748), .B(KEYINPUT95), .ZN(n761) );
  NOR2_X1 U829 ( .A1(G1976), .A2(G288), .ZN(n754) );
  NOR2_X1 U830 ( .A1(G1971), .A2(G303), .ZN(n749) );
  NOR2_X1 U831 ( .A1(n754), .A2(n749), .ZN(n973) );
  NAND2_X1 U832 ( .A1(n761), .A2(n973), .ZN(n750) );
  NAND2_X1 U833 ( .A1(G1976), .A2(G288), .ZN(n969) );
  NAND2_X1 U834 ( .A1(n750), .A2(n969), .ZN(n751) );
  XNOR2_X1 U835 ( .A(KEYINPUT96), .B(n751), .ZN(n752) );
  NOR2_X1 U836 ( .A1(n766), .A2(n752), .ZN(n753) );
  NOR2_X1 U837 ( .A1(KEYINPUT33), .A2(n753), .ZN(n757) );
  NAND2_X1 U838 ( .A1(n754), .A2(KEYINPUT33), .ZN(n755) );
  NOR2_X1 U839 ( .A1(n766), .A2(n755), .ZN(n756) );
  NOR2_X1 U840 ( .A1(n757), .A2(n756), .ZN(n758) );
  XOR2_X1 U841 ( .A(G1981), .B(G305), .Z(n964) );
  NAND2_X1 U842 ( .A1(n758), .A2(n964), .ZN(n770) );
  NAND2_X1 U843 ( .A1(G8), .A2(G166), .ZN(n759) );
  NOR2_X1 U844 ( .A1(G2090), .A2(n759), .ZN(n760) );
  XNOR2_X1 U845 ( .A(n760), .B(KEYINPUT97), .ZN(n762) );
  NAND2_X1 U846 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U847 ( .A1(n763), .A2(n766), .ZN(n769) );
  NOR2_X1 U848 ( .A1(G1981), .A2(G305), .ZN(n764) );
  XNOR2_X1 U849 ( .A(n764), .B(KEYINPUT89), .ZN(n765) );
  XNOR2_X1 U850 ( .A(n765), .B(KEYINPUT24), .ZN(n767) );
  OR2_X1 U851 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U852 ( .A1(n770), .A2(n514), .ZN(n803) );
  NOR2_X1 U853 ( .A1(n772), .A2(n771), .ZN(n816) );
  XNOR2_X1 U854 ( .A(G1986), .B(G290), .ZN(n975) );
  NAND2_X1 U855 ( .A1(n816), .A2(n975), .ZN(n773) );
  XNOR2_X1 U856 ( .A(n773), .B(KEYINPUT82), .ZN(n785) );
  XNOR2_X1 U857 ( .A(KEYINPUT37), .B(G2067), .ZN(n813) );
  NAND2_X1 U858 ( .A1(G104), .A2(n868), .ZN(n775) );
  NAND2_X1 U859 ( .A1(G140), .A2(n533), .ZN(n774) );
  NAND2_X1 U860 ( .A1(n775), .A2(n774), .ZN(n777) );
  XOR2_X1 U861 ( .A(KEYINPUT83), .B(KEYINPUT34), .Z(n776) );
  XNOR2_X1 U862 ( .A(n777), .B(n776), .ZN(n783) );
  NAND2_X1 U863 ( .A1(n872), .A2(G116), .ZN(n778) );
  XNOR2_X1 U864 ( .A(n778), .B(KEYINPUT84), .ZN(n780) );
  NAND2_X1 U865 ( .A1(G128), .A2(n871), .ZN(n779) );
  NAND2_X1 U866 ( .A1(n780), .A2(n779), .ZN(n781) );
  XOR2_X1 U867 ( .A(KEYINPUT35), .B(n781), .Z(n782) );
  NOR2_X1 U868 ( .A1(n783), .A2(n782), .ZN(n784) );
  XNOR2_X1 U869 ( .A(KEYINPUT36), .B(n784), .ZN(n889) );
  NOR2_X1 U870 ( .A1(n813), .A2(n889), .ZN(n940) );
  NAND2_X1 U871 ( .A1(n816), .A2(n940), .ZN(n811) );
  NAND2_X1 U872 ( .A1(G119), .A2(n871), .ZN(n787) );
  NAND2_X1 U873 ( .A1(G131), .A2(n533), .ZN(n786) );
  NAND2_X1 U874 ( .A1(n787), .A2(n786), .ZN(n791) );
  NAND2_X1 U875 ( .A1(G95), .A2(n868), .ZN(n789) );
  NAND2_X1 U876 ( .A1(G107), .A2(n872), .ZN(n788) );
  NAND2_X1 U877 ( .A1(n789), .A2(n788), .ZN(n790) );
  NOR2_X1 U878 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U879 ( .A(n792), .B(KEYINPUT85), .ZN(n866) );
  XNOR2_X1 U880 ( .A(KEYINPUT86), .B(G1991), .ZN(n1004) );
  NAND2_X1 U881 ( .A1(n866), .A2(n1004), .ZN(n801) );
  NAND2_X1 U882 ( .A1(G129), .A2(n871), .ZN(n794) );
  NAND2_X1 U883 ( .A1(G141), .A2(n533), .ZN(n793) );
  NAND2_X1 U884 ( .A1(n794), .A2(n793), .ZN(n797) );
  NAND2_X1 U885 ( .A1(G105), .A2(n868), .ZN(n795) );
  XOR2_X1 U886 ( .A(KEYINPUT38), .B(n795), .Z(n796) );
  NOR2_X1 U887 ( .A1(n797), .A2(n796), .ZN(n799) );
  NAND2_X1 U888 ( .A1(n872), .A2(G117), .ZN(n798) );
  NAND2_X1 U889 ( .A1(n799), .A2(n798), .ZN(n865) );
  NAND2_X1 U890 ( .A1(G1996), .A2(n865), .ZN(n800) );
  NAND2_X1 U891 ( .A1(n801), .A2(n800), .ZN(n802) );
  XOR2_X1 U892 ( .A(KEYINPUT87), .B(n802), .Z(n944) );
  NAND2_X1 U893 ( .A1(n816), .A2(n944), .ZN(n804) );
  NAND2_X1 U894 ( .A1(n803), .A2(n515), .ZN(n819) );
  NOR2_X1 U895 ( .A1(G1996), .A2(n865), .ZN(n949) );
  INV_X1 U896 ( .A(n804), .ZN(n808) );
  NOR2_X1 U897 ( .A1(G1986), .A2(G290), .ZN(n806) );
  NOR2_X1 U898 ( .A1(n1004), .A2(n866), .ZN(n805) );
  XNOR2_X1 U899 ( .A(KEYINPUT98), .B(n805), .ZN(n937) );
  NOR2_X1 U900 ( .A1(n806), .A2(n937), .ZN(n807) );
  NOR2_X1 U901 ( .A1(n808), .A2(n807), .ZN(n809) );
  NOR2_X1 U902 ( .A1(n949), .A2(n809), .ZN(n810) );
  XNOR2_X1 U903 ( .A(n810), .B(KEYINPUT39), .ZN(n812) );
  NAND2_X1 U904 ( .A1(n812), .A2(n811), .ZN(n814) );
  NAND2_X1 U905 ( .A1(n813), .A2(n889), .ZN(n946) );
  NAND2_X1 U906 ( .A1(n814), .A2(n946), .ZN(n815) );
  NAND2_X1 U907 ( .A1(n816), .A2(n815), .ZN(n817) );
  XOR2_X1 U908 ( .A(KEYINPUT99), .B(n817), .Z(n818) );
  NAND2_X1 U909 ( .A1(n819), .A2(n818), .ZN(n820) );
  XNOR2_X1 U910 ( .A(n820), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U911 ( .A1(G2106), .A2(n821), .ZN(G217) );
  AND2_X1 U912 ( .A1(G15), .A2(G2), .ZN(n822) );
  NAND2_X1 U913 ( .A1(G661), .A2(n822), .ZN(G259) );
  NAND2_X1 U914 ( .A1(G3), .A2(G1), .ZN(n823) );
  XOR2_X1 U915 ( .A(KEYINPUT101), .B(n823), .Z(n824) );
  NAND2_X1 U916 ( .A1(n825), .A2(n824), .ZN(G188) );
  XOR2_X1 U917 ( .A(G120), .B(KEYINPUT102), .Z(G236) );
  INV_X1 U919 ( .A(G132), .ZN(G219) );
  INV_X1 U920 ( .A(G108), .ZN(G238) );
  INV_X1 U921 ( .A(G82), .ZN(G220) );
  NOR2_X1 U922 ( .A1(n827), .A2(n826), .ZN(G325) );
  INV_X1 U923 ( .A(G325), .ZN(G261) );
  XOR2_X1 U924 ( .A(KEYINPUT41), .B(G1981), .Z(n829) );
  XNOR2_X1 U925 ( .A(G1961), .B(G1956), .ZN(n828) );
  XNOR2_X1 U926 ( .A(n829), .B(n828), .ZN(n830) );
  XOR2_X1 U927 ( .A(n830), .B(KEYINPUT104), .Z(n832) );
  XNOR2_X1 U928 ( .A(G1996), .B(G1991), .ZN(n831) );
  XNOR2_X1 U929 ( .A(n832), .B(n831), .ZN(n836) );
  XOR2_X1 U930 ( .A(G1986), .B(G1976), .Z(n834) );
  XNOR2_X1 U931 ( .A(G1966), .B(G1971), .ZN(n833) );
  XNOR2_X1 U932 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U933 ( .A(n836), .B(n835), .Z(n838) );
  XNOR2_X1 U934 ( .A(KEYINPUT103), .B(G2474), .ZN(n837) );
  XNOR2_X1 U935 ( .A(n838), .B(n837), .ZN(G229) );
  XOR2_X1 U936 ( .A(G2100), .B(G2096), .Z(n840) );
  XNOR2_X1 U937 ( .A(KEYINPUT42), .B(G2678), .ZN(n839) );
  XNOR2_X1 U938 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U939 ( .A(KEYINPUT43), .B(G2090), .Z(n842) );
  XNOR2_X1 U940 ( .A(G2067), .B(G2072), .ZN(n841) );
  XNOR2_X1 U941 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U942 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U943 ( .A(G2078), .B(G2084), .ZN(n845) );
  XNOR2_X1 U944 ( .A(n846), .B(n845), .ZN(G227) );
  NAND2_X1 U945 ( .A1(G100), .A2(n868), .ZN(n848) );
  NAND2_X1 U946 ( .A1(G112), .A2(n872), .ZN(n847) );
  NAND2_X1 U947 ( .A1(n848), .A2(n847), .ZN(n849) );
  XNOR2_X1 U948 ( .A(KEYINPUT106), .B(n849), .ZN(n855) );
  NAND2_X1 U949 ( .A1(n871), .A2(G124), .ZN(n850) );
  XNOR2_X1 U950 ( .A(n850), .B(KEYINPUT44), .ZN(n852) );
  NAND2_X1 U951 ( .A1(G136), .A2(n533), .ZN(n851) );
  NAND2_X1 U952 ( .A1(n852), .A2(n851), .ZN(n853) );
  XOR2_X1 U953 ( .A(KEYINPUT105), .B(n853), .Z(n854) );
  NOR2_X1 U954 ( .A1(n855), .A2(n854), .ZN(G162) );
  NAND2_X1 U955 ( .A1(G106), .A2(n868), .ZN(n857) );
  NAND2_X1 U956 ( .A1(G142), .A2(n533), .ZN(n856) );
  NAND2_X1 U957 ( .A1(n857), .A2(n856), .ZN(n858) );
  XNOR2_X1 U958 ( .A(n858), .B(KEYINPUT45), .ZN(n860) );
  NAND2_X1 U959 ( .A1(G130), .A2(n871), .ZN(n859) );
  NAND2_X1 U960 ( .A1(n860), .A2(n859), .ZN(n863) );
  NAND2_X1 U961 ( .A1(G118), .A2(n872), .ZN(n861) );
  XNOR2_X1 U962 ( .A(KEYINPUT107), .B(n861), .ZN(n862) );
  NOR2_X1 U963 ( .A1(n863), .A2(n862), .ZN(n864) );
  XNOR2_X1 U964 ( .A(G160), .B(n864), .ZN(n888) );
  XNOR2_X1 U965 ( .A(G162), .B(n865), .ZN(n867) );
  XNOR2_X1 U966 ( .A(n867), .B(n866), .ZN(n881) );
  NAND2_X1 U967 ( .A1(G103), .A2(n868), .ZN(n870) );
  NAND2_X1 U968 ( .A1(G139), .A2(n533), .ZN(n869) );
  NAND2_X1 U969 ( .A1(n870), .A2(n869), .ZN(n878) );
  NAND2_X1 U970 ( .A1(G127), .A2(n871), .ZN(n874) );
  NAND2_X1 U971 ( .A1(G115), .A2(n872), .ZN(n873) );
  NAND2_X1 U972 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U973 ( .A(KEYINPUT47), .B(n875), .ZN(n876) );
  XNOR2_X1 U974 ( .A(KEYINPUT109), .B(n876), .ZN(n877) );
  NOR2_X1 U975 ( .A1(n878), .A2(n877), .ZN(n955) );
  XNOR2_X1 U976 ( .A(G164), .B(n955), .ZN(n879) );
  XNOR2_X1 U977 ( .A(n879), .B(n938), .ZN(n880) );
  XOR2_X1 U978 ( .A(n881), .B(n880), .Z(n886) );
  XOR2_X1 U979 ( .A(KEYINPUT108), .B(KEYINPUT46), .Z(n883) );
  XNOR2_X1 U980 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n882) );
  XNOR2_X1 U981 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U982 ( .A(KEYINPUT48), .B(n884), .ZN(n885) );
  XNOR2_X1 U983 ( .A(n886), .B(n885), .ZN(n887) );
  XNOR2_X1 U984 ( .A(n888), .B(n887), .ZN(n890) );
  XOR2_X1 U985 ( .A(n890), .B(n889), .Z(n891) );
  NOR2_X1 U986 ( .A1(G37), .A2(n891), .ZN(G395) );
  XNOR2_X1 U987 ( .A(G286), .B(n976), .ZN(n893) );
  XNOR2_X1 U988 ( .A(n893), .B(n892), .ZN(n894) );
  XNOR2_X1 U989 ( .A(n894), .B(G301), .ZN(n895) );
  NOR2_X1 U990 ( .A1(G37), .A2(n895), .ZN(G397) );
  XOR2_X1 U991 ( .A(G2451), .B(G2443), .Z(n897) );
  XNOR2_X1 U992 ( .A(G2427), .B(G2454), .ZN(n896) );
  XNOR2_X1 U993 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U994 ( .A(n898), .B(G2446), .Z(n900) );
  XNOR2_X1 U995 ( .A(G1341), .B(G1348), .ZN(n899) );
  XNOR2_X1 U996 ( .A(n900), .B(n899), .ZN(n904) );
  XOR2_X1 U997 ( .A(G2435), .B(KEYINPUT100), .Z(n902) );
  XNOR2_X1 U998 ( .A(G2430), .B(G2438), .ZN(n901) );
  XNOR2_X1 U999 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U1000 ( .A(n904), .B(n903), .Z(n905) );
  NAND2_X1 U1001 ( .A1(G14), .A2(n905), .ZN(n911) );
  NAND2_X1 U1002 ( .A1(G319), .A2(n911), .ZN(n908) );
  NOR2_X1 U1003 ( .A1(G229), .A2(G227), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(KEYINPUT49), .B(n906), .ZN(n907) );
  NOR2_X1 U1005 ( .A1(n908), .A2(n907), .ZN(n910) );
  NOR2_X1 U1006 ( .A1(G395), .A2(G397), .ZN(n909) );
  NAND2_X1 U1007 ( .A1(n910), .A2(n909), .ZN(G225) );
  INV_X1 U1008 ( .A(G225), .ZN(G308) );
  INV_X1 U1009 ( .A(G69), .ZN(G235) );
  INV_X1 U1010 ( .A(G96), .ZN(G221) );
  INV_X1 U1011 ( .A(n911), .ZN(G401) );
  XNOR2_X1 U1012 ( .A(KEYINPUT126), .B(KEYINPUT127), .ZN(n1022) );
  XNOR2_X1 U1013 ( .A(G5), .B(n912), .ZN(n926) );
  XOR2_X1 U1014 ( .A(G1956), .B(G20), .Z(n918) );
  XOR2_X1 U1015 ( .A(G1981), .B(G6), .Z(n913) );
  XNOR2_X1 U1016 ( .A(KEYINPUT123), .B(n913), .ZN(n915) );
  XNOR2_X1 U1017 ( .A(G19), .B(G1341), .ZN(n914) );
  NOR2_X1 U1018 ( .A1(n915), .A2(n914), .ZN(n916) );
  XNOR2_X1 U1019 ( .A(KEYINPUT124), .B(n916), .ZN(n917) );
  NAND2_X1 U1020 ( .A1(n918), .A2(n917), .ZN(n921) );
  XOR2_X1 U1021 ( .A(KEYINPUT59), .B(G1348), .Z(n919) );
  XNOR2_X1 U1022 ( .A(G4), .B(n919), .ZN(n920) );
  NOR2_X1 U1023 ( .A1(n921), .A2(n920), .ZN(n922) );
  XOR2_X1 U1024 ( .A(KEYINPUT60), .B(n922), .Z(n924) );
  XNOR2_X1 U1025 ( .A(G1966), .B(G21), .ZN(n923) );
  NOR2_X1 U1026 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1027 ( .A1(n926), .A2(n925), .ZN(n934) );
  XNOR2_X1 U1028 ( .A(G1971), .B(G22), .ZN(n928) );
  XNOR2_X1 U1029 ( .A(G23), .B(G1976), .ZN(n927) );
  NOR2_X1 U1030 ( .A1(n928), .A2(n927), .ZN(n931) );
  XNOR2_X1 U1031 ( .A(G1986), .B(KEYINPUT125), .ZN(n929) );
  XNOR2_X1 U1032 ( .A(n929), .B(G24), .ZN(n930) );
  NAND2_X1 U1033 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1034 ( .A(KEYINPUT58), .B(n932), .ZN(n933) );
  NOR2_X1 U1035 ( .A1(n934), .A2(n933), .ZN(n935) );
  XOR2_X1 U1036 ( .A(KEYINPUT61), .B(n935), .Z(n936) );
  NOR2_X1 U1037 ( .A1(G16), .A2(n936), .ZN(n1020) );
  NOR2_X1 U1038 ( .A1(n938), .A2(n937), .ZN(n942) );
  XOR2_X1 U1039 ( .A(G160), .B(G2084), .Z(n939) );
  NOR2_X1 U1040 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1041 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1042 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1043 ( .A(n945), .B(KEYINPUT112), .ZN(n947) );
  NAND2_X1 U1044 ( .A1(n947), .A2(n946), .ZN(n953) );
  XNOR2_X1 U1045 ( .A(G2090), .B(G162), .ZN(n948) );
  XNOR2_X1 U1046 ( .A(n948), .B(KEYINPUT113), .ZN(n950) );
  NOR2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1048 ( .A(KEYINPUT51), .B(n951), .ZN(n952) );
  NOR2_X1 U1049 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1050 ( .A(n954), .B(KEYINPUT114), .ZN(n961) );
  XNOR2_X1 U1051 ( .A(KEYINPUT50), .B(KEYINPUT115), .ZN(n959) );
  XNOR2_X1 U1052 ( .A(G2072), .B(n955), .ZN(n957) );
  XNOR2_X1 U1053 ( .A(G164), .B(G2078), .ZN(n956) );
  NAND2_X1 U1054 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1055 ( .A(n959), .B(n958), .ZN(n960) );
  NAND2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1057 ( .A(n962), .B(KEYINPUT52), .ZN(n963) );
  NAND2_X1 U1058 ( .A1(n963), .A2(G29), .ZN(n991) );
  XNOR2_X1 U1059 ( .A(G1966), .B(G168), .ZN(n965) );
  NAND2_X1 U1060 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1061 ( .A(n966), .B(KEYINPUT120), .ZN(n967) );
  XOR2_X1 U1062 ( .A(KEYINPUT57), .B(n967), .Z(n986) );
  NAND2_X1 U1063 ( .A1(G1971), .A2(G303), .ZN(n968) );
  NAND2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n971) );
  XNOR2_X1 U1065 ( .A(G1956), .B(G299), .ZN(n970) );
  NOR2_X1 U1066 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n974) );
  NOR2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n980) );
  XNOR2_X1 U1069 ( .A(G301), .B(G1961), .ZN(n978) );
  XNOR2_X1 U1070 ( .A(n976), .B(G1348), .ZN(n977) );
  NOR2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n983) );
  XNOR2_X1 U1073 ( .A(G1341), .B(n981), .ZN(n982) );
  NOR2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1075 ( .A(KEYINPUT121), .B(n984), .ZN(n985) );
  NOR2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n987) );
  XOR2_X1 U1077 ( .A(KEYINPUT122), .B(n987), .Z(n989) );
  XNOR2_X1 U1078 ( .A(G16), .B(KEYINPUT56), .ZN(n988) );
  NAND2_X1 U1079 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n1017) );
  XNOR2_X1 U1081 ( .A(G27), .B(n992), .ZN(n996) );
  XNOR2_X1 U1082 ( .A(KEYINPUT116), .B(G32), .ZN(n994) );
  XNOR2_X1 U1083 ( .A(n994), .B(n993), .ZN(n995) );
  NAND2_X1 U1084 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1085 ( .A(KEYINPUT117), .B(n997), .ZN(n999) );
  XOR2_X1 U1086 ( .A(G2072), .B(G33), .Z(n998) );
  NAND2_X1 U1087 ( .A1(n999), .A2(n998), .ZN(n1001) );
  XNOR2_X1 U1088 ( .A(G26), .B(G2067), .ZN(n1000) );
  NOR2_X1 U1089 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1090 ( .A(KEYINPUT118), .B(n1002), .ZN(n1003) );
  NAND2_X1 U1091 ( .A1(n1003), .A2(G28), .ZN(n1006) );
  XNOR2_X1 U1092 ( .A(G25), .B(n1004), .ZN(n1005) );
  NOR2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XOR2_X1 U1094 ( .A(KEYINPUT53), .B(n1007), .Z(n1010) );
  XOR2_X1 U1095 ( .A(KEYINPUT54), .B(G34), .Z(n1008) );
  XNOR2_X1 U1096 ( .A(G2084), .B(n1008), .ZN(n1009) );
  NAND2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  XNOR2_X1 U1098 ( .A(G35), .B(G2090), .ZN(n1011) );
  NOR2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XOR2_X1 U1100 ( .A(KEYINPUT119), .B(n1013), .Z(n1014) );
  NOR2_X1 U1101 ( .A1(G29), .A2(n1014), .ZN(n1015) );
  XOR2_X1 U1102 ( .A(KEYINPUT55), .B(n1015), .Z(n1016) );
  NOR2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1104 ( .A1(n1018), .A2(G11), .ZN(n1019) );
  NOR2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1106 ( .A(n1022), .B(n1021), .ZN(n1023) );
  XNOR2_X1 U1107 ( .A(KEYINPUT62), .B(n1023), .ZN(G150) );
  INV_X1 U1108 ( .A(G150), .ZN(G311) );
endmodule

