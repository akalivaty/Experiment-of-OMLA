//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 0 0 0 1 1 1 0 1 0 1 0 1 0 0 0 0 1 0 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 0 0 0 0 0 1 1 1 1 0 0 0 1 1 1 0 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:45 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n772, new_n773, new_n774, new_n775, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034;
  XNOR2_X1  g000(.A(G125), .B(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT16), .ZN(new_n188));
  INV_X1    g002(.A(G140), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G125), .ZN(new_n190));
  OAI211_X1 g004(.A(new_n188), .B(G146), .C1(KEYINPUT16), .C2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G119), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G128), .ZN(new_n193));
  INV_X1    g007(.A(G128), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G119), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT24), .B(G110), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n194), .A2(KEYINPUT23), .A3(G119), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n192), .A2(G128), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n193), .B(new_n199), .C1(new_n200), .C2(KEYINPUT23), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n198), .B1(new_n201), .B2(G110), .ZN(new_n202));
  INV_X1    g016(.A(G146), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n187), .A2(new_n203), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n191), .A2(new_n202), .A3(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT76), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n191), .A2(new_n202), .A3(KEYINPUT76), .A4(new_n204), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n188), .B1(KEYINPUT16), .B2(new_n190), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(new_n203), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(new_n191), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n196), .A2(new_n197), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n213), .B1(G110), .B2(new_n201), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g029(.A(KEYINPUT22), .B(G137), .ZN(new_n216));
  INV_X1    g030(.A(G953), .ZN(new_n217));
  AND3_X1   g031(.A1(new_n217), .A2(G221), .A3(G234), .ZN(new_n218));
  XOR2_X1   g032(.A(new_n216), .B(new_n218), .Z(new_n219));
  NAND3_X1  g033(.A1(new_n209), .A2(new_n215), .A3(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n219), .B1(new_n209), .B2(new_n215), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G902), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n223), .A2(KEYINPUT25), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n209), .A2(new_n215), .ZN(new_n226));
  INV_X1    g040(.A(new_n219), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(new_n224), .A3(new_n220), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT25), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n225), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G217), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n233), .B1(G234), .B2(new_n224), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT77), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n234), .A2(G902), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n223), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n235), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n234), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n240), .B1(new_n225), .B2(new_n231), .ZN(new_n241));
  INV_X1    g055(.A(new_n238), .ZN(new_n242));
  OAI21_X1  g056(.A(KEYINPUT77), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n239), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  NOR2_X1   g059(.A1(G237), .A2(G953), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G210), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n247), .B(KEYINPUT27), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT26), .B(G101), .ZN(new_n249));
  XNOR2_X1  g063(.A(new_n248), .B(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT70), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n203), .A2(G143), .ZN(new_n252));
  INV_X1    g066(.A(G143), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G146), .ZN(new_n254));
  AND2_X1   g068(.A1(KEYINPUT0), .A2(G128), .ZN(new_n255));
  AND3_X1   g069(.A1(new_n252), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  NOR2_X1   g070(.A1(KEYINPUT0), .A2(G128), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT64), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n257), .B(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n255), .B1(new_n252), .B2(new_n254), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n256), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G137), .ZN(new_n262));
  AOI21_X1  g076(.A(KEYINPUT65), .B1(new_n262), .B2(G134), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT11), .ZN(new_n264));
  OAI22_X1  g078(.A1(new_n263), .A2(new_n264), .B1(G134), .B2(new_n262), .ZN(new_n265));
  AOI211_X1 g079(.A(KEYINPUT65), .B(KEYINPUT11), .C1(new_n262), .C2(G134), .ZN(new_n266));
  NOR3_X1   g080(.A1(new_n265), .A2(G131), .A3(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(G131), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n262), .A2(G134), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT65), .ZN(new_n270));
  INV_X1    g084(.A(G134), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n270), .B1(new_n271), .B2(G137), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n269), .B1(new_n272), .B2(KEYINPUT11), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n263), .A2(new_n264), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n268), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n251), .B(new_n261), .C1(new_n267), .C2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(G131), .B1(new_n265), .B2(new_n266), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n273), .A2(new_n268), .A3(new_n274), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n251), .B1(new_n280), .B2(new_n261), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n277), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT72), .ZN(new_n283));
  INV_X1    g097(.A(G116), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(KEYINPUT68), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT68), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(G116), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n285), .A2(new_n287), .A3(G119), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n284), .A2(G119), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT69), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT67), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT2), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n294), .A2(G113), .ZN(new_n295));
  INV_X1    g109(.A(G113), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n296), .A2(KEYINPUT2), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n293), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n296), .A2(KEYINPUT2), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n294), .A2(G113), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n299), .A2(new_n300), .A3(KEYINPUT67), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n291), .A2(new_n292), .A3(new_n298), .A4(new_n301), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n288), .B(new_n290), .C1(new_n295), .C2(new_n297), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AND3_X1   g118(.A1(new_n299), .A2(new_n300), .A3(KEYINPUT67), .ZN(new_n305));
  AOI21_X1  g119(.A(KEYINPUT67), .B1(new_n299), .B2(new_n300), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n292), .B1(new_n307), .B2(new_n291), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n283), .B1(new_n304), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n298), .A2(new_n301), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT68), .B(G116), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n289), .B1(new_n311), .B2(G119), .ZN(new_n312));
  OAI21_X1  g126(.A(KEYINPUT69), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n313), .A2(KEYINPUT72), .A3(new_n303), .A4(new_n302), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n252), .A2(new_n254), .ZN(new_n315));
  OAI211_X1 g129(.A(KEYINPUT66), .B(KEYINPUT1), .C1(new_n253), .C2(G146), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G128), .ZN(new_n317));
  AOI21_X1  g131(.A(KEYINPUT66), .B1(new_n252), .B2(KEYINPUT1), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n315), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT1), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n252), .A2(new_n254), .A3(new_n320), .A4(G128), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(KEYINPUT71), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n271), .A2(G137), .ZN(new_n324));
  OAI21_X1  g138(.A(G131), .B1(new_n269), .B2(new_n324), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n279), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT71), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n319), .A2(new_n327), .A3(new_n321), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n323), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n282), .A2(new_n309), .A3(new_n314), .A4(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n322), .A2(new_n325), .A3(new_n279), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT30), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n261), .B1(new_n267), .B2(new_n275), .ZN(new_n333));
  AND3_X1   g147(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(KEYINPUT70), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n329), .A2(new_n335), .A3(new_n276), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n334), .B1(new_n336), .B2(KEYINPUT30), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n304), .A2(new_n308), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n250), .B(new_n330), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(KEYINPUT31), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT73), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n339), .A2(KEYINPUT73), .A3(KEYINPUT31), .ZN(new_n343));
  OR2_X1    g157(.A1(new_n337), .A2(new_n338), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT31), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n344), .A2(new_n345), .A3(new_n250), .A4(new_n330), .ZN(new_n346));
  INV_X1    g160(.A(new_n250), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT28), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n331), .A2(new_n333), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n313), .A2(new_n303), .A3(new_n302), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n348), .B1(new_n330), .B2(new_n351), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n329), .A2(new_n333), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n309), .A2(new_n314), .ZN(new_n354));
  AOI21_X1  g168(.A(KEYINPUT28), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n347), .B1(new_n352), .B2(new_n355), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n342), .A2(new_n343), .A3(new_n346), .A4(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G472), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n358), .A3(new_n224), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(KEYINPUT32), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT32), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n357), .A2(new_n361), .A3(new_n358), .A4(new_n224), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n309), .A2(new_n314), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n351), .B1(new_n336), .B2(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n355), .B1(KEYINPUT28), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(new_n250), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT29), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n337), .A2(new_n338), .ZN(new_n369));
  INV_X1    g183(.A(new_n330), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n347), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n367), .A2(new_n368), .A3(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT74), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n367), .A2(KEYINPUT74), .A3(new_n368), .A4(new_n371), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT75), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n355), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n336), .A2(new_n364), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n348), .B1(new_n330), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n329), .A2(new_n333), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n348), .B1(new_n380), .B2(new_n364), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT75), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n377), .B1(new_n379), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n347), .A2(new_n368), .ZN(new_n384));
  AOI21_X1  g198(.A(G902), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n374), .A2(new_n375), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G472), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n245), .B1(new_n363), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G221), .ZN(new_n389));
  XNOR2_X1  g203(.A(KEYINPUT9), .B(G234), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n390), .B(KEYINPUT78), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n389), .B1(new_n391), .B2(new_n224), .ZN(new_n392));
  INV_X1    g206(.A(G478), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n393), .A2(KEYINPUT15), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n391), .A2(G217), .A3(new_n217), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n194), .A2(G143), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT95), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n398), .B1(new_n194), .B2(G143), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n253), .A2(KEYINPUT95), .A3(G128), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT13), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n397), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n401), .A2(new_n402), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT96), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n401), .A2(KEYINPUT96), .A3(new_n402), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n403), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n408), .A2(new_n271), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n401), .A2(new_n271), .A3(new_n397), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n311), .A2(G122), .ZN(new_n411));
  INV_X1    g225(.A(G107), .ZN(new_n412));
  OAI21_X1  g226(.A(KEYINPUT94), .B1(new_n284), .B2(G122), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT94), .ZN(new_n414));
  INV_X1    g228(.A(G122), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n414), .A2(new_n415), .A3(G116), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n411), .A2(new_n412), .A3(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n412), .B1(new_n411), .B2(new_n417), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n410), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n409), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n401), .A2(new_n397), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(G134), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n410), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n418), .ZN(new_n426));
  OAI21_X1  g240(.A(KEYINPUT97), .B1(new_n411), .B2(KEYINPUT14), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT97), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT14), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n311), .A2(new_n428), .A3(new_n429), .A4(G122), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n411), .A2(KEYINPUT14), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n427), .A2(new_n417), .A3(new_n430), .A4(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n426), .B1(new_n432), .B2(G107), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n396), .B1(new_n422), .B2(new_n433), .ZN(new_n434));
  OAI221_X1 g248(.A(new_n410), .B1(new_n419), .B2(new_n420), .C1(new_n408), .C2(new_n271), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n432), .A2(G107), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n419), .B1(new_n410), .B2(new_n424), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n396), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n435), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(G902), .B1(new_n434), .B2(new_n440), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n441), .A2(KEYINPUT98), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT98), .ZN(new_n443));
  AOI211_X1 g257(.A(new_n443), .B(G902), .C1(new_n434), .C2(new_n440), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n395), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(G475), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n246), .A2(G214), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n253), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n246), .A2(G143), .A3(G214), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G131), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT17), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n448), .A2(new_n268), .A3(new_n449), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n450), .A2(KEYINPUT17), .A3(G131), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n454), .A2(new_n211), .A3(new_n191), .A4(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n450), .ZN(new_n457));
  NAND2_X1  g271(.A1(KEYINPUT18), .A2(G131), .ZN(new_n458));
  OR2_X1    g272(.A1(new_n187), .A2(new_n203), .ZN(new_n459));
  AOI22_X1  g273(.A1(new_n457), .A2(new_n458), .B1(new_n204), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n458), .ZN(new_n461));
  AND3_X1   g275(.A1(new_n450), .A2(KEYINPUT90), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(KEYINPUT90), .B1(new_n450), .B2(new_n461), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(G113), .B(G122), .ZN(new_n465));
  INV_X1    g279(.A(G104), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n465), .B(new_n466), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n467), .B(KEYINPUT92), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n456), .A2(new_n464), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n467), .B1(new_n456), .B2(new_n464), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n224), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n446), .B1(new_n471), .B2(KEYINPUT93), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT93), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n473), .B(new_n224), .C1(new_n469), .C2(new_n470), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n451), .A2(new_n453), .ZN(new_n475));
  AND2_X1   g289(.A1(KEYINPUT91), .A2(KEYINPUT19), .ZN(new_n476));
  NOR2_X1   g290(.A1(KEYINPUT91), .A2(KEYINPUT19), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n187), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n478), .B1(new_n187), .B2(new_n477), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n475), .B(new_n191), .C1(G146), .C2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n467), .B1(new_n464), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n469), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(G475), .A2(G902), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(KEYINPUT20), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT20), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n486), .B(new_n483), .C1(new_n469), .C2(new_n481), .ZN(new_n487));
  AOI22_X1  g301(.A1(new_n472), .A2(new_n474), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n435), .A2(new_n438), .A3(new_n439), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n439), .B1(new_n435), .B2(new_n438), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n224), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n394), .B1(new_n491), .B2(new_n443), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n445), .A2(new_n488), .A3(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(G952), .ZN(new_n494));
  AOI211_X1 g308(.A(G953), .B(new_n494), .C1(G234), .C2(G237), .ZN(new_n495));
  AOI211_X1 g309(.A(new_n224), .B(new_n217), .C1(G234), .C2(G237), .ZN(new_n496));
  XNOR2_X1  g310(.A(KEYINPUT21), .B(G898), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n493), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(KEYINPUT3), .B1(new_n466), .B2(G107), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT3), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n502), .A2(new_n412), .A3(G104), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n466), .A2(G107), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n501), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(G101), .ZN(new_n506));
  INV_X1    g320(.A(G101), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n501), .A2(new_n503), .A3(new_n507), .A4(new_n504), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n506), .A2(KEYINPUT4), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT4), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n505), .A2(new_n510), .A3(G101), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n509), .A2(new_n261), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT79), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT79), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n509), .A2(new_n514), .A3(new_n261), .A4(new_n511), .ZN(new_n515));
  AND2_X1   g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n466), .A2(G107), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n412), .A2(G104), .ZN(new_n518));
  OAI21_X1  g332(.A(G101), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n508), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n323), .A2(KEYINPUT10), .A3(new_n328), .A4(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n252), .A2(KEYINPUT1), .ZN(new_n523));
  AOI22_X1  g337(.A1(new_n523), .A2(G128), .B1(new_n252), .B2(new_n254), .ZN(new_n524));
  INV_X1    g338(.A(new_n321), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n508), .B(new_n519), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT10), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n522), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n280), .B1(new_n516), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT80), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g346(.A(KEYINPUT80), .B(new_n280), .C1(new_n516), .C2(new_n529), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n513), .A2(new_n515), .ZN(new_n535));
  INV_X1    g349(.A(new_n280), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n535), .A2(new_n536), .A3(new_n522), .A4(new_n528), .ZN(new_n537));
  XNOR2_X1  g351(.A(G110), .B(G140), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n217), .A2(G227), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n538), .B(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n534), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT81), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n526), .B1(new_n322), .B2(new_n521), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n280), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT12), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n546), .A2(KEYINPUT12), .A3(new_n280), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n541), .B1(new_n537), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n544), .A2(new_n545), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n542), .B1(new_n532), .B2(new_n533), .ZN(new_n555));
  OAI21_X1  g369(.A(KEYINPUT81), .B1(new_n555), .B2(new_n552), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n554), .A2(new_n556), .A3(G469), .ZN(new_n557));
  INV_X1    g371(.A(G469), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n558), .A2(new_n224), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  AND2_X1   g374(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n534), .A2(new_n537), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n540), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n542), .A2(KEYINPUT83), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT83), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n537), .A2(new_n565), .A3(new_n541), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  AND3_X1   g381(.A1(new_n546), .A2(KEYINPUT12), .A3(new_n280), .ZN(new_n568));
  AOI21_X1  g382(.A(KEYINPUT12), .B1(new_n546), .B2(new_n280), .ZN(new_n569));
  OAI21_X1  g383(.A(KEYINPUT82), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT82), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n549), .A2(new_n571), .A3(new_n550), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(KEYINPUT84), .B1(new_n567), .B2(new_n573), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n537), .A2(new_n565), .A3(new_n541), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n565), .B1(new_n537), .B2(new_n541), .ZN(new_n576));
  OAI211_X1 g390(.A(KEYINPUT84), .B(new_n573), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n563), .B1(new_n574), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n579), .A2(new_n558), .A3(new_n224), .ZN(new_n580));
  AOI211_X1 g394(.A(new_n392), .B(new_n500), .C1(new_n561), .C2(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(G214), .B1(G237), .B2(G902), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n509), .A2(new_n511), .ZN(new_n583));
  OAI21_X1  g397(.A(KEYINPUT85), .B1(new_n338), .B2(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(G110), .B(G122), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT5), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n296), .B1(new_n289), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n587), .B1(new_n291), .B2(new_n586), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n588), .A2(new_n521), .A3(new_n303), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT85), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n350), .A2(new_n590), .A3(new_n511), .A4(new_n509), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n584), .A2(new_n585), .A3(new_n589), .A4(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(KEYINPUT86), .ZN(new_n593));
  INV_X1    g407(.A(new_n589), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n302), .A2(new_n303), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n583), .B1(new_n595), .B2(new_n313), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n594), .B1(new_n596), .B2(new_n590), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT86), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n597), .A2(new_n598), .A3(new_n585), .A4(new_n584), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n593), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(G125), .ZN(new_n601));
  OR2_X1    g415(.A1(new_n261), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n319), .A2(new_n601), .A3(new_n321), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(G224), .ZN(new_n605));
  OAI21_X1  g419(.A(KEYINPUT7), .B1(new_n605), .B2(G953), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n602), .A2(new_n603), .A3(new_n606), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n585), .B(KEYINPUT8), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n521), .B1(new_n588), .B2(new_n303), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n611), .B1(new_n594), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n600), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT88), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n616), .A2(new_n617), .A3(new_n224), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n614), .B1(new_n593), .B2(new_n599), .ZN(new_n619));
  OAI21_X1  g433(.A(KEYINPUT88), .B1(new_n619), .B2(G902), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n585), .B1(new_n597), .B2(new_n584), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(KEYINPUT6), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT6), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n623), .B1(new_n593), .B2(new_n599), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n622), .B1(new_n624), .B2(new_n621), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n605), .A2(G953), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(KEYINPUT87), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n604), .B(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  AOI22_X1  g443(.A1(new_n618), .A2(new_n620), .B1(new_n625), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g444(.A(G210), .B1(G237), .B2(G902), .ZN(new_n631));
  OAI21_X1  g445(.A(KEYINPUT89), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT89), .ZN(new_n633));
  INV_X1    g447(.A(new_n631), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n617), .B1(new_n616), .B2(new_n224), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n619), .A2(KEYINPUT88), .A3(G902), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n600), .A2(KEYINPUT6), .ZN(new_n638));
  INV_X1    g452(.A(new_n621), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n628), .B1(new_n640), .B2(new_n622), .ZN(new_n641));
  OAI211_X1 g455(.A(new_n633), .B(new_n634), .C1(new_n637), .C2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n630), .A2(new_n631), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n632), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n388), .A2(new_n581), .A3(new_n582), .A4(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G101), .ZN(G3));
  INV_X1    g460(.A(KEYINPUT100), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n441), .A2(new_n647), .A3(G478), .ZN(new_n648));
  AOI21_X1  g462(.A(KEYINPUT100), .B1(new_n491), .B2(new_n393), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n393), .A2(G902), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT99), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n653), .B1(new_n489), .B2(new_n490), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT33), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n653), .B(KEYINPUT33), .C1(new_n489), .C2(new_n490), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n652), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  OR2_X1    g472(.A1(new_n650), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n472), .A2(new_n474), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n485), .A2(new_n487), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n499), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n618), .A2(new_n620), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n625), .A2(new_n629), .ZN(new_n667));
  AND3_X1   g481(.A1(new_n666), .A2(new_n631), .A3(new_n667), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n631), .B1(new_n666), .B2(new_n667), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n582), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n665), .A2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n392), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n541), .B1(new_n534), .B2(new_n537), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n573), .B1(new_n575), .B2(new_n576), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT84), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n673), .B1(new_n676), .B2(new_n577), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n677), .A2(G469), .A3(G902), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n557), .A2(new_n560), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n672), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  OAI22_X1  g494(.A1(new_n366), .A2(new_n250), .B1(new_n339), .B2(KEYINPUT31), .ZN(new_n681));
  AND3_X1   g495(.A1(new_n339), .A2(KEYINPUT73), .A3(KEYINPUT31), .ZN(new_n682));
  AOI21_X1  g496(.A(KEYINPUT73), .B1(new_n339), .B2(KEYINPUT31), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n681), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g498(.A(G472), .B1(new_n684), .B2(G902), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n685), .A2(new_n244), .A3(new_n359), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n680), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n671), .A2(new_n687), .ZN(new_n688));
  XOR2_X1   g502(.A(KEYINPUT34), .B(G104), .Z(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G6));
  AND2_X1   g504(.A1(new_n445), .A2(new_n492), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n691), .A2(new_n662), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n499), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n670), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n687), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G107), .ZN(new_n696));
  XNOR2_X1  g510(.A(KEYINPUT101), .B(KEYINPUT35), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G9));
  NAND2_X1  g512(.A1(new_n685), .A2(new_n359), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n227), .A2(KEYINPUT36), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n226), .B(new_n700), .ZN(new_n701));
  AND2_X1   g515(.A1(new_n701), .A2(new_n237), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n241), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(KEYINPUT102), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT102), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n705), .B1(new_n241), .B2(new_n702), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n699), .A2(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n581), .A2(new_n582), .A3(new_n644), .A4(new_n708), .ZN(new_n709));
  XOR2_X1   g523(.A(KEYINPUT37), .B(G110), .Z(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G12));
  AOI21_X1  g525(.A(new_n707), .B1(new_n363), .B2(new_n387), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n680), .A2(new_n670), .ZN(new_n713));
  AND2_X1   g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n495), .ZN(new_n715));
  INV_X1    g529(.A(new_n496), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n715), .B1(new_n716), .B2(G900), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n692), .A2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n714), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G128), .ZN(G30));
  XNOR2_X1  g535(.A(new_n717), .B(KEYINPUT39), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n680), .A2(new_n723), .ZN(new_n724));
  XOR2_X1   g538(.A(new_n724), .B(KEYINPUT40), .Z(new_n725));
  XOR2_X1   g539(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n726));
  XNOR2_X1  g540(.A(new_n644), .B(new_n726), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n330), .A2(new_n378), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n339), .B1(new_n728), .B2(new_n250), .ZN(new_n729));
  AND2_X1   g543(.A1(new_n729), .A2(new_n224), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n363), .B1(new_n358), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n691), .A2(new_n488), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n731), .A2(new_n582), .A3(new_n703), .A4(new_n732), .ZN(new_n733));
  OR3_X1    g547(.A1(new_n725), .A2(new_n727), .A3(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G143), .ZN(G45));
  OAI211_X1 g549(.A(new_n662), .B(new_n717), .C1(new_n650), .C2(new_n658), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n714), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G146), .ZN(G48));
  OAI21_X1  g553(.A(G469), .B1(new_n677), .B2(G902), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(new_n580), .A3(new_n672), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT104), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n740), .A2(new_n580), .A3(KEYINPUT104), .A4(new_n672), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n671), .A2(new_n388), .A3(new_n743), .A4(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(KEYINPUT41), .B(G113), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n745), .B(new_n746), .ZN(G15));
  NAND4_X1  g561(.A1(new_n388), .A2(new_n694), .A3(new_n743), .A4(new_n744), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G116), .ZN(G18));
  NAND3_X1  g563(.A1(new_n712), .A2(new_n499), .A3(new_n493), .ZN(new_n750));
  INV_X1    g564(.A(new_n582), .ZN(new_n751));
  INV_X1    g565(.A(new_n669), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n751), .B1(new_n752), .B2(new_n643), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n743), .A2(new_n753), .A3(new_n744), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n750), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(new_n192), .ZN(G21));
  OAI211_X1 g570(.A(new_n582), .B(new_n732), .C1(new_n668), .C2(new_n669), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n757), .A2(new_n498), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n358), .B1(new_n357), .B2(new_n224), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n358), .A2(new_n224), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT105), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n383), .A2(new_n761), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n377), .B(KEYINPUT105), .C1(new_n379), .C2(new_n382), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(new_n347), .A3(new_n763), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n346), .A2(new_n340), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n760), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n241), .A2(new_n242), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n759), .A2(new_n766), .A3(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n758), .A2(new_n743), .A3(new_n744), .A4(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G122), .ZN(G24));
  NOR4_X1   g585(.A1(new_n759), .A2(new_n766), .A3(new_n703), .A4(new_n736), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n743), .A2(new_n772), .A3(new_n753), .A4(new_n744), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT106), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n773), .B(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G125), .ZN(G27));
  INV_X1    g590(.A(KEYINPUT42), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n544), .A2(new_n553), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n558), .B1(new_n778), .B2(new_n224), .ZN(new_n779));
  OAI21_X1  g593(.A(KEYINPUT107), .B1(new_n678), .B2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT107), .ZN(new_n781));
  INV_X1    g595(.A(new_n779), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n580), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n780), .A2(new_n672), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n751), .B1(new_n630), .B2(new_n631), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n632), .A2(new_n785), .A3(new_n642), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT108), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n632), .A2(new_n785), .A3(new_n642), .A4(KEYINPUT108), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n784), .A2(new_n388), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n777), .B1(new_n790), .B2(new_n736), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT109), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n580), .A2(new_n782), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n392), .B1(new_n793), .B2(KEYINPUT107), .ZN(new_n794));
  AND4_X1   g608(.A1(new_n788), .A2(new_n789), .A3(new_n783), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n363), .A2(new_n387), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n736), .A2(new_n777), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(new_n767), .A3(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n792), .B1(new_n795), .B2(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n788), .A2(new_n789), .A3(new_n783), .A4(new_n794), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n801), .A2(KEYINPUT109), .A3(new_n798), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n791), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G131), .ZN(G33));
  NOR2_X1   g618(.A1(new_n790), .A2(new_n718), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(new_n271), .ZN(G36));
  NAND2_X1  g620(.A1(new_n659), .A2(new_n488), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT43), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n807), .B(new_n808), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n809), .B(new_n699), .C1(new_n241), .C2(new_n702), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(KEYINPUT44), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n788), .A2(new_n789), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(KEYINPUT45), .B1(new_n554), .B2(new_n556), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT45), .ZN(new_n816));
  OAI21_X1  g630(.A(G469), .B1(new_n778), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n560), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT46), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n818), .A2(KEYINPUT110), .A3(new_n819), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n820), .B(new_n580), .C1(new_n819), .C2(new_n818), .ZN(new_n821));
  AOI21_X1  g635(.A(KEYINPUT110), .B1(new_n818), .B2(new_n819), .ZN(new_n822));
  OR2_X1    g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(new_n672), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n824), .A2(new_n723), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n814), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(KEYINPUT111), .B(G137), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n826), .B(new_n827), .ZN(G39));
  OR4_X1    g642(.A1(new_n796), .A2(new_n812), .A3(new_n244), .A4(new_n736), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT47), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n824), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n823), .A2(KEYINPUT47), .A3(new_n672), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n829), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(new_n189), .ZN(G42));
  OR4_X1    g648(.A1(new_n768), .A2(new_n807), .A3(new_n751), .A4(new_n392), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n740), .A2(new_n580), .ZN(new_n836));
  AOI211_X1 g650(.A(new_n731), .B(new_n835), .C1(KEYINPUT49), .C2(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n836), .A2(KEYINPUT49), .ZN(new_n838));
  XOR2_X1   g652(.A(new_n838), .B(KEYINPUT112), .Z(new_n839));
  NAND3_X1  g653(.A1(new_n837), .A2(new_n727), .A3(new_n839), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n743), .A2(new_n744), .ZN(new_n841));
  AND4_X1   g655(.A1(new_n495), .A2(new_n813), .A3(new_n841), .A4(new_n809), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(KEYINPUT117), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n759), .A2(new_n766), .A3(new_n703), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n813), .A2(new_n841), .ZN(new_n845));
  NOR4_X1   g659(.A1(new_n845), .A2(new_n245), .A3(new_n715), .A4(new_n731), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n659), .A2(new_n662), .ZN(new_n847));
  AOI22_X1  g661(.A1(new_n843), .A2(new_n844), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n809), .A2(new_n495), .A3(new_n769), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n849), .A2(new_n727), .A3(new_n751), .A4(new_n841), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT50), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n850), .A2(new_n851), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  OR2_X1    g668(.A1(new_n854), .A2(KEYINPUT116), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(KEYINPUT116), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n848), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(KEYINPUT118), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT118), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n848), .A2(new_n859), .A3(new_n855), .A4(new_n856), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n813), .A2(new_n849), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n831), .A2(new_n832), .A3(KEYINPUT115), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n740), .A2(new_n580), .A3(new_n392), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT115), .B1(new_n831), .B2(new_n832), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n861), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n858), .A2(new_n860), .A3(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT51), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT53), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n663), .A2(new_n498), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n687), .A2(new_n582), .A3(new_n644), .A4(new_n871), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n645), .A2(new_n872), .A3(KEYINPUT113), .ZN(new_n873));
  AOI21_X1  g687(.A(KEYINPUT113), .B1(new_n645), .B2(new_n872), .ZN(new_n874));
  INV_X1    g688(.A(new_n693), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n687), .A2(new_n582), .A3(new_n644), .A4(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n770), .A2(new_n876), .A3(new_n709), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n873), .A2(new_n874), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n745), .A2(new_n748), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n879), .A2(new_n755), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n493), .A2(new_n717), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n680), .A2(new_n707), .A3(new_n881), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n882), .A2(new_n788), .A3(new_n796), .A4(new_n789), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n784), .A2(new_n772), .A3(new_n788), .A4(new_n789), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n883), .B(new_n884), .C1(new_n790), .C2(new_n718), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n878), .A2(new_n803), .A3(new_n880), .A4(new_n886), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n773), .B(KEYINPUT106), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n712), .B(new_n713), .C1(new_n719), .C2(new_n737), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n703), .A2(new_n717), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n757), .A2(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n891), .A2(new_n731), .A3(new_n783), .A4(new_n794), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT52), .B1(new_n888), .B2(new_n893), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n889), .A2(new_n892), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT52), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n775), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n870), .B1(new_n887), .B2(new_n898), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n888), .A2(KEYINPUT52), .A3(new_n893), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n896), .B1(new_n775), .B2(new_n895), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n645), .A2(new_n872), .A3(KEYINPUT113), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n645), .A2(new_n872), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT113), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(new_n877), .ZN(new_n907));
  AND4_X1   g721(.A1(new_n880), .A2(new_n903), .A3(new_n906), .A4(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n795), .A2(new_n792), .A3(new_n799), .ZN(new_n909));
  OAI21_X1  g723(.A(KEYINPUT109), .B1(new_n801), .B2(new_n798), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n885), .B1(new_n911), .B2(new_n791), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n902), .A2(KEYINPUT53), .A3(new_n908), .A4(new_n912), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n899), .A2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT54), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT114), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n899), .A2(new_n917), .A3(new_n913), .ZN(new_n918));
  OAI211_X1 g732(.A(KEYINPUT114), .B(new_n870), .C1(new_n887), .C2(new_n898), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT54), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n916), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n849), .A2(new_n753), .A3(new_n841), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n922), .A2(G952), .A3(new_n217), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n923), .B1(new_n846), .B2(new_n664), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n768), .B1(new_n363), .B2(new_n387), .ZN(new_n925));
  NAND2_X1  g739(.A1(KEYINPUT120), .A2(KEYINPUT48), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n843), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  OR2_X1    g741(.A1(KEYINPUT120), .A2(KEYINPUT48), .ZN(new_n928));
  AOI22_X1  g742(.A1(new_n843), .A2(new_n925), .B1(new_n928), .B2(new_n926), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n924), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n831), .A2(new_n832), .A3(new_n863), .ZN(new_n931));
  OR2_X1    g745(.A1(new_n931), .A2(KEYINPUT119), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(KEYINPUT119), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n932), .A2(new_n861), .A3(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n854), .A2(new_n868), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n848), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n930), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n869), .A2(new_n921), .A3(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(G952), .A2(G953), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n840), .B1(new_n938), .B2(new_n939), .ZN(G75));
  NAND2_X1  g754(.A1(new_n918), .A2(new_n919), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n941), .A2(new_n224), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(G210), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT56), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n625), .B(new_n628), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT55), .ZN(new_n946));
  AND3_X1   g760(.A1(new_n943), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n946), .B1(new_n943), .B2(new_n944), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n217), .A2(G952), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(G51));
  AND3_X1   g764(.A1(new_n918), .A2(KEYINPUT54), .A3(new_n919), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n951), .A2(new_n920), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n559), .B(KEYINPUT57), .Z(new_n953));
  OAI21_X1  g767(.A(new_n579), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n815), .A2(new_n817), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n942), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n949), .B1(new_n954), .B2(new_n956), .ZN(G54));
  NAND3_X1  g771(.A1(new_n942), .A2(KEYINPUT58), .A3(G475), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n958), .A2(new_n482), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n958), .A2(new_n482), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n959), .A2(new_n960), .A3(new_n949), .ZN(G60));
  INV_X1    g775(.A(KEYINPUT121), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n656), .A2(new_n657), .ZN(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(G478), .A2(G902), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT59), .Z(new_n966));
  NOR2_X1   g780(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n941), .A2(new_n915), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n918), .A2(KEYINPUT54), .A3(new_n919), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n968), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n962), .B1(new_n971), .B2(new_n949), .ZN(new_n972));
  INV_X1    g786(.A(new_n949), .ZN(new_n973));
  OAI211_X1 g787(.A(KEYINPUT121), .B(new_n973), .C1(new_n952), .C2(new_n968), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n964), .B1(new_n921), .B2(new_n966), .ZN(new_n975));
  AND3_X1   g789(.A1(new_n972), .A2(new_n974), .A3(new_n975), .ZN(G63));
  NAND2_X1  g790(.A1(G217), .A2(G902), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT60), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n918), .A2(new_n701), .A3(new_n919), .A4(new_n979), .ZN(new_n980));
  NOR2_X1   g794(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n949), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n941), .A2(new_n978), .ZN(new_n983));
  OAI211_X1 g797(.A(new_n980), .B(new_n982), .C1(new_n983), .C2(new_n223), .ZN(new_n984));
  NAND2_X1  g798(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n984), .B(new_n985), .ZN(G66));
  INV_X1    g800(.A(new_n497), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n217), .B1(new_n987), .B2(G224), .ZN(new_n988));
  INV_X1    g802(.A(new_n908), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n988), .B1(new_n989), .B2(new_n217), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n640), .B(new_n622), .C1(G898), .C2(new_n217), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT123), .Z(new_n992));
  XNOR2_X1  g806(.A(new_n990), .B(new_n992), .ZN(G69));
  AOI21_X1  g807(.A(new_n217), .B1(G227), .B2(G900), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n994), .A2(KEYINPUT126), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n775), .A2(new_n889), .ZN(new_n996));
  INV_X1    g810(.A(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n734), .A2(new_n997), .ZN(new_n998));
  OR2_X1    g812(.A1(new_n998), .A2(KEYINPUT62), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n833), .B1(new_n825), .B2(new_n814), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n998), .A2(KEYINPUT62), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n663), .B1(new_n691), .B2(new_n662), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n813), .A2(new_n388), .A3(new_n724), .A4(new_n1002), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n1003), .B(KEYINPUT124), .Z(new_n1004));
  NAND4_X1  g818(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .A4(new_n1004), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n337), .B(new_n479), .Z(new_n1006));
  AND2_X1   g820(.A1(new_n1006), .A2(new_n217), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n995), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1008), .ZN(new_n1009));
  INV_X1    g823(.A(KEYINPUT125), .ZN(new_n1010));
  AOI211_X1 g824(.A(new_n768), .B(new_n757), .C1(new_n387), .C2(new_n363), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n805), .B1(new_n825), .B2(new_n1011), .ZN(new_n1012));
  AND2_X1   g826(.A1(new_n1012), .A2(new_n803), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1000), .A2(new_n1013), .A3(new_n997), .ZN(new_n1014));
  AND2_X1   g828(.A1(new_n1014), .A2(new_n217), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n217), .A2(G900), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1010), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1016), .B1(new_n1014), .B2(new_n217), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1006), .B1(new_n1018), .B2(KEYINPUT125), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1009), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n994), .A2(KEYINPUT126), .ZN(new_n1021));
  INV_X1    g835(.A(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g836(.A(new_n1020), .B(new_n1022), .ZN(G72));
  NOR2_X1   g837(.A1(new_n369), .A2(new_n370), .ZN(new_n1024));
  XNOR2_X1  g838(.A(new_n1024), .B(KEYINPUT127), .ZN(new_n1025));
  OR2_X1    g839(.A1(new_n1005), .A2(new_n989), .ZN(new_n1026));
  NAND2_X1  g840(.A1(G472), .A2(G902), .ZN(new_n1027));
  XOR2_X1   g841(.A(new_n1027), .B(KEYINPUT63), .Z(new_n1028));
  AOI211_X1 g842(.A(new_n347), .B(new_n1025), .C1(new_n1026), .C2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n371), .A2(new_n339), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1030), .A2(new_n1028), .ZN(new_n1031));
  NOR2_X1   g845(.A1(new_n914), .A2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g846(.A(new_n1028), .B1(new_n1014), .B2(new_n989), .ZN(new_n1033));
  AND3_X1   g847(.A1(new_n1033), .A2(new_n347), .A3(new_n1025), .ZN(new_n1034));
  NOR4_X1   g848(.A1(new_n1029), .A2(new_n949), .A3(new_n1032), .A4(new_n1034), .ZN(G57));
endmodule


