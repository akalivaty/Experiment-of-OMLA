

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593;

  XNOR2_X1 U324 ( .A(n454), .B(KEYINPUT103), .ZN(n455) );
  XNOR2_X1 U325 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U326 ( .A(n457), .B(KEYINPUT38), .ZN(n504) );
  XNOR2_X1 U327 ( .A(KEYINPUT25), .B(KEYINPUT99), .ZN(n443) );
  XNOR2_X1 U328 ( .A(n444), .B(n443), .ZN(n448) );
  XNOR2_X1 U329 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U330 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n471) );
  XNOR2_X1 U331 ( .A(n325), .B(n324), .ZN(n329) );
  XNOR2_X1 U332 ( .A(n472), .B(n471), .ZN(n549) );
  XNOR2_X1 U333 ( .A(n435), .B(n434), .ZN(n437) );
  XNOR2_X1 U334 ( .A(n456), .B(n455), .ZN(n520) );
  NOR2_X1 U335 ( .A1(n548), .A2(n565), .ZN(n592) );
  XOR2_X1 U336 ( .A(n466), .B(KEYINPUT41), .Z(n555) );
  XOR2_X1 U337 ( .A(n439), .B(n438), .Z(n569) );
  XNOR2_X1 U338 ( .A(n479), .B(KEYINPUT62), .ZN(n480) );
  XNOR2_X1 U339 ( .A(n458), .B(KEYINPUT104), .ZN(n459) );
  XNOR2_X1 U340 ( .A(n481), .B(n480), .ZN(G1355GAT) );
  XNOR2_X1 U341 ( .A(n460), .B(n459), .ZN(G1329GAT) );
  XOR2_X1 U342 ( .A(G15GAT), .B(G113GAT), .Z(n293) );
  XNOR2_X1 U343 ( .A(G141GAT), .B(G22GAT), .ZN(n292) );
  XNOR2_X1 U344 ( .A(n293), .B(n292), .ZN(n297) );
  XOR2_X1 U345 ( .A(KEYINPUT68), .B(KEYINPUT67), .Z(n295) );
  XNOR2_X1 U346 ( .A(G169GAT), .B(KEYINPUT29), .ZN(n294) );
  XNOR2_X1 U347 ( .A(n295), .B(n294), .ZN(n296) );
  XNOR2_X1 U348 ( .A(n297), .B(n296), .ZN(n309) );
  XNOR2_X1 U349 ( .A(G197GAT), .B(G36GAT), .ZN(n298) );
  XNOR2_X1 U350 ( .A(n298), .B(G50GAT), .ZN(n300) );
  XNOR2_X1 U351 ( .A(G1GAT), .B(KEYINPUT70), .ZN(n299) );
  XNOR2_X1 U352 ( .A(n299), .B(G8GAT), .ZN(n332) );
  XOR2_X1 U353 ( .A(n300), .B(n332), .Z(n307) );
  XOR2_X1 U354 ( .A(G29GAT), .B(KEYINPUT8), .Z(n302) );
  XNOR2_X1 U355 ( .A(KEYINPUT7), .B(KEYINPUT69), .ZN(n301) );
  XNOR2_X1 U356 ( .A(n302), .B(n301), .ZN(n350) );
  XOR2_X1 U357 ( .A(n350), .B(KEYINPUT30), .Z(n304) );
  NAND2_X1 U358 ( .A1(G229GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U359 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U360 ( .A(n305), .B(G43GAT), .ZN(n306) );
  XNOR2_X1 U361 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U362 ( .A(n309), .B(n308), .ZN(n583) );
  INV_X1 U363 ( .A(n583), .ZN(n536) );
  XNOR2_X1 U364 ( .A(G204GAT), .B(G92GAT), .ZN(n310) );
  XNOR2_X1 U365 ( .A(n310), .B(G64GAT), .ZN(n388) );
  XOR2_X1 U366 ( .A(G85GAT), .B(G57GAT), .Z(n368) );
  XNOR2_X1 U367 ( .A(n388), .B(n368), .ZN(n314) );
  INV_X1 U368 ( .A(n314), .ZN(n312) );
  AND2_X1 U369 ( .A1(G230GAT), .A2(G233GAT), .ZN(n313) );
  INV_X1 U370 ( .A(n313), .ZN(n311) );
  NAND2_X1 U371 ( .A1(n312), .A2(n311), .ZN(n316) );
  NAND2_X1 U372 ( .A1(n314), .A2(n313), .ZN(n315) );
  NAND2_X1 U373 ( .A1(n316), .A2(n315), .ZN(n317) );
  XOR2_X1 U374 ( .A(n317), .B(KEYINPUT31), .Z(n325) );
  XOR2_X1 U375 ( .A(G78GAT), .B(G148GAT), .Z(n319) );
  XNOR2_X1 U376 ( .A(G106GAT), .B(KEYINPUT74), .ZN(n318) );
  XNOR2_X1 U377 ( .A(n319), .B(n318), .ZN(n418) );
  XNOR2_X1 U378 ( .A(n418), .B(KEYINPUT33), .ZN(n323) );
  XOR2_X1 U379 ( .A(KEYINPUT75), .B(KEYINPUT32), .Z(n321) );
  XNOR2_X1 U380 ( .A(G176GAT), .B(KEYINPUT73), .ZN(n320) );
  XNOR2_X1 U381 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U382 ( .A(G99GAT), .B(G71GAT), .ZN(n326) );
  XNOR2_X1 U383 ( .A(n326), .B(G120GAT), .ZN(n422) );
  XNOR2_X1 U384 ( .A(KEYINPUT13), .B(KEYINPUT72), .ZN(n327) );
  XNOR2_X1 U385 ( .A(n327), .B(KEYINPUT71), .ZN(n343) );
  XNOR2_X1 U386 ( .A(n422), .B(n343), .ZN(n328) );
  XNOR2_X1 U387 ( .A(n329), .B(n328), .ZN(n587) );
  NOR2_X1 U388 ( .A1(n536), .A2(n587), .ZN(n488) );
  XOR2_X1 U389 ( .A(KEYINPUT14), .B(KEYINPUT80), .Z(n331) );
  XNOR2_X1 U390 ( .A(KEYINPUT79), .B(KEYINPUT78), .ZN(n330) );
  XNOR2_X1 U391 ( .A(n331), .B(n330), .ZN(n336) );
  XOR2_X1 U392 ( .A(G22GAT), .B(G155GAT), .Z(n408) );
  XOR2_X1 U393 ( .A(n408), .B(n332), .Z(n334) );
  NAND2_X1 U394 ( .A1(G231GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U395 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U396 ( .A(n336), .B(n335), .ZN(n347) );
  XOR2_X1 U397 ( .A(G64GAT), .B(G57GAT), .Z(n338) );
  XNOR2_X1 U398 ( .A(G211GAT), .B(G78GAT), .ZN(n337) );
  XNOR2_X1 U399 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U400 ( .A(n339), .B(G71GAT), .Z(n341) );
  XOR2_X1 U401 ( .A(G15GAT), .B(G127GAT), .Z(n432) );
  XNOR2_X1 U402 ( .A(G183GAT), .B(n432), .ZN(n340) );
  XNOR2_X1 U403 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U404 ( .A(n342), .B(KEYINPUT12), .Z(n345) );
  XNOR2_X1 U405 ( .A(n343), .B(KEYINPUT15), .ZN(n344) );
  XNOR2_X1 U406 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U407 ( .A(n347), .B(n346), .ZN(n591) );
  INV_X1 U408 ( .A(n591), .ZN(n541) );
  XOR2_X1 U409 ( .A(KEYINPUT77), .B(G85GAT), .Z(n349) );
  XNOR2_X1 U410 ( .A(G218GAT), .B(G106GAT), .ZN(n348) );
  XNOR2_X1 U411 ( .A(n349), .B(n348), .ZN(n354) );
  XOR2_X1 U412 ( .A(G36GAT), .B(G190GAT), .Z(n389) );
  XOR2_X1 U413 ( .A(n350), .B(n389), .Z(n352) );
  NAND2_X1 U414 ( .A1(G232GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U415 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U416 ( .A(n354), .B(n353), .Z(n356) );
  XOR2_X1 U417 ( .A(G43GAT), .B(G134GAT), .Z(n423) );
  XOR2_X1 U418 ( .A(G50GAT), .B(G162GAT), .Z(n409) );
  XNOR2_X1 U419 ( .A(n423), .B(n409), .ZN(n355) );
  XNOR2_X1 U420 ( .A(n356), .B(n355), .ZN(n364) );
  XOR2_X1 U421 ( .A(KEYINPUT11), .B(KEYINPUT65), .Z(n358) );
  XNOR2_X1 U422 ( .A(G92GAT), .B(KEYINPUT9), .ZN(n357) );
  XNOR2_X1 U423 ( .A(n358), .B(n357), .ZN(n362) );
  XOR2_X1 U424 ( .A(KEYINPUT76), .B(KEYINPUT66), .Z(n360) );
  XNOR2_X1 U425 ( .A(G99GAT), .B(KEYINPUT10), .ZN(n359) );
  XNOR2_X1 U426 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U427 ( .A(n362), .B(n361), .Z(n363) );
  XNOR2_X1 U428 ( .A(n364), .B(n363), .ZN(n562) );
  XNOR2_X1 U429 ( .A(KEYINPUT36), .B(n562), .ZN(n478) );
  XOR2_X1 U430 ( .A(G155GAT), .B(G162GAT), .Z(n366) );
  XNOR2_X1 U431 ( .A(G134GAT), .B(G148GAT), .ZN(n365) );
  XNOR2_X1 U432 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U433 ( .A(n367), .B(KEYINPUT77), .Z(n370) );
  XNOR2_X1 U434 ( .A(G29GAT), .B(n368), .ZN(n369) );
  XNOR2_X1 U435 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U436 ( .A(KEYINPUT94), .B(KEYINPUT6), .Z(n372) );
  XNOR2_X1 U437 ( .A(KEYINPUT5), .B(KEYINPUT91), .ZN(n371) );
  XNOR2_X1 U438 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U439 ( .A(n374), .B(n373), .ZN(n378) );
  XOR2_X1 U440 ( .A(KEYINPUT4), .B(G120GAT), .Z(n376) );
  XNOR2_X1 U441 ( .A(G1GAT), .B(G127GAT), .ZN(n375) );
  XNOR2_X1 U442 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U443 ( .A(n378), .B(n377), .ZN(n387) );
  XOR2_X1 U444 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n380) );
  NAND2_X1 U445 ( .A1(G225GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U446 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U447 ( .A(n381), .B(KEYINPUT1), .Z(n385) );
  XNOR2_X1 U448 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n382) );
  XNOR2_X1 U449 ( .A(n382), .B(KEYINPUT83), .ZN(n431) );
  XNOR2_X1 U450 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n383) );
  XNOR2_X1 U451 ( .A(n383), .B(KEYINPUT2), .ZN(n416) );
  XNOR2_X1 U452 ( .A(n431), .B(n416), .ZN(n384) );
  XNOR2_X1 U453 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U454 ( .A(n387), .B(n386), .ZN(n521) );
  XOR2_X1 U455 ( .A(n389), .B(n388), .Z(n391) );
  NAND2_X1 U456 ( .A1(G226GAT), .A2(G233GAT), .ZN(n390) );
  XNOR2_X1 U457 ( .A(n391), .B(n390), .ZN(n395) );
  XOR2_X1 U458 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n393) );
  XNOR2_X1 U459 ( .A(G8GAT), .B(KEYINPUT95), .ZN(n392) );
  XNOR2_X1 U460 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U461 ( .A(n395), .B(n394), .Z(n405) );
  XOR2_X1 U462 ( .A(KEYINPUT85), .B(KEYINPUT17), .Z(n397) );
  XNOR2_X1 U463 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n396) );
  XNOR2_X1 U464 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U465 ( .A(n398), .B(G183GAT), .Z(n400) );
  XNOR2_X1 U466 ( .A(G169GAT), .B(G176GAT), .ZN(n399) );
  XNOR2_X1 U467 ( .A(n400), .B(n399), .ZN(n439) );
  XOR2_X1 U468 ( .A(KEYINPUT90), .B(G218GAT), .Z(n402) );
  XNOR2_X1 U469 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n401) );
  XNOR2_X1 U470 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U471 ( .A(G197GAT), .B(n403), .Z(n419) );
  XNOR2_X1 U472 ( .A(n439), .B(n419), .ZN(n404) );
  XNOR2_X1 U473 ( .A(n405), .B(n404), .ZN(n525) );
  XNOR2_X1 U474 ( .A(n525), .B(KEYINPUT27), .ZN(n446) );
  NOR2_X1 U475 ( .A1(n521), .A2(n446), .ZN(n551) );
  XOR2_X1 U476 ( .A(G204GAT), .B(KEYINPUT23), .Z(n407) );
  XNOR2_X1 U477 ( .A(KEYINPUT89), .B(KEYINPUT88), .ZN(n406) );
  XNOR2_X1 U478 ( .A(n407), .B(n406), .ZN(n413) );
  XOR2_X1 U479 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n411) );
  XNOR2_X1 U480 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U481 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U482 ( .A(n413), .B(n412), .Z(n415) );
  NAND2_X1 U483 ( .A1(G228GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U484 ( .A(n415), .B(n414), .ZN(n417) );
  XOR2_X1 U485 ( .A(n417), .B(n416), .Z(n421) );
  XNOR2_X1 U486 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U487 ( .A(n421), .B(n420), .ZN(n566) );
  XOR2_X1 U488 ( .A(n566), .B(KEYINPUT28), .Z(n529) );
  NAND2_X1 U489 ( .A1(n551), .A2(n529), .ZN(n533) );
  XNOR2_X1 U490 ( .A(n423), .B(n422), .ZN(n427) );
  INV_X1 U491 ( .A(n427), .ZN(n425) );
  AND2_X1 U492 ( .A1(G227GAT), .A2(G233GAT), .ZN(n426) );
  INV_X1 U493 ( .A(n426), .ZN(n424) );
  NAND2_X1 U494 ( .A1(n425), .A2(n424), .ZN(n429) );
  NAND2_X1 U495 ( .A1(n427), .A2(n426), .ZN(n428) );
  NAND2_X1 U496 ( .A1(n429), .A2(n428), .ZN(n430) );
  XNOR2_X1 U497 ( .A(n430), .B(KEYINPUT20), .ZN(n435) );
  XOR2_X1 U498 ( .A(KEYINPUT84), .B(n431), .Z(n433) );
  XOR2_X1 U499 ( .A(G190GAT), .B(KEYINPUT86), .Z(n436) );
  XNOR2_X1 U500 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U501 ( .A(KEYINPUT87), .B(n569), .ZN(n440) );
  NOR2_X1 U502 ( .A1(n533), .A2(n440), .ZN(n452) );
  NOR2_X1 U503 ( .A1(n569), .A2(n525), .ZN(n441) );
  XNOR2_X1 U504 ( .A(n441), .B(KEYINPUT98), .ZN(n442) );
  NOR2_X1 U505 ( .A1(n566), .A2(n442), .ZN(n444) );
  NAND2_X1 U506 ( .A1(n566), .A2(n569), .ZN(n445) );
  XNOR2_X1 U507 ( .A(n445), .B(KEYINPUT26), .ZN(n548) );
  NOR2_X1 U508 ( .A1(n548), .A2(n446), .ZN(n447) );
  NOR2_X1 U509 ( .A1(n448), .A2(n447), .ZN(n450) );
  INV_X1 U510 ( .A(n521), .ZN(n449) );
  NOR2_X1 U511 ( .A1(n450), .A2(n449), .ZN(n451) );
  NOR2_X1 U512 ( .A1(n452), .A2(n451), .ZN(n486) );
  NOR2_X1 U513 ( .A1(n478), .A2(n486), .ZN(n453) );
  NAND2_X1 U514 ( .A1(n541), .A2(n453), .ZN(n456) );
  INV_X1 U515 ( .A(KEYINPUT37), .ZN(n454) );
  NAND2_X1 U516 ( .A1(n488), .A2(n520), .ZN(n457) );
  NOR2_X1 U517 ( .A1(n504), .A2(n525), .ZN(n460) );
  INV_X1 U518 ( .A(G36GAT), .ZN(n458) );
  INV_X1 U519 ( .A(n587), .ZN(n466) );
  NOR2_X1 U520 ( .A1(n555), .A2(n536), .ZN(n461) );
  XNOR2_X1 U521 ( .A(n461), .B(KEYINPUT46), .ZN(n462) );
  NOR2_X1 U522 ( .A1(n591), .A2(n462), .ZN(n463) );
  NAND2_X1 U523 ( .A1(n463), .A2(n562), .ZN(n464) );
  XNOR2_X1 U524 ( .A(n464), .B(KEYINPUT47), .ZN(n470) );
  NOR2_X1 U525 ( .A1(n478), .A2(n541), .ZN(n465) );
  XNOR2_X1 U526 ( .A(KEYINPUT45), .B(n465), .ZN(n467) );
  NAND2_X1 U527 ( .A1(n467), .A2(n466), .ZN(n468) );
  NOR2_X1 U528 ( .A1(n468), .A2(n583), .ZN(n469) );
  NOR2_X1 U529 ( .A1(n470), .A2(n469), .ZN(n472) );
  XOR2_X1 U530 ( .A(KEYINPUT121), .B(n525), .Z(n473) );
  NOR2_X1 U531 ( .A1(n549), .A2(n473), .ZN(n474) );
  XNOR2_X1 U532 ( .A(KEYINPUT122), .B(n474), .ZN(n475) );
  XNOR2_X1 U533 ( .A(n475), .B(KEYINPUT54), .ZN(n476) );
  NAND2_X1 U534 ( .A1(n476), .A2(n521), .ZN(n565) );
  INV_X1 U535 ( .A(n592), .ZN(n477) );
  NOR2_X1 U536 ( .A1(n478), .A2(n477), .ZN(n481) );
  INV_X1 U537 ( .A(G218GAT), .ZN(n479) );
  XOR2_X1 U538 ( .A(KEYINPUT16), .B(KEYINPUT82), .Z(n483) );
  NAND2_X1 U539 ( .A1(n591), .A2(n562), .ZN(n482) );
  XNOR2_X1 U540 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U541 ( .A(n484), .B(KEYINPUT81), .ZN(n485) );
  NOR2_X1 U542 ( .A1(n486), .A2(n485), .ZN(n487) );
  XNOR2_X1 U543 ( .A(KEYINPUT100), .B(n487), .ZN(n508) );
  NAND2_X1 U544 ( .A1(n488), .A2(n508), .ZN(n496) );
  NOR2_X1 U545 ( .A1(n521), .A2(n496), .ZN(n490) );
  XNOR2_X1 U546 ( .A(KEYINPUT34), .B(KEYINPUT101), .ZN(n489) );
  XNOR2_X1 U547 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U548 ( .A(G1GAT), .B(n491), .ZN(G1324GAT) );
  NOR2_X1 U549 ( .A1(n525), .A2(n496), .ZN(n492) );
  XOR2_X1 U550 ( .A(G8GAT), .B(n492), .Z(G1325GAT) );
  NOR2_X1 U551 ( .A1(n569), .A2(n496), .ZN(n494) );
  XNOR2_X1 U552 ( .A(KEYINPUT102), .B(KEYINPUT35), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U554 ( .A(G15GAT), .B(n495), .ZN(G1326GAT) );
  NOR2_X1 U555 ( .A1(n529), .A2(n496), .ZN(n497) );
  XOR2_X1 U556 ( .A(G22GAT), .B(n497), .Z(G1327GAT) );
  NOR2_X1 U557 ( .A1(n504), .A2(n521), .ZN(n498) );
  XNOR2_X1 U558 ( .A(n498), .B(KEYINPUT39), .ZN(n499) );
  XNOR2_X1 U559 ( .A(G29GAT), .B(n499), .ZN(G1328GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n501) );
  XNOR2_X1 U561 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n501), .B(n500), .ZN(n503) );
  NOR2_X1 U563 ( .A1(n569), .A2(n504), .ZN(n502) );
  XOR2_X1 U564 ( .A(n503), .B(n502), .Z(G1330GAT) );
  XNOR2_X1 U565 ( .A(G50GAT), .B(KEYINPUT107), .ZN(n506) );
  NOR2_X1 U566 ( .A1(n529), .A2(n504), .ZN(n505) );
  XNOR2_X1 U567 ( .A(n506), .B(n505), .ZN(G1331GAT) );
  NOR2_X1 U568 ( .A1(n555), .A2(n583), .ZN(n507) );
  XNOR2_X1 U569 ( .A(n507), .B(KEYINPUT108), .ZN(n519) );
  NAND2_X1 U570 ( .A1(n508), .A2(n519), .ZN(n515) );
  NOR2_X1 U571 ( .A1(n521), .A2(n515), .ZN(n509) );
  XOR2_X1 U572 ( .A(n509), .B(KEYINPUT42), .Z(n510) );
  XNOR2_X1 U573 ( .A(G57GAT), .B(n510), .ZN(G1332GAT) );
  NOR2_X1 U574 ( .A1(n525), .A2(n515), .ZN(n511) );
  XOR2_X1 U575 ( .A(G64GAT), .B(n511), .Z(G1333GAT) );
  NOR2_X1 U576 ( .A1(n569), .A2(n515), .ZN(n513) );
  XNOR2_X1 U577 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n512) );
  XNOR2_X1 U578 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U579 ( .A(G71GAT), .B(n514), .ZN(G1334GAT) );
  NOR2_X1 U580 ( .A1(n529), .A2(n515), .ZN(n517) );
  XNOR2_X1 U581 ( .A(KEYINPUT43), .B(KEYINPUT111), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n517), .B(n516), .ZN(n518) );
  XOR2_X1 U583 ( .A(G78GAT), .B(n518), .Z(G1335GAT) );
  NAND2_X1 U584 ( .A1(n520), .A2(n519), .ZN(n528) );
  NOR2_X1 U585 ( .A1(n521), .A2(n528), .ZN(n523) );
  XNOR2_X1 U586 ( .A(KEYINPUT112), .B(KEYINPUT113), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U588 ( .A(G85GAT), .B(n524), .ZN(G1336GAT) );
  NOR2_X1 U589 ( .A1(n525), .A2(n528), .ZN(n526) );
  XOR2_X1 U590 ( .A(G92GAT), .B(n526), .Z(G1337GAT) );
  NOR2_X1 U591 ( .A1(n569), .A2(n528), .ZN(n527) );
  XOR2_X1 U592 ( .A(G99GAT), .B(n527), .Z(G1338GAT) );
  NOR2_X1 U593 ( .A1(n529), .A2(n528), .ZN(n531) );
  XNOR2_X1 U594 ( .A(KEYINPUT114), .B(KEYINPUT44), .ZN(n530) );
  XNOR2_X1 U595 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U596 ( .A(G106GAT), .B(n532), .Z(G1339GAT) );
  NOR2_X1 U597 ( .A1(n549), .A2(n533), .ZN(n535) );
  INV_X1 U598 ( .A(n569), .ZN(n534) );
  NAND2_X1 U599 ( .A1(n535), .A2(n534), .ZN(n545) );
  NOR2_X1 U600 ( .A1(n536), .A2(n545), .ZN(n538) );
  XNOR2_X1 U601 ( .A(G113GAT), .B(KEYINPUT115), .ZN(n537) );
  XNOR2_X1 U602 ( .A(n538), .B(n537), .ZN(G1340GAT) );
  NOR2_X1 U603 ( .A1(n555), .A2(n545), .ZN(n540) );
  XNOR2_X1 U604 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n540), .B(n539), .ZN(G1341GAT) );
  NOR2_X1 U606 ( .A1(n541), .A2(n545), .ZN(n543) );
  XNOR2_X1 U607 ( .A(KEYINPUT50), .B(KEYINPUT116), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U609 ( .A(G127GAT), .B(n544), .Z(G1342GAT) );
  NOR2_X1 U610 ( .A1(n562), .A2(n545), .ZN(n547) );
  XNOR2_X1 U611 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n547), .B(n546), .ZN(G1343GAT) );
  NOR2_X1 U613 ( .A1(n549), .A2(n548), .ZN(n550) );
  NAND2_X1 U614 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U615 ( .A(KEYINPUT117), .B(n552), .ZN(n563) );
  NAND2_X1 U616 ( .A1(n563), .A2(n583), .ZN(n553) );
  XNOR2_X1 U617 ( .A(n553), .B(KEYINPUT118), .ZN(n554) );
  XNOR2_X1 U618 ( .A(G141GAT), .B(n554), .ZN(G1344GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT52), .B(KEYINPUT119), .Z(n557) );
  INV_X1 U620 ( .A(n555), .ZN(n574) );
  NAND2_X1 U621 ( .A1(n563), .A2(n574), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n557), .B(n556), .ZN(n559) );
  XOR2_X1 U623 ( .A(G148GAT), .B(KEYINPUT53), .Z(n558) );
  XNOR2_X1 U624 ( .A(n559), .B(n558), .ZN(G1345GAT) );
  NAND2_X1 U625 ( .A1(n563), .A2(n591), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(KEYINPUT120), .ZN(n561) );
  XNOR2_X1 U627 ( .A(G155GAT), .B(n561), .ZN(G1346GAT) );
  INV_X1 U628 ( .A(n562), .ZN(n580) );
  NAND2_X1 U629 ( .A1(n563), .A2(n580), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U632 ( .A(n567), .B(KEYINPUT55), .ZN(n568) );
  NOR2_X1 U633 ( .A1(n569), .A2(n568), .ZN(n579) );
  NAND2_X1 U634 ( .A1(n583), .A2(n579), .ZN(n570) );
  XNOR2_X1 U635 ( .A(G169GAT), .B(n570), .ZN(G1348GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT57), .B(KEYINPUT124), .Z(n572) );
  XNOR2_X1 U637 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XOR2_X1 U639 ( .A(KEYINPUT123), .B(n573), .Z(n576) );
  NAND2_X1 U640 ( .A1(n579), .A2(n574), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1349GAT) );
  XOR2_X1 U642 ( .A(G183GAT), .B(KEYINPUT125), .Z(n578) );
  NAND2_X1 U643 ( .A1(n579), .A2(n591), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(G1350GAT) );
  XNOR2_X1 U645 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n582) );
  NAND2_X1 U646 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1351GAT) );
  XOR2_X1 U648 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n585) );
  NAND2_X1 U649 ( .A1(n592), .A2(n583), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(G197GAT), .B(n586), .ZN(G1352GAT) );
  XOR2_X1 U652 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n589) );
  NAND2_X1 U653 ( .A1(n592), .A2(n587), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U655 ( .A(G204GAT), .B(n590), .ZN(G1353GAT) );
  NAND2_X1 U656 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U657 ( .A(n593), .B(G211GAT), .ZN(G1354GAT) );
endmodule

