

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U556 ( .A1(n599), .A2(n598), .ZN(n989) );
  NOR2_X2 U557 ( .A1(n597), .A2(n596), .ZN(n599) );
  OR2_X1 U558 ( .A1(n790), .A2(n789), .ZN(n791) );
  BUF_X1 U559 ( .A(n763), .Z(n779) );
  NOR2_X4 U560 ( .A1(G651), .A2(n651), .ZN(n662) );
  NOR2_X2 U561 ( .A1(G1384), .A2(G164), .ZN(n724) );
  NOR2_X4 U562 ( .A1(G2105), .A2(n531), .ZN(n566) );
  INV_X2 U563 ( .A(G2104), .ZN(n531) );
  NAND2_X1 U564 ( .A1(n528), .A2(n531), .ZN(n529) );
  INV_X1 U565 ( .A(G2105), .ZN(n528) );
  XOR2_X1 U566 ( .A(n762), .B(KEYINPUT29), .Z(n523) );
  AND2_X1 U567 ( .A1(G138), .A2(n900), .ZN(n524) );
  NOR2_X1 U568 ( .A1(n813), .A2(n812), .ZN(n525) );
  AND2_X1 U569 ( .A1(n814), .A2(n525), .ZN(n526) );
  NAND2_X1 U570 ( .A1(n772), .A2(n788), .ZN(n527) );
  INV_X1 U571 ( .A(n977), .ZN(n812) );
  AND2_X1 U572 ( .A1(n777), .A2(n776), .ZN(n778) );
  NAND2_X1 U573 ( .A1(n527), .A2(n778), .ZN(n797) );
  XOR2_X1 U574 ( .A(KEYINPUT83), .B(n530), .Z(n533) );
  XOR2_X1 U575 ( .A(KEYINPUT1), .B(n549), .Z(n668) );
  AND2_X1 U576 ( .A1(G2105), .A2(G2104), .ZN(n896) );
  NAND2_X1 U577 ( .A1(n896), .A2(G114), .ZN(n536) );
  XNOR2_X2 U578 ( .A(n529), .B(KEYINPUT17), .ZN(n900) );
  NAND2_X1 U579 ( .A1(G102), .A2(n566), .ZN(n530) );
  AND2_X1 U580 ( .A1(n531), .A2(G2105), .ZN(n570) );
  NAND2_X1 U581 ( .A1(G126), .A2(n570), .ZN(n532) );
  NAND2_X1 U582 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X1 U583 ( .A1(n524), .A2(n534), .ZN(n535) );
  NAND2_X1 U584 ( .A1(n536), .A2(n535), .ZN(n538) );
  INV_X1 U585 ( .A(KEYINPUT84), .ZN(n537) );
  XNOR2_X2 U586 ( .A(n538), .B(n537), .ZN(G164) );
  XOR2_X1 U587 ( .A(G2427), .B(G2435), .Z(n540) );
  XNOR2_X1 U588 ( .A(G2454), .B(G2443), .ZN(n539) );
  XNOR2_X1 U589 ( .A(n540), .B(n539), .ZN(n547) );
  XOR2_X1 U590 ( .A(G2451), .B(KEYINPUT101), .Z(n542) );
  XNOR2_X1 U591 ( .A(G2430), .B(G2438), .ZN(n541) );
  XNOR2_X1 U592 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U593 ( .A(n543), .B(G2446), .Z(n545) );
  XNOR2_X1 U594 ( .A(G1341), .B(G1348), .ZN(n544) );
  XNOR2_X1 U595 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U596 ( .A(n547), .B(n546), .ZN(n548) );
  AND2_X1 U597 ( .A1(n548), .A2(G14), .ZN(G401) );
  INV_X1 U598 ( .A(G57), .ZN(G237) );
  INV_X1 U599 ( .A(G132), .ZN(G219) );
  INV_X1 U600 ( .A(G82), .ZN(G220) );
  INV_X1 U601 ( .A(G651), .ZN(n552) );
  NOR2_X1 U602 ( .A1(G543), .A2(n552), .ZN(n549) );
  NAND2_X1 U603 ( .A1(G64), .A2(n668), .ZN(n550) );
  XNOR2_X1 U604 ( .A(n550), .B(KEYINPUT67), .ZN(n559) );
  NOR2_X1 U605 ( .A1(G651), .A2(G543), .ZN(n663) );
  NAND2_X1 U606 ( .A1(G90), .A2(n663), .ZN(n554) );
  XNOR2_X1 U607 ( .A(G543), .B(KEYINPUT0), .ZN(n551) );
  XNOR2_X1 U608 ( .A(n551), .B(KEYINPUT65), .ZN(n651) );
  NOR2_X1 U609 ( .A1(n651), .A2(n552), .ZN(n664) );
  NAND2_X1 U610 ( .A1(G77), .A2(n664), .ZN(n553) );
  NAND2_X1 U611 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U612 ( .A(n555), .B(KEYINPUT9), .ZN(n557) );
  NAND2_X1 U613 ( .A1(G52), .A2(n662), .ZN(n556) );
  NAND2_X1 U614 ( .A1(n557), .A2(n556), .ZN(n558) );
  NOR2_X1 U615 ( .A1(n559), .A2(n558), .ZN(G171) );
  NAND2_X1 U616 ( .A1(G88), .A2(n663), .ZN(n561) );
  NAND2_X1 U617 ( .A1(G75), .A2(n664), .ZN(n560) );
  NAND2_X1 U618 ( .A1(n561), .A2(n560), .ZN(n565) );
  NAND2_X1 U619 ( .A1(G62), .A2(n668), .ZN(n563) );
  NAND2_X1 U620 ( .A1(G50), .A2(n662), .ZN(n562) );
  NAND2_X1 U621 ( .A1(n563), .A2(n562), .ZN(n564) );
  NOR2_X1 U622 ( .A1(n565), .A2(n564), .ZN(G166) );
  NAND2_X1 U623 ( .A1(n900), .A2(G137), .ZN(n569) );
  NAND2_X1 U624 ( .A1(G101), .A2(n566), .ZN(n567) );
  XOR2_X1 U625 ( .A(KEYINPUT23), .B(n567), .Z(n568) );
  NAND2_X1 U626 ( .A1(n569), .A2(n568), .ZN(n574) );
  NAND2_X1 U627 ( .A1(G125), .A2(n570), .ZN(n572) );
  NAND2_X1 U628 ( .A1(G113), .A2(n896), .ZN(n571) );
  NAND2_X1 U629 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U630 ( .A1(n574), .A2(n573), .ZN(G160) );
  XNOR2_X1 U631 ( .A(KEYINPUT74), .B(KEYINPUT7), .ZN(n586) );
  NAND2_X1 U632 ( .A1(n663), .A2(G89), .ZN(n575) );
  XNOR2_X1 U633 ( .A(n575), .B(KEYINPUT4), .ZN(n577) );
  NAND2_X1 U634 ( .A1(G76), .A2(n664), .ZN(n576) );
  NAND2_X1 U635 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U636 ( .A(KEYINPUT5), .B(n578), .ZN(n584) );
  NAND2_X1 U637 ( .A1(n668), .A2(G63), .ZN(n579) );
  XOR2_X1 U638 ( .A(KEYINPUT73), .B(n579), .Z(n581) );
  NAND2_X1 U639 ( .A1(n662), .A2(G51), .ZN(n580) );
  NAND2_X1 U640 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U641 ( .A(KEYINPUT6), .B(n582), .Z(n583) );
  NAND2_X1 U642 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U643 ( .A(n586), .B(n585), .ZN(G168) );
  XOR2_X1 U644 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U645 ( .A1(G94), .A2(G452), .ZN(n587) );
  XOR2_X1 U646 ( .A(KEYINPUT68), .B(n587), .Z(G173) );
  NAND2_X1 U647 ( .A1(G7), .A2(G661), .ZN(n588) );
  XNOR2_X1 U648 ( .A(n588), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U649 ( .A(G223), .ZN(n842) );
  NAND2_X1 U650 ( .A1(n842), .A2(G567), .ZN(n589) );
  XOR2_X1 U651 ( .A(KEYINPUT11), .B(n589), .Z(G234) );
  NAND2_X1 U652 ( .A1(n663), .A2(G81), .ZN(n590) );
  XNOR2_X1 U653 ( .A(n590), .B(KEYINPUT12), .ZN(n592) );
  NAND2_X1 U654 ( .A1(G68), .A2(n664), .ZN(n591) );
  NAND2_X1 U655 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U656 ( .A(KEYINPUT13), .B(n593), .Z(n597) );
  NAND2_X1 U657 ( .A1(G56), .A2(n668), .ZN(n594) );
  XNOR2_X1 U658 ( .A(n594), .B(KEYINPUT14), .ZN(n595) );
  XNOR2_X1 U659 ( .A(n595), .B(KEYINPUT71), .ZN(n596) );
  NAND2_X1 U660 ( .A1(n662), .A2(G43), .ZN(n598) );
  INV_X1 U661 ( .A(G860), .ZN(n621) );
  OR2_X1 U662 ( .A1(n989), .A2(n621), .ZN(G153) );
  INV_X1 U663 ( .A(G171), .ZN(G301) );
  NAND2_X1 U664 ( .A1(G868), .A2(G301), .ZN(n609) );
  NAND2_X1 U665 ( .A1(G79), .A2(n664), .ZN(n606) );
  NAND2_X1 U666 ( .A1(G66), .A2(n668), .ZN(n601) );
  NAND2_X1 U667 ( .A1(G92), .A2(n663), .ZN(n600) );
  NAND2_X1 U668 ( .A1(n601), .A2(n600), .ZN(n604) );
  NAND2_X1 U669 ( .A1(n662), .A2(G54), .ZN(n602) );
  XOR2_X1 U670 ( .A(KEYINPUT72), .B(n602), .Z(n603) );
  NOR2_X1 U671 ( .A1(n604), .A2(n603), .ZN(n605) );
  NAND2_X1 U672 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X2 U673 ( .A(n607), .B(KEYINPUT15), .ZN(n988) );
  INV_X1 U674 ( .A(G868), .ZN(n679) );
  NAND2_X1 U675 ( .A1(n736), .A2(n679), .ZN(n608) );
  NAND2_X1 U676 ( .A1(n609), .A2(n608), .ZN(G284) );
  NAND2_X1 U677 ( .A1(G91), .A2(n663), .ZN(n611) );
  NAND2_X1 U678 ( .A1(G78), .A2(n664), .ZN(n610) );
  NAND2_X1 U679 ( .A1(n611), .A2(n610), .ZN(n616) );
  NAND2_X1 U680 ( .A1(G65), .A2(n668), .ZN(n613) );
  NAND2_X1 U681 ( .A1(G53), .A2(n662), .ZN(n612) );
  NAND2_X1 U682 ( .A1(n613), .A2(n612), .ZN(n614) );
  XOR2_X1 U683 ( .A(KEYINPUT69), .B(n614), .Z(n615) );
  NOR2_X1 U684 ( .A1(n616), .A2(n615), .ZN(n617) );
  XOR2_X1 U685 ( .A(KEYINPUT70), .B(n617), .Z(G299) );
  NOR2_X1 U686 ( .A1(G286), .A2(n679), .ZN(n618) );
  XOR2_X1 U687 ( .A(KEYINPUT75), .B(n618), .Z(n620) );
  NOR2_X1 U688 ( .A1(G299), .A2(G868), .ZN(n619) );
  NOR2_X1 U689 ( .A1(n620), .A2(n619), .ZN(G297) );
  NAND2_X1 U690 ( .A1(n621), .A2(G559), .ZN(n622) );
  NAND2_X1 U691 ( .A1(n622), .A2(n988), .ZN(n623) );
  XNOR2_X1 U692 ( .A(n623), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U693 ( .A1(G868), .A2(n989), .ZN(n624) );
  XNOR2_X1 U694 ( .A(KEYINPUT76), .B(n624), .ZN(n627) );
  NAND2_X1 U695 ( .A1(G868), .A2(n988), .ZN(n625) );
  NOR2_X1 U696 ( .A1(G559), .A2(n625), .ZN(n626) );
  NOR2_X1 U697 ( .A1(n627), .A2(n626), .ZN(G282) );
  NAND2_X1 U698 ( .A1(G123), .A2(n570), .ZN(n628) );
  XNOR2_X1 U699 ( .A(n628), .B(KEYINPUT18), .ZN(n630) );
  BUF_X1 U700 ( .A(n566), .Z(n899) );
  NAND2_X1 U701 ( .A1(n899), .A2(G99), .ZN(n629) );
  NAND2_X1 U702 ( .A1(n630), .A2(n629), .ZN(n634) );
  NAND2_X1 U703 ( .A1(G135), .A2(n900), .ZN(n632) );
  NAND2_X1 U704 ( .A1(G111), .A2(n896), .ZN(n631) );
  NAND2_X1 U705 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U706 ( .A1(n634), .A2(n633), .ZN(n1008) );
  XNOR2_X1 U707 ( .A(n1008), .B(G2096), .ZN(n636) );
  INV_X1 U708 ( .A(G2100), .ZN(n635) );
  NAND2_X1 U709 ( .A1(n636), .A2(n635), .ZN(G156) );
  NAND2_X1 U710 ( .A1(G61), .A2(n668), .ZN(n638) );
  NAND2_X1 U711 ( .A1(G86), .A2(n663), .ZN(n637) );
  NAND2_X1 U712 ( .A1(n638), .A2(n637), .ZN(n641) );
  NAND2_X1 U713 ( .A1(n664), .A2(G73), .ZN(n639) );
  XOR2_X1 U714 ( .A(KEYINPUT2), .B(n639), .Z(n640) );
  NOR2_X1 U715 ( .A1(n641), .A2(n640), .ZN(n643) );
  NAND2_X1 U716 ( .A1(n662), .A2(G48), .ZN(n642) );
  NAND2_X1 U717 ( .A1(n643), .A2(n642), .ZN(G305) );
  NAND2_X1 U718 ( .A1(n662), .A2(G47), .ZN(n645) );
  NAND2_X1 U719 ( .A1(n668), .A2(G60), .ZN(n644) );
  NAND2_X1 U720 ( .A1(n645), .A2(n644), .ZN(n646) );
  XOR2_X1 U721 ( .A(KEYINPUT66), .B(n646), .Z(n650) );
  NAND2_X1 U722 ( .A1(G85), .A2(n663), .ZN(n648) );
  NAND2_X1 U723 ( .A1(G72), .A2(n664), .ZN(n647) );
  AND2_X1 U724 ( .A1(n648), .A2(n647), .ZN(n649) );
  NAND2_X1 U725 ( .A1(n650), .A2(n649), .ZN(G290) );
  NAND2_X1 U726 ( .A1(G49), .A2(n662), .ZN(n653) );
  NAND2_X1 U727 ( .A1(G87), .A2(n651), .ZN(n652) );
  NAND2_X1 U728 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U729 ( .A1(n668), .A2(n654), .ZN(n656) );
  NAND2_X1 U730 ( .A1(G651), .A2(G74), .ZN(n655) );
  NAND2_X1 U731 ( .A1(n656), .A2(n655), .ZN(G288) );
  XNOR2_X1 U732 ( .A(KEYINPUT81), .B(KEYINPUT19), .ZN(n658) );
  XOR2_X1 U733 ( .A(G290), .B(G288), .Z(n657) );
  XNOR2_X1 U734 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U735 ( .A(G305), .B(n659), .ZN(n661) );
  XNOR2_X1 U736 ( .A(G166), .B(G299), .ZN(n660) );
  XNOR2_X1 U737 ( .A(n661), .B(n660), .ZN(n675) );
  NAND2_X1 U738 ( .A1(n662), .A2(G55), .ZN(n673) );
  NAND2_X1 U739 ( .A1(G93), .A2(n663), .ZN(n666) );
  NAND2_X1 U740 ( .A1(G80), .A2(n664), .ZN(n665) );
  NAND2_X1 U741 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U742 ( .A(KEYINPUT78), .B(n667), .ZN(n671) );
  NAND2_X1 U743 ( .A1(G67), .A2(n668), .ZN(n669) );
  XNOR2_X1 U744 ( .A(KEYINPUT79), .B(n669), .ZN(n670) );
  NOR2_X1 U745 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U746 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U747 ( .A(KEYINPUT80), .B(n674), .ZN(n853) );
  XOR2_X1 U748 ( .A(n675), .B(n853), .Z(n856) );
  NAND2_X1 U749 ( .A1(G559), .A2(n988), .ZN(n676) );
  XOR2_X1 U750 ( .A(n989), .B(n676), .Z(n851) );
  XNOR2_X1 U751 ( .A(n856), .B(n851), .ZN(n677) );
  NAND2_X1 U752 ( .A1(n677), .A2(G868), .ZN(n678) );
  XNOR2_X1 U753 ( .A(n678), .B(KEYINPUT82), .ZN(n681) );
  NAND2_X1 U754 ( .A1(n853), .A2(n679), .ZN(n680) );
  NAND2_X1 U755 ( .A1(n681), .A2(n680), .ZN(G295) );
  NAND2_X1 U756 ( .A1(G2078), .A2(G2084), .ZN(n682) );
  XOR2_X1 U757 ( .A(KEYINPUT20), .B(n682), .Z(n683) );
  NAND2_X1 U758 ( .A1(G2090), .A2(n683), .ZN(n684) );
  XNOR2_X1 U759 ( .A(KEYINPUT21), .B(n684), .ZN(n685) );
  NAND2_X1 U760 ( .A1(n685), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U761 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U762 ( .A1(G220), .A2(G219), .ZN(n686) );
  XOR2_X1 U763 ( .A(KEYINPUT22), .B(n686), .Z(n687) );
  NOR2_X1 U764 ( .A1(G218), .A2(n687), .ZN(n688) );
  NAND2_X1 U765 ( .A1(G96), .A2(n688), .ZN(n849) );
  NAND2_X1 U766 ( .A1(n849), .A2(G2106), .ZN(n692) );
  NAND2_X1 U767 ( .A1(G69), .A2(G120), .ZN(n689) );
  NOR2_X1 U768 ( .A1(G237), .A2(n689), .ZN(n690) );
  NAND2_X1 U769 ( .A1(G108), .A2(n690), .ZN(n850) );
  NAND2_X1 U770 ( .A1(n850), .A2(G567), .ZN(n691) );
  NAND2_X1 U771 ( .A1(n692), .A2(n691), .ZN(n928) );
  NAND2_X1 U772 ( .A1(G483), .A2(G661), .ZN(n693) );
  NOR2_X1 U773 ( .A1(n928), .A2(n693), .ZN(n847) );
  NAND2_X1 U774 ( .A1(n847), .A2(G36), .ZN(G176) );
  INV_X1 U775 ( .A(G166), .ZN(G303) );
  NAND2_X1 U776 ( .A1(G95), .A2(n899), .ZN(n695) );
  NAND2_X1 U777 ( .A1(G131), .A2(n900), .ZN(n694) );
  NAND2_X1 U778 ( .A1(n695), .A2(n694), .ZN(n699) );
  NAND2_X1 U779 ( .A1(G119), .A2(n570), .ZN(n697) );
  NAND2_X1 U780 ( .A1(G107), .A2(n896), .ZN(n696) );
  NAND2_X1 U781 ( .A1(n697), .A2(n696), .ZN(n698) );
  OR2_X1 U782 ( .A1(n699), .A2(n698), .ZN(n916) );
  AND2_X1 U783 ( .A1(n916), .A2(G1991), .ZN(n708) );
  NAND2_X1 U784 ( .A1(G129), .A2(n570), .ZN(n701) );
  NAND2_X1 U785 ( .A1(G141), .A2(n900), .ZN(n700) );
  NAND2_X1 U786 ( .A1(n701), .A2(n700), .ZN(n704) );
  NAND2_X1 U787 ( .A1(n566), .A2(G105), .ZN(n702) );
  XOR2_X1 U788 ( .A(KEYINPUT38), .B(n702), .Z(n703) );
  NOR2_X1 U789 ( .A1(n704), .A2(n703), .ZN(n706) );
  NAND2_X1 U790 ( .A1(n896), .A2(G117), .ZN(n705) );
  NAND2_X1 U791 ( .A1(n706), .A2(n705), .ZN(n909) );
  AND2_X1 U792 ( .A1(G1996), .A2(n909), .ZN(n707) );
  NOR2_X1 U793 ( .A1(n708), .A2(n707), .ZN(n1014) );
  NAND2_X1 U794 ( .A1(G160), .A2(G40), .ZN(n723) );
  NOR2_X1 U795 ( .A1(n724), .A2(n723), .ZN(n837) );
  INV_X1 U796 ( .A(n837), .ZN(n709) );
  NOR2_X1 U797 ( .A1(n1014), .A2(n709), .ZN(n829) );
  XOR2_X1 U798 ( .A(KEYINPUT88), .B(n829), .Z(n721) );
  NAND2_X1 U799 ( .A1(G104), .A2(n566), .ZN(n711) );
  NAND2_X1 U800 ( .A1(G140), .A2(n900), .ZN(n710) );
  NAND2_X1 U801 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U802 ( .A(KEYINPUT34), .B(n712), .ZN(n719) );
  NAND2_X1 U803 ( .A1(n570), .A2(G128), .ZN(n713) );
  XNOR2_X1 U804 ( .A(n713), .B(KEYINPUT86), .ZN(n715) );
  NAND2_X1 U805 ( .A1(G116), .A2(n896), .ZN(n714) );
  NAND2_X1 U806 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U807 ( .A(KEYINPUT87), .B(n716), .ZN(n717) );
  XNOR2_X1 U808 ( .A(KEYINPUT35), .B(n717), .ZN(n718) );
  NOR2_X1 U809 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U810 ( .A(KEYINPUT36), .B(n720), .ZN(n919) );
  XNOR2_X1 U811 ( .A(KEYINPUT37), .B(G2067), .ZN(n834) );
  NOR2_X1 U812 ( .A1(n919), .A2(n834), .ZN(n1012) );
  NAND2_X1 U813 ( .A1(n837), .A2(n1012), .ZN(n832) );
  NAND2_X1 U814 ( .A1(n721), .A2(n832), .ZN(n821) );
  NOR2_X1 U815 ( .A1(G2090), .A2(G303), .ZN(n722) );
  NAND2_X1 U816 ( .A1(G8), .A2(n722), .ZN(n799) );
  INV_X1 U817 ( .A(n723), .ZN(n725) );
  NAND2_X1 U818 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X2 U819 ( .A(n726), .B(KEYINPUT64), .ZN(n763) );
  INV_X1 U820 ( .A(n763), .ZN(n752) );
  NOR2_X1 U821 ( .A1(G1961), .A2(n752), .ZN(n727) );
  XOR2_X1 U822 ( .A(KEYINPUT90), .B(n727), .Z(n729) );
  XNOR2_X1 U823 ( .A(G2078), .B(KEYINPUT25), .ZN(n934) );
  NAND2_X1 U824 ( .A1(n752), .A2(n934), .ZN(n728) );
  NAND2_X1 U825 ( .A1(n729), .A2(n728), .ZN(n767) );
  NAND2_X1 U826 ( .A1(n767), .A2(G171), .ZN(n784) );
  INV_X1 U827 ( .A(G2067), .ZN(n730) );
  OR2_X1 U828 ( .A1(n763), .A2(n730), .ZN(n731) );
  XNOR2_X1 U829 ( .A(n731), .B(KEYINPUT92), .ZN(n733) );
  NAND2_X1 U830 ( .A1(G1348), .A2(n779), .ZN(n732) );
  NAND2_X1 U831 ( .A1(n733), .A2(n732), .ZN(n735) );
  INV_X1 U832 ( .A(KEYINPUT93), .ZN(n734) );
  XNOR2_X1 U833 ( .A(n735), .B(n734), .ZN(n743) );
  INV_X1 U834 ( .A(n988), .ZN(n736) );
  OR2_X1 U835 ( .A1(n736), .A2(n989), .ZN(n738) );
  NAND2_X1 U836 ( .A1(n779), .A2(G1341), .ZN(n745) );
  INV_X1 U837 ( .A(n745), .ZN(n737) );
  NOR2_X1 U838 ( .A1(n738), .A2(n737), .ZN(n741) );
  AND2_X1 U839 ( .A1(n752), .A2(G1996), .ZN(n740) );
  XNOR2_X1 U840 ( .A(KEYINPUT26), .B(KEYINPUT91), .ZN(n739) );
  XNOR2_X1 U841 ( .A(n740), .B(n739), .ZN(n746) );
  NAND2_X1 U842 ( .A1(n741), .A2(n746), .ZN(n742) );
  NAND2_X1 U843 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U844 ( .A(n744), .B(KEYINPUT94), .ZN(n750) );
  NAND2_X1 U845 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U846 ( .A1(n989), .A2(n747), .ZN(n748) );
  OR2_X1 U847 ( .A1(n748), .A2(n988), .ZN(n749) );
  NAND2_X1 U848 ( .A1(n750), .A2(n749), .ZN(n756) );
  NAND2_X1 U849 ( .A1(G2072), .A2(n752), .ZN(n751) );
  XNOR2_X1 U850 ( .A(n751), .B(KEYINPUT27), .ZN(n754) );
  INV_X1 U851 ( .A(G1956), .ZN(n951) );
  NOR2_X1 U852 ( .A1(n752), .A2(n951), .ZN(n753) );
  NOR2_X1 U853 ( .A1(n754), .A2(n753), .ZN(n758) );
  INV_X1 U854 ( .A(G299), .ZN(n757) );
  NAND2_X1 U855 ( .A1(n758), .A2(n757), .ZN(n755) );
  NAND2_X1 U856 ( .A1(n756), .A2(n755), .ZN(n761) );
  NOR2_X1 U857 ( .A1(n758), .A2(n757), .ZN(n759) );
  XOR2_X1 U858 ( .A(n759), .B(KEYINPUT28), .Z(n760) );
  NAND2_X1 U859 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U860 ( .A1(n784), .A2(n523), .ZN(n772) );
  NAND2_X1 U861 ( .A1(G8), .A2(n763), .ZN(n816) );
  NOR2_X1 U862 ( .A1(G1966), .A2(n816), .ZN(n775) );
  NOR2_X1 U863 ( .A1(n779), .A2(G2084), .ZN(n773) );
  NOR2_X1 U864 ( .A1(n775), .A2(n773), .ZN(n764) );
  NAND2_X1 U865 ( .A1(G8), .A2(n764), .ZN(n765) );
  XNOR2_X1 U866 ( .A(KEYINPUT30), .B(n765), .ZN(n766) );
  NOR2_X1 U867 ( .A1(G168), .A2(n766), .ZN(n769) );
  NOR2_X1 U868 ( .A1(G171), .A2(n767), .ZN(n768) );
  NOR2_X1 U869 ( .A1(n769), .A2(n768), .ZN(n771) );
  INV_X1 U870 ( .A(KEYINPUT31), .ZN(n770) );
  XNOR2_X1 U871 ( .A(n771), .B(n770), .ZN(n788) );
  NAND2_X1 U872 ( .A1(G8), .A2(n773), .ZN(n774) );
  XOR2_X1 U873 ( .A(KEYINPUT89), .B(n774), .Z(n777) );
  INV_X1 U874 ( .A(n775), .ZN(n776) );
  NOR2_X1 U875 ( .A1(G1971), .A2(n816), .ZN(n781) );
  NOR2_X1 U876 ( .A1(n779), .A2(G2090), .ZN(n780) );
  NOR2_X1 U877 ( .A1(n781), .A2(n780), .ZN(n782) );
  NAND2_X1 U878 ( .A1(n782), .A2(G303), .ZN(n787) );
  INV_X1 U879 ( .A(n787), .ZN(n783) );
  OR2_X1 U880 ( .A1(n783), .A2(G286), .ZN(n786) );
  AND2_X1 U881 ( .A1(n784), .A2(n786), .ZN(n785) );
  NAND2_X1 U882 ( .A1(n523), .A2(n785), .ZN(n792) );
  INV_X1 U883 ( .A(n786), .ZN(n790) );
  AND2_X1 U884 ( .A1(n788), .A2(n787), .ZN(n789) );
  NAND2_X1 U885 ( .A1(n792), .A2(n791), .ZN(n793) );
  NAND2_X1 U886 ( .A1(n793), .A2(G8), .ZN(n795) );
  XOR2_X1 U887 ( .A(KEYINPUT95), .B(KEYINPUT32), .Z(n794) );
  XNOR2_X1 U888 ( .A(n795), .B(n794), .ZN(n796) );
  NAND2_X1 U889 ( .A1(n797), .A2(n796), .ZN(n798) );
  XNOR2_X1 U890 ( .A(n798), .B(KEYINPUT96), .ZN(n811) );
  NAND2_X1 U891 ( .A1(n799), .A2(n811), .ZN(n800) );
  NAND2_X1 U892 ( .A1(n800), .A2(n816), .ZN(n806) );
  XNOR2_X1 U893 ( .A(KEYINPUT97), .B(G1981), .ZN(n801) );
  XNOR2_X1 U894 ( .A(n801), .B(G305), .ZN(n983) );
  NOR2_X1 U895 ( .A1(G288), .A2(G1976), .ZN(n809) );
  INV_X1 U896 ( .A(n809), .ZN(n976) );
  NOR2_X1 U897 ( .A1(n816), .A2(n976), .ZN(n802) );
  NAND2_X1 U898 ( .A1(KEYINPUT33), .A2(n802), .ZN(n803) );
  NAND2_X1 U899 ( .A1(n983), .A2(n803), .ZN(n813) );
  INV_X1 U900 ( .A(n813), .ZN(n804) );
  NAND2_X1 U901 ( .A1(KEYINPUT33), .A2(n804), .ZN(n805) );
  NAND2_X1 U902 ( .A1(n806), .A2(n805), .ZN(n819) );
  NOR2_X1 U903 ( .A1(G1981), .A2(G305), .ZN(n807) );
  XNOR2_X1 U904 ( .A(KEYINPUT24), .B(n807), .ZN(n815) );
  NOR2_X1 U905 ( .A1(G1971), .A2(G303), .ZN(n808) );
  NOR2_X1 U906 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U907 ( .A1(n811), .A2(n810), .ZN(n814) );
  NAND2_X1 U908 ( .A1(G1976), .A2(G288), .ZN(n977) );
  NOR2_X1 U909 ( .A1(n815), .A2(n526), .ZN(n817) );
  NOR2_X1 U910 ( .A1(n817), .A2(n816), .ZN(n818) );
  NOR2_X1 U911 ( .A1(n819), .A2(n818), .ZN(n820) );
  NOR2_X1 U912 ( .A1(n821), .A2(n820), .ZN(n822) );
  XNOR2_X1 U913 ( .A(n822), .B(KEYINPUT98), .ZN(n825) );
  XNOR2_X1 U914 ( .A(G1986), .B(G290), .ZN(n980) );
  NAND2_X1 U915 ( .A1(n837), .A2(n980), .ZN(n823) );
  XOR2_X1 U916 ( .A(KEYINPUT85), .B(n823), .Z(n824) );
  NAND2_X1 U917 ( .A1(n825), .A2(n824), .ZN(n840) );
  NOR2_X1 U918 ( .A1(G1996), .A2(n909), .ZN(n826) );
  XOR2_X1 U919 ( .A(KEYINPUT99), .B(n826), .Z(n1005) );
  NOR2_X1 U920 ( .A1(G1991), .A2(n916), .ZN(n1009) );
  NOR2_X1 U921 ( .A1(G1986), .A2(G290), .ZN(n827) );
  NOR2_X1 U922 ( .A1(n1009), .A2(n827), .ZN(n828) );
  NOR2_X1 U923 ( .A1(n829), .A2(n828), .ZN(n830) );
  NOR2_X1 U924 ( .A1(n1005), .A2(n830), .ZN(n831) );
  XNOR2_X1 U925 ( .A(KEYINPUT39), .B(n831), .ZN(n833) );
  NAND2_X1 U926 ( .A1(n833), .A2(n832), .ZN(n836) );
  NAND2_X1 U927 ( .A1(n919), .A2(n834), .ZN(n835) );
  XNOR2_X1 U928 ( .A(KEYINPUT100), .B(n835), .ZN(n1024) );
  NAND2_X1 U929 ( .A1(n836), .A2(n1024), .ZN(n838) );
  NAND2_X1 U930 ( .A1(n838), .A2(n837), .ZN(n839) );
  NAND2_X1 U931 ( .A1(n840), .A2(n839), .ZN(n841) );
  XNOR2_X1 U932 ( .A(n841), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U933 ( .A1(n842), .A2(G2106), .ZN(n843) );
  XNOR2_X1 U934 ( .A(n843), .B(KEYINPUT102), .ZN(G217) );
  NAND2_X1 U935 ( .A1(G15), .A2(G2), .ZN(n844) );
  XNOR2_X1 U936 ( .A(KEYINPUT103), .B(n844), .ZN(n845) );
  NAND2_X1 U937 ( .A1(n845), .A2(G661), .ZN(G259) );
  NAND2_X1 U938 ( .A1(G3), .A2(G1), .ZN(n846) );
  XNOR2_X1 U939 ( .A(KEYINPUT104), .B(n846), .ZN(n848) );
  NAND2_X1 U940 ( .A1(n848), .A2(n847), .ZN(G188) );
  NOR2_X1 U941 ( .A1(n850), .A2(n849), .ZN(G325) );
  XNOR2_X1 U942 ( .A(KEYINPUT105), .B(G325), .ZN(G261) );
  XNOR2_X1 U944 ( .A(KEYINPUT77), .B(n851), .ZN(n852) );
  NOR2_X1 U945 ( .A1(G860), .A2(n852), .ZN(n854) );
  XOR2_X1 U946 ( .A(n854), .B(n853), .Z(G145) );
  INV_X1 U947 ( .A(G120), .ZN(G236) );
  INV_X1 U948 ( .A(G96), .ZN(G221) );
  INV_X1 U949 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U950 ( .A(G171), .B(n989), .ZN(n855) );
  XNOR2_X1 U951 ( .A(n855), .B(G286), .ZN(n858) );
  XOR2_X1 U952 ( .A(n736), .B(n856), .Z(n857) );
  XNOR2_X1 U953 ( .A(n858), .B(n857), .ZN(n859) );
  NOR2_X1 U954 ( .A1(G37), .A2(n859), .ZN(G397) );
  XOR2_X1 U955 ( .A(G2474), .B(G1976), .Z(n861) );
  XNOR2_X1 U956 ( .A(G1986), .B(G1956), .ZN(n860) );
  XNOR2_X1 U957 ( .A(n861), .B(n860), .ZN(n862) );
  XOR2_X1 U958 ( .A(n862), .B(KEYINPUT106), .Z(n864) );
  XNOR2_X1 U959 ( .A(G1996), .B(G1991), .ZN(n863) );
  XNOR2_X1 U960 ( .A(n864), .B(n863), .ZN(n868) );
  XOR2_X1 U961 ( .A(G1981), .B(G1971), .Z(n866) );
  XNOR2_X1 U962 ( .A(G1966), .B(G1961), .ZN(n865) );
  XNOR2_X1 U963 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U964 ( .A(n868), .B(n867), .Z(n870) );
  XNOR2_X1 U965 ( .A(KEYINPUT107), .B(KEYINPUT41), .ZN(n869) );
  XNOR2_X1 U966 ( .A(n870), .B(n869), .ZN(G229) );
  XOR2_X1 U967 ( .A(G2100), .B(G2096), .Z(n872) );
  XNOR2_X1 U968 ( .A(KEYINPUT42), .B(G2678), .ZN(n871) );
  XNOR2_X1 U969 ( .A(n872), .B(n871), .ZN(n876) );
  XOR2_X1 U970 ( .A(KEYINPUT43), .B(G2072), .Z(n874) );
  XNOR2_X1 U971 ( .A(G2067), .B(G2090), .ZN(n873) );
  XNOR2_X1 U972 ( .A(n874), .B(n873), .ZN(n875) );
  XOR2_X1 U973 ( .A(n876), .B(n875), .Z(n878) );
  XNOR2_X1 U974 ( .A(G2078), .B(G2084), .ZN(n877) );
  XNOR2_X1 U975 ( .A(n878), .B(n877), .ZN(G227) );
  XOR2_X1 U976 ( .A(KEYINPUT44), .B(KEYINPUT109), .Z(n880) );
  NAND2_X1 U977 ( .A1(G124), .A2(n570), .ZN(n879) );
  XNOR2_X1 U978 ( .A(n880), .B(n879), .ZN(n881) );
  XNOR2_X1 U979 ( .A(n881), .B(KEYINPUT108), .ZN(n883) );
  NAND2_X1 U980 ( .A1(n566), .A2(G100), .ZN(n882) );
  NAND2_X1 U981 ( .A1(n883), .A2(n882), .ZN(n887) );
  NAND2_X1 U982 ( .A1(G136), .A2(n900), .ZN(n885) );
  NAND2_X1 U983 ( .A1(G112), .A2(n896), .ZN(n884) );
  NAND2_X1 U984 ( .A1(n885), .A2(n884), .ZN(n886) );
  NOR2_X1 U985 ( .A1(n887), .A2(n886), .ZN(G162) );
  NAND2_X1 U986 ( .A1(G103), .A2(n899), .ZN(n889) );
  NAND2_X1 U987 ( .A1(G139), .A2(n900), .ZN(n888) );
  NAND2_X1 U988 ( .A1(n889), .A2(n888), .ZN(n895) );
  NAND2_X1 U989 ( .A1(G127), .A2(n570), .ZN(n891) );
  NAND2_X1 U990 ( .A1(G115), .A2(n896), .ZN(n890) );
  NAND2_X1 U991 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U992 ( .A(KEYINPUT47), .B(n892), .Z(n893) );
  XNOR2_X1 U993 ( .A(KEYINPUT110), .B(n893), .ZN(n894) );
  NOR2_X1 U994 ( .A1(n895), .A2(n894), .ZN(n1020) );
  XNOR2_X1 U995 ( .A(G160), .B(n1008), .ZN(n907) );
  NAND2_X1 U996 ( .A1(G130), .A2(n570), .ZN(n898) );
  NAND2_X1 U997 ( .A1(G118), .A2(n896), .ZN(n897) );
  NAND2_X1 U998 ( .A1(n898), .A2(n897), .ZN(n905) );
  NAND2_X1 U999 ( .A1(G106), .A2(n899), .ZN(n902) );
  NAND2_X1 U1000 ( .A1(G142), .A2(n900), .ZN(n901) );
  NAND2_X1 U1001 ( .A1(n902), .A2(n901), .ZN(n903) );
  XOR2_X1 U1002 ( .A(KEYINPUT45), .B(n903), .Z(n904) );
  NOR2_X1 U1003 ( .A1(n905), .A2(n904), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(n1020), .B(n908), .ZN(n911) );
  XOR2_X1 U1006 ( .A(G164), .B(n909), .Z(n910) );
  XNOR2_X1 U1007 ( .A(n911), .B(n910), .ZN(n915) );
  XOR2_X1 U1008 ( .A(KEYINPUT112), .B(KEYINPUT46), .Z(n913) );
  XNOR2_X1 U1009 ( .A(KEYINPUT111), .B(KEYINPUT48), .ZN(n912) );
  XNOR2_X1 U1010 ( .A(n913), .B(n912), .ZN(n914) );
  XOR2_X1 U1011 ( .A(n915), .B(n914), .Z(n918) );
  XOR2_X1 U1012 ( .A(n916), .B(G162), .Z(n917) );
  XNOR2_X1 U1013 ( .A(n918), .B(n917), .ZN(n920) );
  XOR2_X1 U1014 ( .A(n920), .B(n919), .Z(n921) );
  NOR2_X1 U1015 ( .A1(G37), .A2(n921), .ZN(G395) );
  NOR2_X1 U1016 ( .A1(G401), .A2(n928), .ZN(n925) );
  NOR2_X1 U1017 ( .A1(G229), .A2(G227), .ZN(n922) );
  XNOR2_X1 U1018 ( .A(KEYINPUT49), .B(n922), .ZN(n923) );
  NOR2_X1 U1019 ( .A1(G397), .A2(n923), .ZN(n924) );
  NAND2_X1 U1020 ( .A1(n925), .A2(n924), .ZN(n926) );
  NOR2_X1 U1021 ( .A1(n926), .A2(G395), .ZN(n927) );
  XNOR2_X1 U1022 ( .A(n927), .B(KEYINPUT113), .ZN(G225) );
  XOR2_X1 U1023 ( .A(KEYINPUT114), .B(G225), .Z(G308) );
  INV_X1 U1024 ( .A(n928), .ZN(G319) );
  INV_X1 U1025 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1026 ( .A(KEYINPUT119), .B(G34), .Z(n930) );
  XNOR2_X1 U1027 ( .A(G2084), .B(KEYINPUT54), .ZN(n929) );
  XNOR2_X1 U1028 ( .A(n930), .B(n929), .ZN(n946) );
  XOR2_X1 U1029 ( .A(G2090), .B(G35), .Z(n944) );
  XOR2_X1 U1030 ( .A(G2067), .B(G26), .Z(n931) );
  NAND2_X1 U1031 ( .A1(n931), .A2(G28), .ZN(n940) );
  XNOR2_X1 U1032 ( .A(G1996), .B(G32), .ZN(n933) );
  XNOR2_X1 U1033 ( .A(G33), .B(G2072), .ZN(n932) );
  NOR2_X1 U1034 ( .A1(n933), .A2(n932), .ZN(n938) );
  XOR2_X1 U1035 ( .A(n934), .B(G27), .Z(n936) );
  XNOR2_X1 U1036 ( .A(G1991), .B(G25), .ZN(n935) );
  NOR2_X1 U1037 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1038 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1040 ( .A(KEYINPUT118), .B(n941), .Z(n942) );
  XNOR2_X1 U1041 ( .A(n942), .B(KEYINPUT53), .ZN(n943) );
  NAND2_X1 U1042 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1043 ( .A1(n946), .A2(n945), .ZN(n947) );
  XOR2_X1 U1044 ( .A(KEYINPUT55), .B(n947), .Z(n948) );
  NOR2_X1 U1045 ( .A1(G29), .A2(n948), .ZN(n949) );
  XOR2_X1 U1046 ( .A(KEYINPUT120), .B(n949), .Z(n950) );
  NAND2_X1 U1047 ( .A1(G11), .A2(n950), .ZN(n1035) );
  XOR2_X1 U1048 ( .A(G1961), .B(G5), .Z(n961) );
  XNOR2_X1 U1049 ( .A(G20), .B(n951), .ZN(n955) );
  XNOR2_X1 U1050 ( .A(G1341), .B(G19), .ZN(n953) );
  XNOR2_X1 U1051 ( .A(G6), .B(G1981), .ZN(n952) );
  NOR2_X1 U1052 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1053 ( .A1(n955), .A2(n954), .ZN(n958) );
  XOR2_X1 U1054 ( .A(KEYINPUT59), .B(G1348), .Z(n956) );
  XNOR2_X1 U1055 ( .A(G4), .B(n956), .ZN(n957) );
  NOR2_X1 U1056 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1057 ( .A(KEYINPUT60), .B(n959), .ZN(n960) );
  NAND2_X1 U1058 ( .A1(n961), .A2(n960), .ZN(n963) );
  XNOR2_X1 U1059 ( .A(G21), .B(G1966), .ZN(n962) );
  NOR2_X1 U1060 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1061 ( .A(KEYINPUT124), .B(n964), .ZN(n972) );
  XOR2_X1 U1062 ( .A(G1986), .B(G24), .Z(n965) );
  XNOR2_X1 U1063 ( .A(KEYINPUT125), .B(n965), .ZN(n969) );
  XOR2_X1 U1064 ( .A(G1971), .B(G22), .Z(n967) );
  XOR2_X1 U1065 ( .A(G1976), .B(G23), .Z(n966) );
  NAND2_X1 U1066 ( .A1(n967), .A2(n966), .ZN(n968) );
  NOR2_X1 U1067 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1068 ( .A(KEYINPUT58), .B(n970), .ZN(n971) );
  NAND2_X1 U1069 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1070 ( .A(n973), .B(KEYINPUT126), .ZN(n974) );
  XNOR2_X1 U1071 ( .A(KEYINPUT61), .B(n974), .ZN(n975) );
  NOR2_X1 U1072 ( .A1(G16), .A2(n975), .ZN(n1003) );
  XNOR2_X1 U1073 ( .A(G16), .B(KEYINPUT56), .ZN(n1000) );
  XNOR2_X1 U1074 ( .A(G166), .B(G1971), .ZN(n982) );
  NAND2_X1 U1075 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1076 ( .A(KEYINPUT122), .B(n978), .ZN(n979) );
  NOR2_X1 U1077 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1078 ( .A1(n982), .A2(n981), .ZN(n987) );
  XNOR2_X1 U1079 ( .A(G1966), .B(G168), .ZN(n984) );
  NAND2_X1 U1080 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1081 ( .A(KEYINPUT57), .B(n985), .Z(n986) );
  NOR2_X1 U1082 ( .A1(n987), .A2(n986), .ZN(n998) );
  XNOR2_X1 U1083 ( .A(n988), .B(G1348), .ZN(n993) );
  XNOR2_X1 U1084 ( .A(G301), .B(G1961), .ZN(n991) );
  XNOR2_X1 U1085 ( .A(n989), .B(G1341), .ZN(n990) );
  NOR2_X1 U1086 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1087 ( .A1(n993), .A2(n992), .ZN(n996) );
  XOR2_X1 U1088 ( .A(G1956), .B(G299), .Z(n994) );
  XNOR2_X1 U1089 ( .A(KEYINPUT121), .B(n994), .ZN(n995) );
  NOR2_X1 U1090 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1091 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1093 ( .A(KEYINPUT123), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1033) );
  XOR2_X1 U1095 ( .A(G2090), .B(G162), .Z(n1004) );
  NOR2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1097 ( .A(KEYINPUT117), .B(n1006), .Z(n1007) );
  XOR2_X1 U1098 ( .A(KEYINPUT51), .B(n1007), .Z(n1019) );
  NOR2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1100 ( .A(KEYINPUT115), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1016) );
  XOR2_X1 U1103 ( .A(G160), .B(G2084), .Z(n1015) );
  NOR2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1105 ( .A(KEYINPUT116), .B(n1017), .ZN(n1018) );
  NAND2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1027) );
  XOR2_X1 U1107 ( .A(G2072), .B(n1020), .Z(n1022) );
  XOR2_X1 U1108 ( .A(G164), .B(G2078), .Z(n1021) );
  NOR2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1110 ( .A(KEYINPUT50), .B(n1023), .ZN(n1025) );
  NAND2_X1 U1111 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NOR2_X1 U1112 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1113 ( .A(KEYINPUT52), .B(n1028), .ZN(n1030) );
  INV_X1 U1114 ( .A(KEYINPUT55), .ZN(n1029) );
  NAND2_X1 U1115 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1116 ( .A1(n1031), .A2(G29), .ZN(n1032) );
  NAND2_X1 U1117 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NOR2_X1 U1118 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XOR2_X1 U1119 ( .A(KEYINPUT127), .B(n1036), .Z(n1037) );
  XNOR2_X1 U1120 ( .A(KEYINPUT62), .B(n1037), .ZN(G311) );
  INV_X1 U1121 ( .A(G311), .ZN(G150) );
endmodule

