//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 1 0 1 0 1 1 0 0 1 0 0 1 1 0 1 0 0 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n759, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n851, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941;
  XOR2_X1   g000(.A(G15gat), .B(G22gat), .Z(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT96), .ZN(new_n203));
  INV_X1    g002(.A(G1gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  AOI21_X1  g004(.A(G8gat), .B1(new_n205), .B2(KEYINPUT97), .ZN(new_n206));
  AND2_X1   g005(.A1(new_n204), .A2(KEYINPUT16), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n205), .B1(new_n203), .B2(new_n207), .ZN(new_n208));
  OR2_X1    g007(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n206), .A2(new_n208), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT14), .ZN(new_n211));
  OR3_X1    g010(.A1(new_n211), .A2(G29gat), .A3(G36gat), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n211), .B1(G29gat), .B2(G36gat), .ZN(new_n213));
  XNOR2_X1  g012(.A(KEYINPUT95), .B(G36gat), .ZN(new_n214));
  INV_X1    g013(.A(G29gat), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n212), .B(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G43gat), .B(G50gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n217), .A2(KEYINPUT15), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT15), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n220), .B1(new_n217), .B2(KEYINPUT94), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(KEYINPUT94), .B2(new_n217), .ZN(new_n222));
  MUX2_X1   g021(.A(new_n216), .B(new_n219), .S(new_n222), .Z(new_n223));
  AND3_X1   g022(.A1(new_n209), .A2(new_n210), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n209), .A2(new_n210), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n223), .B(KEYINPUT17), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G229gat), .A2(G233gat), .ZN(new_n228));
  AND2_X1   g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OR2_X1    g028(.A1(new_n229), .A2(KEYINPUT18), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n227), .A2(KEYINPUT18), .A3(new_n228), .ZN(new_n231));
  XOR2_X1   g030(.A(new_n225), .B(new_n223), .Z(new_n232));
  XOR2_X1   g031(.A(new_n228), .B(KEYINPUT13), .Z(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n230), .A2(new_n231), .A3(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(G113gat), .B(G141gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(KEYINPUT93), .B(G197gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g037(.A(KEYINPUT11), .B(G169gat), .Z(new_n239));
  XNOR2_X1  g038(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g039(.A(new_n240), .B(KEYINPUT12), .Z(new_n241));
  OR2_X1    g040(.A1(new_n235), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n235), .A2(new_n241), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(G226gat), .A2(G233gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(KEYINPUT27), .B(G183gat), .ZN(new_n247));
  INV_X1    g046(.A(G190gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(KEYINPUT28), .ZN(new_n250));
  INV_X1    g049(.A(G169gat), .ZN(new_n251));
  INV_X1    g050(.A(G176gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT26), .ZN(new_n254));
  NAND2_X1  g053(.A1(G169gat), .A2(G176gat), .ZN(new_n255));
  AND3_X1   g054(.A1(new_n253), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(G183gat), .A2(G190gat), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n257), .B1(new_n253), .B2(new_n254), .ZN(new_n258));
  NOR3_X1   g057(.A1(new_n250), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT64), .ZN(new_n260));
  NAND3_X1  g059(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n261), .B1(G183gat), .B2(G190gat), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n260), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n263), .ZN(new_n265));
  OR2_X1    g064(.A1(G183gat), .A2(G190gat), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n265), .A2(new_n266), .A3(KEYINPUT64), .A4(new_n261), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n251), .A2(new_n252), .A3(KEYINPUT23), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT23), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n269), .B1(G169gat), .B2(G176gat), .ZN(new_n270));
  AND3_X1   g069(.A1(new_n268), .A2(new_n270), .A3(new_n255), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n264), .A2(new_n267), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT25), .ZN(new_n273));
  AOI21_X1  g072(.A(KEYINPUT65), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT66), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n257), .B1(new_n275), .B2(KEYINPUT24), .ZN(new_n276));
  AND2_X1   g075(.A1(new_n275), .A2(KEYINPUT24), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n266), .B(new_n261), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n278), .A2(new_n271), .A3(KEYINPUT25), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n274), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n272), .A2(KEYINPUT65), .A3(new_n273), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n259), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n246), .B1(new_n283), .B2(KEYINPUT29), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT73), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G197gat), .B(G204gat), .ZN(new_n287));
  INV_X1    g086(.A(G211gat), .ZN(new_n288));
  INV_X1    g087(.A(G218gat), .ZN(new_n289));
  OAI22_X1  g088(.A1(new_n288), .A2(new_n289), .B1(KEYINPUT71), .B2(KEYINPUT22), .ZN(new_n290));
  AND2_X1   g089(.A1(KEYINPUT71), .A2(KEYINPUT22), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n287), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n292), .B(KEYINPUT72), .ZN(new_n293));
  XOR2_X1   g092(.A(G211gat), .B(G218gat), .Z(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  OR2_X1    g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n293), .A2(new_n295), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n272), .A2(new_n273), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT65), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n301), .A2(new_n282), .A3(new_n279), .ZN(new_n302));
  OR3_X1    g101(.A1(new_n250), .A2(new_n256), .A3(new_n258), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n246), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT29), .ZN(new_n305));
  INV_X1    g104(.A(new_n282), .ZN(new_n306));
  NOR3_X1   g105(.A1(new_n306), .A2(new_n274), .A3(new_n280), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n305), .B1(new_n307), .B2(new_n259), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n304), .B1(new_n308), .B2(new_n246), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n286), .B(new_n298), .C1(new_n309), .C2(new_n285), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n284), .B1(new_n283), .B2(new_n246), .ZN(new_n311));
  INV_X1    g110(.A(new_n298), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  XOR2_X1   g112(.A(G8gat), .B(G36gat), .Z(new_n314));
  XNOR2_X1  g113(.A(G64gat), .B(G92gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n314), .B(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n317));
  XOR2_X1   g116(.A(new_n316), .B(new_n317), .Z(new_n318));
  NAND3_X1  g117(.A1(new_n310), .A2(new_n313), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT30), .ZN(new_n320));
  OR2_X1    g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n310), .A2(new_n313), .ZN(new_n322));
  INV_X1    g121(.A(new_n318), .ZN(new_n323));
  AOI21_X1  g122(.A(KEYINPUT76), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT76), .ZN(new_n325));
  AOI211_X1 g124(.A(new_n325), .B(new_n318), .C1(new_n310), .C2(new_n313), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n321), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT77), .ZN(new_n328));
  AND3_X1   g127(.A1(new_n319), .A2(new_n328), .A3(new_n320), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n328), .B1(new_n319), .B2(new_n320), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT35), .ZN(new_n333));
  XNOR2_X1  g132(.A(G127gat), .B(G134gat), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT67), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n334), .B(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(G113gat), .ZN(new_n337));
  INV_X1    g136(.A(G120gat), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT1), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n339), .B1(new_n337), .B2(new_n338), .ZN(new_n340));
  AND2_X1   g139(.A1(new_n334), .A2(new_n339), .ZN(new_n341));
  XNOR2_X1  g140(.A(KEYINPUT68), .B(G113gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(G120gat), .ZN(new_n343));
  AOI22_X1  g142(.A1(new_n336), .A2(new_n340), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  NOR2_X1   g143(.A1(G155gat), .A2(G162gat), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G155gat), .A2(G162gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  XOR2_X1   g147(.A(G141gat), .B(G148gat), .Z(new_n349));
  INV_X1    g148(.A(KEYINPUT2), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n348), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT79), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n345), .A2(new_n350), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT78), .ZN(new_n355));
  INV_X1    g154(.A(G141gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(KEYINPUT78), .A2(G141gat), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n357), .A2(G148gat), .A3(new_n358), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n356), .A2(G148gat), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  AOI221_X4 g160(.A(new_n353), .B1(new_n354), .B2(new_n347), .C1(new_n359), .C2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n359), .A2(new_n361), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n354), .A2(new_n347), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT79), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n352), .B1(new_n362), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n344), .B1(new_n366), .B2(KEYINPUT3), .ZN(new_n367));
  NOR3_X1   g166(.A1(new_n366), .A2(KEYINPUT80), .A3(KEYINPUT3), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT80), .ZN(new_n369));
  AND2_X1   g168(.A1(KEYINPUT78), .A2(G141gat), .ZN(new_n370));
  NOR2_X1   g169(.A1(KEYINPUT78), .A2(G141gat), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n360), .B1(new_n372), .B2(G148gat), .ZN(new_n373));
  AND2_X1   g172(.A1(new_n354), .A2(new_n347), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n353), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n363), .A2(KEYINPUT79), .A3(new_n364), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n351), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT3), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n369), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n367), .B1(new_n368), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT5), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n341), .A2(new_n343), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n334), .B(KEYINPUT67), .ZN(new_n383));
  INV_X1    g182(.A(new_n340), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n382), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT4), .ZN(new_n386));
  NOR3_X1   g185(.A1(new_n366), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT4), .B1(new_n377), .B2(new_n344), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(G225gat), .A2(G233gat), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n380), .A2(new_n381), .A3(new_n389), .A4(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n385), .B1(new_n377), .B2(new_n378), .ZN(new_n392));
  OAI21_X1  g191(.A(KEYINPUT80), .B1(new_n366), .B2(KEYINPUT3), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n377), .A2(new_n369), .A3(new_n378), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n390), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n386), .B1(new_n366), .B2(new_n385), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n377), .A2(KEYINPUT4), .A3(new_n344), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NOR3_X1   g198(.A1(new_n395), .A2(new_n396), .A3(new_n399), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n366), .A2(new_n385), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n377), .A2(new_n344), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n396), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT5), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n391), .B1(new_n400), .B2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(G1gat), .B(G29gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n406), .B(KEYINPUT0), .ZN(new_n407));
  XNOR2_X1  g206(.A(G57gat), .B(G85gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n407), .B(new_n408), .ZN(new_n409));
  AND4_X1   g208(.A1(KEYINPUT81), .A2(new_n405), .A3(KEYINPUT6), .A4(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n409), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n380), .A2(new_n390), .A3(new_n389), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n377), .B(new_n344), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n381), .B1(new_n413), .B2(new_n396), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n411), .B1(new_n415), .B2(new_n391), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT81), .B1(new_n416), .B2(KEYINPUT6), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n410), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT88), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n409), .B(KEYINPUT85), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT6), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n415), .A2(new_n411), .A3(new_n391), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(KEYINPUT88), .B1(new_n410), .B2(new_n417), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n420), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n332), .A2(new_n333), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT32), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT69), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n302), .A2(new_n303), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n430), .B1(new_n431), .B2(new_n385), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n283), .A2(KEYINPUT69), .A3(new_n344), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n431), .A2(new_n385), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(G227gat), .A2(G233gat), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n429), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT33), .B1(new_n435), .B2(new_n437), .ZN(new_n439));
  XOR2_X1   g238(.A(G15gat), .B(G43gat), .Z(new_n440));
  XNOR2_X1  g239(.A(G71gat), .B(G99gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n440), .B(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  NOR3_X1   g242(.A1(new_n438), .A2(new_n439), .A3(new_n443), .ZN(new_n444));
  AOI221_X4 g243(.A(new_n429), .B1(KEYINPUT33), .B2(new_n442), .C1(new_n435), .C2(new_n437), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n432), .A2(new_n433), .A3(new_n436), .A4(new_n434), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT34), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n447), .A2(KEYINPUT34), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n446), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n435), .A2(new_n437), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT33), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n443), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n438), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n445), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n457), .A2(new_n458), .A3(new_n451), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n452), .A2(new_n460), .ZN(new_n461));
  XNOR2_X1  g260(.A(G78gat), .B(G106gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n462), .B(G50gat), .ZN(new_n463));
  XNOR2_X1  g262(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n463), .B(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n465), .B(KEYINPUT84), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT29), .B1(new_n296), .B2(new_n297), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n366), .B1(new_n468), .B2(KEYINPUT3), .ZN(new_n469));
  AOI21_X1  g268(.A(KEYINPUT29), .B1(new_n393), .B2(new_n394), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n469), .B1(new_n470), .B2(new_n298), .ZN(new_n471));
  NAND2_X1  g270(.A1(G228gat), .A2(G233gat), .ZN(new_n472));
  XOR2_X1   g271(.A(new_n472), .B(G22gat), .Z(new_n473));
  NAND2_X1  g272(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n473), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n469), .B(new_n475), .C1(new_n470), .C2(new_n298), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n467), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT84), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n465), .A2(new_n478), .ZN(new_n479));
  AND2_X1   g278(.A1(new_n474), .A2(new_n476), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n461), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n428), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n393), .A2(new_n394), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n399), .B1(new_n485), .B2(new_n367), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n404), .B1(new_n486), .B2(new_n390), .ZN(new_n487));
  INV_X1    g286(.A(new_n391), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n409), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n489), .A2(new_n423), .A3(new_n424), .ZN(new_n490));
  OAI211_X1 g289(.A(KEYINPUT6), .B(new_n409), .C1(new_n487), .C2(new_n488), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT81), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n416), .A2(KEYINPUT81), .A3(KEYINPUT6), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n490), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n495), .B(new_n321), .C1(new_n324), .C2(new_n326), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT82), .B1(new_n496), .B2(new_n331), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n319), .A2(new_n320), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n498), .B1(new_n418), .B2(new_n490), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT82), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n319), .A2(new_n320), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT77), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n319), .A2(new_n328), .A3(new_n320), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n322), .A2(new_n323), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(new_n325), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n322), .A2(KEYINPUT76), .A3(new_n323), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n499), .A2(new_n500), .A3(new_n504), .A4(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT70), .B1(new_n449), .B2(new_n450), .ZN(new_n510));
  OR2_X1    g309(.A1(new_n447), .A2(KEYINPUT34), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT70), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n511), .A2(new_n512), .A3(new_n448), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n510), .B(new_n513), .C1(new_n444), .C2(new_n445), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n514), .A2(new_n459), .A3(new_n481), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT91), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n514), .A2(KEYINPUT91), .A3(new_n459), .A4(new_n481), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n497), .A2(new_n509), .A3(new_n517), .A4(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT92), .ZN(new_n520));
  AND3_X1   g319(.A1(new_n519), .A2(new_n520), .A3(KEYINPUT35), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n520), .B1(new_n519), .B2(KEYINPUT35), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n484), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT90), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n498), .B1(new_n506), .B2(new_n507), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(new_n504), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n396), .B1(new_n395), .B2(new_n399), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n527), .A2(KEYINPUT39), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n527), .B(KEYINPUT39), .C1(new_n396), .C2(new_n413), .ZN(new_n529));
  INV_X1    g328(.A(new_n421), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT40), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n528), .A2(new_n529), .A3(KEYINPUT40), .A4(new_n530), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n533), .A2(new_n422), .A3(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT86), .B1(new_n526), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT86), .ZN(new_n538));
  AOI211_X1 g337(.A(new_n538), .B(new_n535), .C1(new_n525), .C2(new_n504), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT37), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n541), .B1(new_n311), .B2(new_n298), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n286), .B(new_n312), .C1(new_n309), .C2(new_n285), .ZN(new_n543));
  AOI21_X1  g342(.A(KEYINPUT38), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(KEYINPUT37), .B1(new_n311), .B2(new_n312), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n318), .B1(new_n545), .B2(new_n310), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT87), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT87), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n544), .A2(new_n546), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n545), .A2(new_n310), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(new_n323), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n541), .B1(new_n310), .B2(new_n313), .ZN(new_n554));
  OAI21_X1  g353(.A(KEYINPUT38), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n551), .B1(KEYINPUT89), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(KEYINPUT89), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n425), .A2(new_n319), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n557), .A2(new_n559), .A3(new_n426), .A4(new_n420), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n481), .B1(new_n556), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n524), .B1(new_n540), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n481), .ZN(new_n563));
  INV_X1    g362(.A(new_n560), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n555), .A2(KEYINPUT89), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n565), .B1(new_n548), .B2(new_n550), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n563), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n538), .B1(new_n332), .B2(new_n535), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n526), .A2(KEYINPUT86), .A3(new_n536), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n567), .A2(new_n570), .A3(KEYINPUT90), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n481), .B1(new_n497), .B2(new_n509), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT36), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n573), .B1(new_n452), .B2(new_n460), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n514), .A2(KEYINPUT36), .A3(new_n459), .ZN(new_n575));
  AND2_X1   g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n562), .A2(new_n571), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n245), .B1(new_n523), .B2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n495), .ZN(new_n580));
  XOR2_X1   g379(.A(G57gat), .B(G64gat), .Z(new_n581));
  INV_X1    g380(.A(KEYINPUT9), .ZN(new_n582));
  INV_X1    g381(.A(G71gat), .ZN(new_n583));
  INV_X1    g382(.A(G78gat), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  XOR2_X1   g385(.A(G71gat), .B(G78gat), .Z(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT21), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(G231gat), .A2(G233gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(G127gat), .B(G155gat), .Z(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  XOR2_X1   g395(.A(G183gat), .B(G211gat), .Z(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n225), .B1(new_n589), .B2(new_n588), .ZN(new_n599));
  XOR2_X1   g398(.A(KEYINPUT98), .B(KEYINPUT99), .Z(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  AND2_X1   g400(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n598), .A2(new_n601), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT8), .ZN(new_n605));
  NAND2_X1  g404(.A1(G99gat), .A2(G106gat), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n605), .B1(new_n606), .B2(KEYINPUT101), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n607), .B1(KEYINPUT101), .B2(new_n606), .ZN(new_n608));
  AND3_X1   g407(.A1(KEYINPUT100), .A2(G85gat), .A3(G92gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(KEYINPUT7), .ZN(new_n610));
  AND2_X1   g409(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT7), .ZN(new_n612));
  XOR2_X1   g411(.A(KEYINPUT102), .B(G85gat), .Z(new_n613));
  INV_X1    g412(.A(G92gat), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n612), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n611), .B1(new_n609), .B2(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(G99gat), .B(G106gat), .Z(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n617), .ZN(new_n619));
  OAI211_X1 g418(.A(new_n611), .B(new_n619), .C1(new_n609), .C2(new_n615), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  AND2_X1   g421(.A1(G232gat), .A2(G233gat), .ZN(new_n623));
  AOI22_X1  g422(.A1(new_n622), .A2(new_n223), .B1(KEYINPUT41), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT103), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n226), .B1(new_n625), .B2(new_n622), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n621), .A2(KEYINPUT103), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n624), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(G134gat), .B(G162gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XOR2_X1   g429(.A(G190gat), .B(G218gat), .Z(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(KEYINPUT104), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n623), .A2(KEYINPUT41), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  OR2_X1    g434(.A1(new_n630), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n630), .A2(new_n635), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT105), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n588), .B1(new_n620), .B2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n621), .B(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT10), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  OR3_X1    g443(.A1(new_n621), .A2(new_n643), .A3(new_n588), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(G230gat), .ZN(new_n647));
  INV_X1    g446(.A(G233gat), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n651), .B1(new_n650), .B2(new_n642), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT106), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(G120gat), .B(G148gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(G176gat), .B(G204gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  AND2_X1   g456(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n654), .A2(new_n657), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n604), .A2(new_n639), .A3(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n579), .A2(new_n580), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(G1gat), .ZN(G1324gat));
  NAND3_X1  g464(.A1(new_n579), .A2(new_n526), .A3(new_n663), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT16), .B(G8gat), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n668), .B(KEYINPUT42), .Z(new_n669));
  NAND2_X1  g468(.A1(new_n666), .A2(G8gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT107), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(KEYINPUT108), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT108), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n669), .A2(new_n674), .A3(new_n671), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n673), .A2(new_n675), .ZN(G1325gat));
  AND2_X1   g475(.A1(new_n579), .A2(new_n663), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n576), .ZN(new_n679));
  OAI21_X1  g478(.A(G15gat), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n662), .A2(G15gat), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n579), .A2(new_n461), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n680), .A2(new_n682), .ZN(G1326gat));
  NAND2_X1  g482(.A1(new_n677), .A2(new_n563), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT109), .ZN(new_n685));
  XNOR2_X1  g484(.A(KEYINPUT43), .B(G22gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(G1327gat));
  INV_X1    g486(.A(new_n604), .ZN(new_n688));
  AND4_X1   g487(.A1(new_n579), .A2(new_n688), .A3(new_n638), .A4(new_n661), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n689), .A2(new_n215), .A3(new_n580), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT110), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT45), .ZN(new_n692));
  OR2_X1    g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n245), .A2(new_n604), .A3(new_n660), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT111), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT114), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT112), .ZN(new_n698));
  AND3_X1   g497(.A1(new_n523), .A2(new_n578), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n698), .B1(new_n523), .B2(new_n578), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n638), .B(KEYINPUT113), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n702), .A2(KEYINPUT44), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n697), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  AND3_X1   g503(.A1(new_n562), .A2(new_n571), .A3(new_n577), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n519), .A2(KEYINPUT35), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(KEYINPUT92), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n519), .A2(new_n520), .A3(KEYINPUT35), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n483), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(KEYINPUT112), .B1(new_n705), .B2(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n523), .A2(new_n578), .A3(new_n698), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n710), .A2(new_n697), .A3(new_n711), .A4(new_n703), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n638), .B1(new_n705), .B2(new_n709), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(KEYINPUT44), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n696), .B1(new_n704), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(G29gat), .B1(new_n716), .B2(new_n495), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n693), .A2(new_n694), .A3(new_n717), .ZN(G1328gat));
  NAND3_X1  g517(.A1(new_n689), .A2(new_n214), .A3(new_n526), .ZN(new_n719));
  AND2_X1   g518(.A1(KEYINPUT115), .A2(KEYINPUT46), .ZN(new_n720));
  OR2_X1    g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(KEYINPUT115), .A2(KEYINPUT46), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n719), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  OR2_X1    g522(.A1(new_n716), .A2(new_n332), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  OAI211_X1 g524(.A(new_n721), .B(new_n723), .C1(new_n725), .C2(new_n214), .ZN(G1329gat));
  OAI211_X1 g525(.A(new_n576), .B(new_n696), .C1(new_n704), .C2(new_n715), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(G43gat), .ZN(new_n728));
  INV_X1    g527(.A(G43gat), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n689), .A2(new_n729), .A3(new_n461), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT47), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n728), .A2(KEYINPUT47), .A3(new_n730), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(G1330gat));
  OAI211_X1 g534(.A(new_n563), .B(new_n696), .C1(new_n704), .C2(new_n715), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(G50gat), .ZN(new_n737));
  INV_X1    g536(.A(G50gat), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n689), .A2(new_n738), .A3(new_n563), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT48), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n737), .A2(KEYINPUT48), .A3(new_n739), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(G1331gat));
  NAND4_X1  g543(.A1(new_n245), .A2(new_n604), .A3(new_n639), .A4(new_n660), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n699), .A2(new_n700), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n580), .ZN(new_n747));
  XOR2_X1   g546(.A(KEYINPUT116), .B(G57gat), .Z(new_n748));
  XNOR2_X1  g547(.A(new_n747), .B(new_n748), .ZN(G1332gat));
  NAND2_X1  g548(.A1(new_n746), .A2(new_n526), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n750), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n751));
  XOR2_X1   g550(.A(KEYINPUT49), .B(G64gat), .Z(new_n752));
  OAI21_X1  g551(.A(new_n751), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  XOR2_X1   g552(.A(new_n753), .B(KEYINPUT117), .Z(G1333gat));
  NAND3_X1  g553(.A1(new_n746), .A2(new_n583), .A3(new_n461), .ZN(new_n755));
  AND2_X1   g554(.A1(new_n746), .A2(new_n576), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n755), .B1(new_n583), .B2(new_n756), .ZN(new_n757));
  XOR2_X1   g556(.A(new_n757), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g557(.A1(new_n746), .A2(new_n563), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g559(.A1(new_n244), .A2(new_n604), .A3(new_n661), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n580), .B(new_n761), .C1(new_n704), .C2(new_n715), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT51), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT118), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n765), .B(new_n638), .C1(new_n705), .C2(new_n709), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n244), .A2(new_n604), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n523), .A2(new_n578), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n765), .B1(new_n769), .B2(new_n638), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n764), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n713), .A2(KEYINPUT118), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n772), .A2(KEYINPUT51), .A3(new_n767), .A4(new_n766), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n660), .A2(new_n580), .A3(new_n613), .ZN(new_n775));
  OAI22_X1  g574(.A1(new_n763), .A2(new_n613), .B1(new_n774), .B2(new_n775), .ZN(G1336gat));
  OAI211_X1 g575(.A(new_n526), .B(new_n761), .C1(new_n704), .C2(new_n715), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(G92gat), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT119), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n771), .A2(new_n773), .A3(new_n779), .ZN(new_n780));
  OAI211_X1 g579(.A(KEYINPUT119), .B(new_n764), .C1(new_n768), .C2(new_n770), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n661), .A2(G92gat), .A3(new_n332), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n778), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(KEYINPUT52), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n786));
  INV_X1    g585(.A(new_n782), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n778), .B(new_n786), .C1(new_n774), .C2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n785), .A2(new_n788), .ZN(G1337gat));
  OAI21_X1  g588(.A(new_n761), .B1(new_n704), .B2(new_n715), .ZN(new_n790));
  OAI21_X1  g589(.A(G99gat), .B1(new_n790), .B2(new_n679), .ZN(new_n791));
  INV_X1    g590(.A(G99gat), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n461), .A2(new_n660), .A3(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n791), .B1(new_n774), .B2(new_n793), .ZN(G1338gat));
  OAI211_X1 g593(.A(new_n563), .B(new_n761), .C1(new_n704), .C2(new_n715), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(G106gat), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n661), .A2(G106gat), .A3(new_n481), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n780), .A2(new_n781), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT53), .ZN(new_n800));
  XNOR2_X1  g599(.A(KEYINPUT120), .B(KEYINPUT53), .ZN(new_n801));
  INV_X1    g600(.A(new_n797), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n796), .B(new_n801), .C1(new_n774), .C2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n800), .A2(new_n803), .ZN(G1339gat));
  NOR2_X1   g603(.A1(new_n232), .A2(new_n233), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n227), .A2(new_n228), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n240), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n242), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n660), .ZN(new_n809));
  OR2_X1    g608(.A1(new_n651), .A2(KEYINPUT54), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n644), .A2(new_n649), .A3(new_n645), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n651), .A2(KEYINPUT54), .A3(new_n811), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n810), .A2(new_n657), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(KEYINPUT55), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n814), .B1(new_n652), .B2(new_n657), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n813), .A2(KEYINPUT55), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n244), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n809), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n702), .ZN(new_n820));
  INV_X1    g619(.A(new_n702), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n821), .A2(new_n808), .A3(new_n817), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n604), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n662), .A2(new_n244), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n825), .A2(new_n526), .A3(new_n495), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n517), .A2(new_n518), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OR3_X1    g627(.A1(new_n828), .A2(new_n245), .A3(new_n342), .ZN(new_n829));
  INV_X1    g628(.A(new_n825), .ZN(new_n830));
  INV_X1    g629(.A(new_n482), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n526), .A2(new_n495), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT121), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n826), .A2(KEYINPUT121), .A3(new_n831), .ZN(new_n836));
  AND3_X1   g635(.A1(new_n835), .A2(new_n836), .A3(new_n244), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n829), .B1(new_n837), .B2(new_n337), .ZN(G1340gat));
  NAND3_X1  g637(.A1(new_n835), .A2(new_n836), .A3(new_n660), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT122), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n839), .A2(new_n840), .A3(G120gat), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n840), .B1(new_n839), .B2(G120gat), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n660), .A2(new_n338), .ZN(new_n843));
  OAI22_X1  g642(.A1(new_n841), .A2(new_n842), .B1(new_n828), .B2(new_n843), .ZN(G1341gat));
  NAND4_X1  g643(.A1(new_n835), .A2(new_n836), .A3(G127gat), .A4(new_n604), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n845), .A2(KEYINPUT123), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n845), .A2(KEYINPUT123), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n828), .A2(new_n688), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n848), .A2(G127gat), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n846), .A2(new_n847), .A3(new_n849), .ZN(G1342gat));
  NOR3_X1   g649(.A1(new_n828), .A2(G134gat), .A3(new_n639), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(KEYINPUT56), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n835), .A2(new_n836), .A3(new_n638), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(G134gat), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n852), .A2(new_n854), .ZN(G1343gat));
  NOR2_X1   g654(.A1(new_n576), .A2(new_n481), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n826), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n857), .A2(new_n356), .A3(new_n244), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT58), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n679), .A2(new_n832), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT124), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n638), .B1(new_n819), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n809), .A2(new_n818), .A3(KEYINPUT124), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n604), .B1(new_n864), .B2(new_n822), .ZN(new_n865));
  OAI211_X1 g664(.A(KEYINPUT57), .B(new_n563), .C1(new_n865), .C2(new_n824), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n867), .B1(new_n825), .B2(new_n481), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n860), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n869), .A2(new_n244), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n858), .B(new_n859), .C1(new_n870), .C2(new_n372), .ZN(new_n871));
  INV_X1    g670(.A(new_n858), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n372), .B1(new_n869), .B2(new_n244), .ZN(new_n873));
  OAI21_X1  g672(.A(KEYINPUT58), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n871), .A2(new_n874), .ZN(G1344gat));
  INV_X1    g674(.A(G148gat), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n857), .A2(new_n876), .A3(new_n660), .ZN(new_n877));
  AOI211_X1 g676(.A(KEYINPUT59), .B(new_n876), .C1(new_n869), .C2(new_n660), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT59), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n860), .A2(new_n661), .ZN(new_n880));
  AND3_X1   g679(.A1(new_n808), .A2(new_n817), .A3(new_n638), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n881), .B1(new_n862), .B2(new_n863), .ZN(new_n882));
  OAI22_X1  g681(.A1(new_n882), .A2(new_n604), .B1(new_n244), .B2(new_n662), .ZN(new_n883));
  AOI21_X1  g682(.A(KEYINPUT57), .B1(new_n883), .B2(new_n563), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n825), .A2(new_n867), .A3(new_n481), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n880), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n879), .B1(new_n886), .B2(G148gat), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n877), .B1(new_n878), .B2(new_n887), .ZN(G1345gat));
  INV_X1    g687(.A(G155gat), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n857), .A2(new_n889), .A3(new_n604), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n869), .A2(new_n604), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n890), .B1(new_n891), .B2(new_n889), .ZN(G1346gat));
  INV_X1    g691(.A(G162gat), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n857), .A2(new_n893), .A3(new_n638), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n869), .A2(new_n821), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT125), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(G162gat), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n895), .A2(new_n896), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n894), .B1(new_n898), .B2(new_n899), .ZN(G1347gat));
  NOR3_X1   g699(.A1(new_n825), .A2(new_n332), .A3(new_n580), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n901), .A2(new_n827), .ZN(new_n902));
  AOI21_X1  g701(.A(G169gat), .B1(new_n902), .B2(new_n244), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n831), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n904), .A2(new_n251), .A3(new_n245), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n903), .A2(new_n905), .ZN(G1348gat));
  NAND3_X1  g705(.A1(new_n902), .A2(new_n252), .A3(new_n660), .ZN(new_n907));
  OAI21_X1  g706(.A(G176gat), .B1(new_n904), .B2(new_n661), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(G1349gat));
  NAND3_X1  g708(.A1(new_n902), .A2(new_n247), .A3(new_n604), .ZN(new_n910));
  OAI21_X1  g709(.A(G183gat), .B1(new_n904), .B2(new_n688), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g712(.A1(new_n902), .A2(new_n248), .A3(new_n821), .ZN(new_n914));
  OAI21_X1  g713(.A(G190gat), .B1(new_n904), .B2(new_n639), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n915), .A2(KEYINPUT61), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n915), .A2(KEYINPUT61), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n914), .B1(new_n916), .B2(new_n917), .ZN(G1351gat));
  NOR3_X1   g717(.A1(new_n576), .A2(new_n332), .A3(new_n580), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n919), .B1(new_n884), .B2(new_n885), .ZN(new_n920));
  OAI21_X1  g719(.A(G197gat), .B1(new_n920), .B2(new_n245), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n901), .A2(new_n856), .ZN(new_n922));
  INV_X1    g721(.A(G197gat), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n922), .A2(new_n923), .A3(new_n244), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n924), .A2(KEYINPUT126), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n924), .A2(KEYINPUT126), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n921), .B1(new_n925), .B2(new_n926), .ZN(G1352gat));
  INV_X1    g726(.A(G204gat), .ZN(new_n928));
  OAI211_X1 g727(.A(new_n660), .B(new_n919), .C1(new_n884), .C2(new_n885), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n928), .B1(new_n929), .B2(KEYINPUT127), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n930), .B1(KEYINPUT127), .B2(new_n929), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n901), .A2(new_n928), .A3(new_n660), .A4(new_n856), .ZN(new_n932));
  XOR2_X1   g731(.A(new_n932), .B(KEYINPUT62), .Z(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(new_n933), .ZN(G1353gat));
  NAND3_X1  g733(.A1(new_n922), .A2(new_n288), .A3(new_n604), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n604), .B(new_n919), .C1(new_n884), .C2(new_n885), .ZN(new_n936));
  AND3_X1   g735(.A1(new_n936), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n937));
  AOI21_X1  g736(.A(KEYINPUT63), .B1(new_n936), .B2(G211gat), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n935), .B1(new_n937), .B2(new_n938), .ZN(G1354gat));
  OAI21_X1  g738(.A(G218gat), .B1(new_n920), .B2(new_n639), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n922), .A2(new_n289), .A3(new_n821), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(G1355gat));
endmodule


