//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 0 1 1 0 1 0 0 1 0 0 0 1 1 0 0 0 0 0 1 1 0 1 0 0 1 0 0 1 0 1 0 0 0 0 1 0 0 1 0 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:17 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n552, new_n553, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n579, new_n580, new_n581, new_n582,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n623, new_n625, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT66), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT67), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(G325));
  XOR2_X1   g030(.A(new_n454), .B(KEYINPUT68), .Z(G261));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n452), .A2(new_n457), .B1(new_n458), .B2(new_n453), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT69), .Z(G319));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n464), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  INV_X1    g046(.A(G137), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n462), .A2(KEYINPUT70), .A3(G2104), .ZN(new_n473));
  AND2_X1   g048(.A1(new_n473), .A2(new_n465), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT70), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n463), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n474), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n469), .B(new_n471), .C1(new_n472), .C2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n475), .ZN(new_n482));
  INV_X1    g057(.A(G136), .ZN(new_n483));
  INV_X1    g058(.A(G124), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n474), .A2(G2105), .A3(new_n477), .ZN(new_n485));
  OAI221_X1 g060(.A(new_n482), .B1(new_n478), .B2(new_n483), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  INV_X1    g062(.A(KEYINPUT71), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(G114), .ZN(new_n489));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(KEYINPUT71), .ZN(new_n491));
  OAI21_X1  g066(.A(G2105), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(G126), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n495), .B1(new_n485), .B2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(G138), .ZN(new_n498));
  OAI21_X1  g073(.A(KEYINPUT4), .B1(new_n478), .B2(new_n498), .ZN(new_n499));
  OR4_X1    g074(.A1(KEYINPUT4), .A2(new_n466), .A3(new_n498), .A4(G2105), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n497), .B1(new_n499), .B2(new_n500), .ZN(G164));
  AND2_X1   g076(.A1(G75), .A2(G543), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n503), .B1(new_n504), .B2(KEYINPUT72), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT72), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(KEYINPUT5), .A3(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n502), .B1(new_n508), .B2(G62), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT73), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  OR3_X1    g086(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(G50), .A2(G543), .ZN(new_n513));
  AND2_X1   g088(.A1(new_n505), .A2(new_n507), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT6), .B(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n510), .B1(new_n509), .B2(new_n511), .ZN(new_n519));
  AND3_X1   g094(.A1(new_n512), .A2(new_n518), .A3(new_n519), .ZN(G166));
  OR2_X1    g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n521), .A2(KEYINPUT74), .A3(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT74), .ZN(new_n524));
  AND2_X1   g099(.A1(KEYINPUT6), .A2(G651), .ZN(new_n525));
  NOR2_X1   g100(.A1(KEYINPUT6), .A2(G651), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n523), .A2(new_n527), .A3(G51), .A4(G543), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n508), .A2(G89), .A3(new_n517), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n508), .A2(G63), .A3(G651), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  AND4_X1   g107(.A1(new_n528), .A2(new_n529), .A3(new_n530), .A4(new_n532), .ZN(G168));
  INV_X1    g108(.A(G64), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n534), .B1(new_n505), .B2(new_n507), .ZN(new_n535));
  AND2_X1   g110(.A1(G77), .A2(G543), .ZN(new_n536));
  OAI21_X1  g111(.A(G651), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n523), .A2(new_n527), .A3(G52), .A4(G543), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n508), .A2(G90), .A3(new_n517), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  AOI21_X1  g116(.A(new_n504), .B1(new_n517), .B2(new_n524), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n542), .A2(G43), .A3(new_n523), .ZN(new_n543));
  INV_X1    g118(.A(G56), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n544), .B1(new_n505), .B2(new_n507), .ZN(new_n545));
  AND2_X1   g120(.A1(G68), .A2(G543), .ZN(new_n546));
  OAI21_X1  g121(.A(G651), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n508), .A2(G81), .A3(new_n517), .ZN(new_n548));
  AND3_X1   g123(.A1(new_n543), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  INV_X1    g129(.A(KEYINPUT77), .ZN(new_n555));
  NAND4_X1  g130(.A1(new_n523), .A2(new_n527), .A3(G53), .A4(G543), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT9), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n557), .A2(KEYINPUT75), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n558), .ZN(new_n560));
  NAND4_X1  g135(.A1(new_n542), .A2(G53), .A3(new_n523), .A4(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(KEYINPUT76), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT76), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n559), .A2(new_n561), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G65), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n514), .B2(new_n568), .ZN(new_n569));
  AND2_X1   g144(.A1(new_n508), .A2(new_n517), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n569), .A2(G651), .B1(new_n570), .B2(G91), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n555), .B1(new_n566), .B2(new_n571), .ZN(new_n572));
  AND3_X1   g147(.A1(new_n559), .A2(new_n561), .A3(new_n564), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n564), .B1(new_n559), .B2(new_n561), .ZN(new_n574));
  OAI211_X1 g149(.A(new_n555), .B(new_n571), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n572), .A2(new_n576), .ZN(G299));
  INV_X1    g152(.A(G168), .ZN(G286));
  INV_X1    g153(.A(KEYINPUT78), .ZN(new_n579));
  NAND2_X1  g154(.A1(G166), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n512), .A2(new_n518), .A3(new_n519), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(KEYINPUT78), .ZN(new_n582));
  AND2_X1   g157(.A1(new_n580), .A2(new_n582), .ZN(G303));
  AND2_X1   g158(.A1(new_n542), .A2(new_n523), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(G49), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n570), .A2(G87), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(G288));
  AND2_X1   g163(.A1(new_n508), .A2(G61), .ZN(new_n589));
  NAND2_X1  g164(.A1(G73), .A2(G543), .ZN(new_n590));
  XOR2_X1   g165(.A(new_n590), .B(KEYINPUT79), .Z(new_n591));
  OAI21_X1  g166(.A(G651), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(G48), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G86), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n514), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(new_n517), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n592), .A2(new_n596), .ZN(G305));
  NAND2_X1  g172(.A1(new_n584), .A2(G47), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n570), .A2(G85), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  OAI211_X1 g175(.A(new_n598), .B(new_n599), .C1(new_n511), .C2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT80), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n601), .B(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(G301), .A2(G868), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT81), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n570), .A2(new_n605), .A3(G92), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n508), .A2(new_n517), .ZN(new_n607));
  INV_X1    g182(.A(G92), .ZN(new_n608));
  OAI21_X1  g183(.A(KEYINPUT81), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n606), .A2(KEYINPUT10), .A3(new_n609), .ZN(new_n613));
  NAND2_X1  g188(.A1(G79), .A2(G543), .ZN(new_n614));
  INV_X1    g189(.A(G66), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n514), .B2(new_n615), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n584), .A2(G54), .B1(new_n616), .B2(G651), .ZN(new_n617));
  AND3_X1   g192(.A1(new_n612), .A2(new_n613), .A3(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n604), .B1(new_n618), .B2(G868), .ZN(G284));
  OAI21_X1  g194(.A(new_n604), .B1(new_n618), .B2(G868), .ZN(G321));
  MUX2_X1   g195(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g196(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n618), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND3_X1  g199(.A1(new_n543), .A2(new_n547), .A3(new_n548), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n618), .A2(new_n623), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT82), .Z(new_n627));
  MUX2_X1   g202(.A(new_n625), .B(new_n627), .S(G868), .Z(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g204(.A(G123), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n485), .A2(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(KEYINPUT84), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n634));
  INV_X1    g209(.A(G111), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n634), .B1(new_n635), .B2(G2105), .ZN(new_n636));
  INV_X1    g211(.A(new_n478), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n636), .B1(new_n637), .B2(G135), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n633), .A2(new_n638), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n639), .A2(G2096), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(G2096), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n475), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT12), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2100), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT83), .B(KEYINPUT13), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n640), .A2(new_n641), .A3(new_n646), .ZN(G156));
  XNOR2_X1  g222(.A(KEYINPUT15), .B(G2435), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT85), .B(G2438), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G2427), .B(G2430), .Z(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(KEYINPUT14), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2443), .B(G2446), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1341), .B(G1348), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2451), .B(G2454), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT16), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT86), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n662), .A2(G14), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n658), .A2(new_n661), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT87), .Z(G401));
  INV_X1    g241(.A(KEYINPUT18), .ZN(new_n667));
  XOR2_X1   g242(.A(G2084), .B(G2090), .Z(new_n668));
  XNOR2_X1  g243(.A(G2067), .B(G2678), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n670), .A2(KEYINPUT17), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n668), .A2(new_n669), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n667), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(G2100), .ZN(new_n674));
  XOR2_X1   g249(.A(G2072), .B(G2078), .Z(new_n675));
  AOI21_X1  g250(.A(new_n675), .B1(new_n670), .B2(KEYINPUT18), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(G2096), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n674), .B(new_n677), .ZN(G227));
  XNOR2_X1  g253(.A(G1971), .B(G1976), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n682), .A2(KEYINPUT90), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1956), .B(G2474), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1961), .B(G1966), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n684), .A2(new_n685), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n686), .B1(new_n681), .B2(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n683), .B(new_n688), .Z(new_n689));
  INV_X1    g264(.A(KEYINPUT89), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n687), .A2(new_n690), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n691), .A2(new_n681), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT20), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n689), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1991), .B(G1996), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1981), .B(G1986), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n699), .B(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(G229));
  INV_X1    g278(.A(G16), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G21), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G168), .B2(new_n704), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT96), .Z(new_n707));
  INV_X1    g282(.A(G1966), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT97), .ZN(new_n710));
  INV_X1    g285(.A(G29), .ZN(new_n711));
  OR3_X1    g286(.A1(new_n639), .A2(KEYINPUT98), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g287(.A(KEYINPUT98), .B1(new_n639), .B2(new_n711), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT31), .B(G11), .Z(new_n714));
  INV_X1    g289(.A(KEYINPUT30), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n711), .B1(new_n715), .B2(G28), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n716), .A2(KEYINPUT99), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(new_n715), .B2(G28), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n716), .A2(KEYINPUT99), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n714), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(G5), .A2(G16), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT100), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G301), .B2(new_n704), .ZN(new_n723));
  INV_X1    g298(.A(G1961), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g300(.A1(new_n712), .A2(new_n713), .A3(new_n720), .A4(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(new_n708), .B2(new_n707), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n710), .A2(new_n727), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT101), .Z(new_n729));
  NAND2_X1  g304(.A1(G299), .A2(G16), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n704), .A2(G20), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT23), .ZN(new_n732));
  AND3_X1   g307(.A1(new_n730), .A2(G1956), .A3(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(G1956), .B1(new_n730), .B2(new_n732), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n711), .A2(G33), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT25), .Z(new_n738));
  INV_X1    g313(.A(G139), .ZN(new_n739));
  INV_X1    g314(.A(G127), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n466), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G115), .B2(G2104), .ZN(new_n742));
  OAI221_X1 g317(.A(new_n738), .B1(new_n739), .B2(new_n478), .C1(new_n742), .C2(new_n475), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n736), .B1(new_n743), .B2(G29), .ZN(new_n744));
  INV_X1    g319(.A(G2072), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT95), .Z(new_n747));
  XOR2_X1   g322(.A(KEYINPUT103), .B(G2078), .Z(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT104), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n711), .A2(G27), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT102), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n499), .A2(new_n500), .ZN(new_n752));
  INV_X1    g327(.A(new_n497), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n751), .B1(new_n754), .B2(G29), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n747), .B1(new_n749), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n704), .A2(G4), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n618), .B2(new_n704), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT93), .B(G1348), .Z(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n756), .B(new_n760), .C1(new_n749), .C2(new_n755), .ZN(new_n761));
  XOR2_X1   g336(.A(KEYINPUT94), .B(KEYINPUT24), .Z(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G34), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n763), .A2(new_n711), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n479), .B2(new_n711), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G2084), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n723), .A2(new_n724), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n744), .A2(new_n745), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n711), .A2(G35), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G162), .B2(new_n711), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT105), .B(KEYINPUT29), .ZN(new_n772));
  INV_X1    g347(.A(G2090), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n771), .B(new_n774), .Z(new_n775));
  NAND2_X1  g350(.A1(new_n711), .A2(G26), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT28), .ZN(new_n777));
  OR2_X1    g352(.A1(G104), .A2(G2105), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n778), .B(G2104), .C1(G116), .C2(new_n475), .ZN(new_n779));
  INV_X1    g354(.A(G140), .ZN(new_n780));
  INV_X1    g355(.A(G128), .ZN(new_n781));
  OAI221_X1 g356(.A(new_n779), .B1(new_n478), .B2(new_n780), .C1(new_n781), .C2(new_n485), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n777), .B1(new_n783), .B2(new_n711), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(G2067), .Z(new_n785));
  NAND2_X1  g360(.A1(new_n704), .A2(G19), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(new_n549), .B2(new_n704), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(G1341), .Z(new_n788));
  NAND2_X1  g363(.A1(new_n711), .A2(G32), .ZN(new_n789));
  NAND3_X1  g364(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT26), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n790), .A2(new_n791), .ZN(new_n793));
  AOI22_X1  g368(.A1(new_n792), .A2(new_n793), .B1(G105), .B2(new_n470), .ZN(new_n794));
  INV_X1    g369(.A(G129), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(new_n485), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G141), .B2(new_n637), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n789), .B1(new_n797), .B2(new_n711), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT27), .B(G1996), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n775), .A2(new_n785), .A3(new_n788), .A4(new_n800), .ZN(new_n801));
  NOR3_X1   g376(.A1(new_n761), .A2(new_n769), .A3(new_n801), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n729), .A2(new_n735), .A3(new_n802), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n704), .A2(G24), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(G290), .B2(G16), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n806), .A2(G1986), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n711), .A2(G25), .ZN(new_n808));
  INV_X1    g383(.A(G119), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n485), .A2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT91), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  OAI21_X1  g387(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n813));
  INV_X1    g388(.A(G107), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n813), .B1(new_n814), .B2(G2105), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(new_n637), .B2(G131), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n812), .A2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n808), .B1(new_n818), .B2(new_n711), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT35), .B(G1991), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n806), .A2(G1986), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n807), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(G6), .A2(G16), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n592), .A2(new_n596), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n824), .B1(new_n825), .B2(G16), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT32), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(G1981), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n704), .A2(G23), .ZN(new_n829));
  INV_X1    g404(.A(G288), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n829), .B1(new_n830), .B2(new_n704), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT33), .B(G1976), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(G166), .A2(G16), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(G16), .B2(G22), .ZN(new_n835));
  INV_X1    g410(.A(G1971), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n835), .A2(new_n836), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n833), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  OR3_X1    g414(.A1(new_n828), .A2(KEYINPUT92), .A3(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(KEYINPUT92), .B1(new_n828), .B2(new_n839), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT34), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n823), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n840), .A2(KEYINPUT34), .A3(new_n841), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(KEYINPUT36), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT36), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n844), .A2(new_n848), .A3(new_n845), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n803), .B1(new_n847), .B2(new_n849), .ZN(G311));
  INV_X1    g425(.A(G311), .ZN(G150));
  NAND2_X1  g426(.A1(new_n618), .A2(G559), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT38), .ZN(new_n853));
  AOI22_X1  g428(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n854), .A2(new_n511), .ZN(new_n855));
  NAND4_X1  g430(.A1(new_n523), .A2(new_n527), .A3(G55), .A4(G543), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n508), .A2(G93), .A3(new_n517), .ZN(new_n857));
  AND3_X1   g432(.A1(new_n856), .A2(KEYINPUT106), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(KEYINPUT106), .B1(new_n856), .B2(new_n857), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n855), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(new_n625), .ZN(new_n861));
  OAI211_X1 g436(.A(new_n549), .B(new_n855), .C1(new_n859), .C2(new_n858), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n853), .B(new_n864), .ZN(new_n865));
  AND2_X1   g440(.A1(new_n865), .A2(KEYINPUT39), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(KEYINPUT39), .ZN(new_n867));
  NOR3_X1   g442(.A1(new_n866), .A2(new_n867), .A3(G860), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n860), .A2(G860), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT37), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n868), .A2(new_n870), .ZN(G145));
  XNOR2_X1  g446(.A(G164), .B(new_n782), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n872), .A2(new_n797), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n743), .A2(KEYINPUT108), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n797), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n743), .A2(KEYINPUT108), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n877), .ZN(new_n879));
  NAND4_X1  g454(.A1(new_n873), .A2(new_n879), .A3(new_n874), .A4(new_n875), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n817), .B(new_n643), .ZN(new_n882));
  INV_X1    g457(.A(G130), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT109), .ZN(new_n884));
  NOR3_X1   g459(.A1(new_n884), .A2(new_n475), .A3(G118), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n884), .B1(new_n475), .B2(G118), .ZN(new_n886));
  OR2_X1    g461(.A1(G106), .A2(G2105), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n886), .A2(G2104), .A3(new_n887), .ZN(new_n888));
  OAI22_X1  g463(.A1(new_n485), .A2(new_n883), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n889), .B1(G142), .B2(new_n637), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n882), .B(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n881), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n891), .A2(new_n878), .A3(new_n880), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  XOR2_X1   g470(.A(new_n479), .B(KEYINPUT107), .Z(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(new_n486), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(new_n639), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(G37), .B1(new_n895), .B2(new_n899), .ZN(new_n900));
  AND2_X1   g475(.A1(new_n893), .A2(new_n894), .ZN(new_n901));
  AOI21_X1  g476(.A(KEYINPUT110), .B1(new_n901), .B2(new_n898), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT110), .ZN(new_n903));
  NOR3_X1   g478(.A1(new_n895), .A2(new_n903), .A3(new_n899), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n900), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g481(.A(G290), .B(new_n581), .ZN(new_n907));
  XNOR2_X1  g482(.A(G288), .B(G305), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n907), .B(new_n908), .ZN(new_n909));
  XOR2_X1   g484(.A(new_n909), .B(KEYINPUT42), .Z(new_n910));
  XNOR2_X1  g485(.A(new_n627), .B(new_n864), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT111), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT41), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n571), .B1(new_n573), .B2(new_n574), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT77), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n915), .A2(new_n575), .A3(new_n618), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n618), .B1(new_n915), .B2(new_n575), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n913), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n618), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n919), .B1(new_n572), .B2(new_n576), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n915), .A2(new_n575), .A3(new_n618), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n920), .A2(KEYINPUT41), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n912), .B1(new_n918), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n916), .A2(new_n917), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT111), .B1(new_n924), .B2(KEYINPUT41), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n911), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n926), .B1(new_n911), .B2(new_n924), .ZN(new_n927));
  AND2_X1   g502(.A1(new_n910), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n910), .A2(new_n927), .ZN(new_n929));
  OAI21_X1  g504(.A(G868), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n860), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n930), .B1(G868), .B2(new_n931), .ZN(G295));
  OAI21_X1  g507(.A(new_n930), .B1(G868), .B2(new_n931), .ZN(G331));
  NAND4_X1  g508(.A1(new_n537), .A2(KEYINPUT112), .A3(new_n538), .A4(new_n539), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT113), .ZN(new_n935));
  AND3_X1   g510(.A1(G168), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n935), .B1(G168), .B2(new_n934), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n863), .A2(new_n938), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n861), .B(new_n862), .C1(new_n937), .C2(new_n936), .ZN(new_n940));
  NOR2_X1   g515(.A1(G171), .A2(KEYINPUT112), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n941), .B1(new_n939), .B2(new_n940), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n945), .B1(new_n923), .B2(new_n925), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n939), .A2(new_n940), .ZN(new_n947));
  INV_X1    g522(.A(new_n941), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AOI22_X1  g524(.A1(new_n949), .A2(new_n942), .B1(new_n921), .B2(new_n920), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n946), .A2(new_n909), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT114), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT114), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n946), .A2(new_n909), .A3(new_n954), .A4(new_n951), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n909), .B1(new_n946), .B2(new_n951), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n957), .A2(G37), .ZN(new_n958));
  AOI21_X1  g533(.A(KEYINPUT43), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT43), .ZN(new_n960));
  INV_X1    g535(.A(G37), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n918), .A2(new_n922), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n950), .B1(new_n962), .B2(new_n945), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n961), .B1(new_n963), .B2(new_n909), .ZN(new_n964));
  AOI211_X1 g539(.A(new_n960), .B(new_n964), .C1(new_n953), .C2(new_n955), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT44), .B1(new_n959), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT44), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n960), .B1(new_n956), .B2(new_n958), .ZN(new_n968));
  AOI211_X1 g543(.A(KEYINPUT43), .B(new_n964), .C1(new_n953), .C2(new_n955), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n966), .A2(new_n970), .ZN(G397));
  INV_X1    g546(.A(KEYINPUT45), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n972), .B1(G164), .B2(G1384), .ZN(new_n973));
  INV_X1    g548(.A(G40), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n479), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n782), .B(G2067), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n979), .B(KEYINPUT115), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n797), .B(G1996), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n817), .B(new_n820), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n978), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  XNOR2_X1  g559(.A(G290), .B(G1986), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n984), .B1(new_n977), .B2(new_n985), .ZN(new_n986));
  XOR2_X1   g561(.A(new_n986), .B(KEYINPUT116), .Z(new_n987));
  INV_X1    g562(.A(KEYINPUT117), .ZN(new_n988));
  AOI21_X1  g563(.A(G1384), .B1(new_n752), .B2(new_n753), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n975), .B1(new_n989), .B2(KEYINPUT45), .ZN(new_n990));
  NOR3_X1   g565(.A1(G164), .A2(new_n972), .A3(G1384), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n988), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n989), .A2(KEYINPUT45), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n993), .A2(new_n973), .A3(KEYINPUT117), .A4(new_n975), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n992), .A2(new_n836), .A3(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(G1384), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n754), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT50), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT50), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n989), .A2(new_n999), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n998), .A2(new_n773), .A3(new_n1000), .A4(new_n975), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n995), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(G8), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n580), .A2(G8), .A3(new_n582), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n1005));
  OR3_X1    g580(.A1(new_n1004), .A2(KEYINPUT118), .A3(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT118), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1008));
  AND3_X1   g583(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1003), .A2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g585(.A(KEYINPUT119), .B(G1981), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n825), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(G305), .A2(G1981), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT49), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G8), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1017), .B1(new_n989), .B2(new_n975), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1012), .A2(KEYINPUT49), .A3(new_n1013), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1016), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n830), .A2(G1976), .ZN(new_n1021));
  INV_X1    g596(.A(G1976), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT52), .B1(G288), .B2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1018), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1020), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(KEYINPUT52), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1025), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1030), .A2(new_n1002), .A3(G8), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n1010), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT54), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT53), .ZN(new_n1034));
  AND2_X1   g609(.A1(new_n992), .A2(new_n994), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1034), .B1(new_n1035), .B2(G2078), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n993), .A2(new_n975), .A3(new_n973), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1034), .A2(G2078), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n998), .A2(new_n1000), .A3(new_n975), .ZN(new_n1040));
  AOI22_X1  g615(.A1(new_n1038), .A2(new_n1039), .B1(new_n1040), .B2(new_n724), .ZN(new_n1041));
  AOI21_X1  g616(.A(G301), .B1(new_n1036), .B2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(G2078), .B1(new_n992), .B2(new_n994), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n1041), .B(G301), .C1(new_n1043), .C2(KEYINPUT53), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1033), .B1(new_n1042), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT126), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1037), .A2(new_n708), .ZN(new_n1048));
  XNOR2_X1  g623(.A(KEYINPUT122), .B(G2084), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n998), .A2(new_n1000), .A3(new_n975), .A4(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1047), .B(G8), .C1(new_n1051), .C2(G286), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT51), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1017), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1055));
  NOR2_X1   g630(.A1(G168), .A2(new_n1017), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1047), .B(KEYINPUT51), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1054), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1051), .A2(new_n1056), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1041), .B1(new_n1043), .B2(KEYINPUT53), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(G171), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1062), .A2(KEYINPUT54), .A3(new_n1044), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1032), .A2(new_n1046), .A3(new_n1060), .A4(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT125), .ZN(new_n1065));
  INV_X1    g640(.A(G1996), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1038), .A2(KEYINPUT124), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT124), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1068), .B1(new_n1037), .B2(G1996), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n989), .A2(new_n975), .ZN(new_n1071));
  XOR2_X1   g646(.A(KEYINPUT58), .B(G1341), .Z(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1065), .B1(new_n1070), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1073), .ZN(new_n1075));
  AOI211_X1 g650(.A(KEYINPUT125), .B(new_n1075), .C1(new_n1067), .C2(new_n1069), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n549), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT59), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT61), .ZN(new_n1080));
  XNOR2_X1  g655(.A(KEYINPUT56), .B(G2072), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1038), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n571), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1083), .A2(KEYINPUT57), .ZN(new_n1084));
  AOI22_X1  g659(.A1(new_n914), .A2(KEYINPUT57), .B1(new_n1084), .B2(new_n562), .ZN(new_n1085));
  INV_X1    g660(.A(G1956), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1040), .A2(new_n1086), .ZN(new_n1087));
  AND3_X1   g662(.A1(new_n1082), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1085), .B1(new_n1082), .B2(new_n1087), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1080), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1071), .A2(G2067), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1091), .B1(new_n1040), .B2(new_n759), .ZN(new_n1092));
  OR2_X1    g667(.A1(new_n1092), .A2(new_n618), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n618), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1093), .A2(KEYINPUT60), .A3(new_n1094), .ZN(new_n1095));
  OR2_X1    g670(.A1(new_n1094), .A2(KEYINPUT60), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n1090), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1082), .A2(new_n1087), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT123), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1085), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1100), .B1(new_n1099), .B2(new_n1098), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1088), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1101), .A2(KEYINPUT61), .A3(new_n1102), .ZN(new_n1103));
  OAI211_X1 g678(.A(KEYINPUT59), .B(new_n549), .C1(new_n1074), .C2(new_n1076), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1079), .A2(new_n1097), .A3(new_n1103), .A4(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1101), .B1(new_n919), .B2(new_n1092), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n1102), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1064), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  XOR2_X1   g683(.A(new_n1018), .B(KEYINPUT121), .Z(new_n1109));
  AND3_X1   g684(.A1(new_n1020), .A2(new_n1022), .A3(new_n830), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1012), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1109), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(KEYINPUT120), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT120), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1027), .A2(new_n1020), .A3(new_n1114), .A4(new_n1024), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1112), .B1(new_n1116), .B2(new_n1031), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n1055), .A2(G168), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1010), .A2(new_n1029), .A3(new_n1031), .A4(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT63), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1055), .A2(KEYINPUT63), .A3(G168), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1122), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1123), .A2(new_n1031), .A3(new_n1010), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1117), .B1(new_n1121), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1060), .A2(KEYINPUT62), .ZN(new_n1126));
  AND4_X1   g701(.A1(new_n1029), .A2(new_n1042), .A3(new_n1010), .A4(new_n1031), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT62), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1058), .A2(new_n1128), .A3(new_n1059), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1126), .A2(new_n1127), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1125), .A2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n987), .B1(new_n1108), .B2(new_n1131), .ZN(new_n1132));
  NOR3_X1   g707(.A1(new_n978), .A2(G290), .A3(G1986), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1133), .B(KEYINPUT48), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n984), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n977), .A2(KEYINPUT46), .A3(new_n1066), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT46), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1137), .B1(new_n978), .B2(G1996), .ZN(new_n1138));
  AND2_X1   g713(.A1(new_n980), .A2(new_n797), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1136), .B(new_n1138), .C1(new_n1139), .C2(new_n978), .ZN(new_n1140));
  XOR2_X1   g715(.A(new_n1140), .B(KEYINPUT47), .Z(new_n1141));
  NAND3_X1  g716(.A1(new_n982), .A2(new_n820), .A3(new_n818), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1142), .B1(G2067), .B2(new_n782), .ZN(new_n1143));
  AOI211_X1 g718(.A(new_n1135), .B(new_n1141), .C1(new_n977), .C2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1132), .A2(new_n1144), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g720(.A1(G227), .A2(new_n459), .ZN(new_n1147));
  OAI21_X1  g721(.A(new_n1147), .B1(new_n663), .B2(new_n664), .ZN(new_n1148));
  OR2_X1    g722(.A1(new_n1148), .A2(KEYINPUT127), .ZN(new_n1149));
  NAND2_X1  g723(.A1(new_n1148), .A2(KEYINPUT127), .ZN(new_n1150));
  AND3_X1   g724(.A1(new_n702), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  OAI211_X1 g725(.A(new_n905), .B(new_n1151), .C1(new_n968), .C2(new_n969), .ZN(G225));
  INV_X1    g726(.A(G225), .ZN(G308));
endmodule


