

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590;

  INV_X1 U324 ( .A(KEYINPUT32), .ZN(n335) );
  XNOR2_X1 U325 ( .A(n391), .B(n390), .ZN(n453) );
  XNOR2_X1 U326 ( .A(n357), .B(n356), .ZN(n360) );
  XNOR2_X1 U327 ( .A(n355), .B(G92GAT), .ZN(n356) );
  NOR2_X1 U328 ( .A1(n495), .A2(n448), .ZN(n546) );
  XNOR2_X1 U329 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U330 ( .A(n395), .B(n351), .ZN(n353) );
  XNOR2_X1 U331 ( .A(n454), .B(KEYINPUT118), .ZN(n455) );
  XNOR2_X1 U332 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U333 ( .A(n456), .B(n455), .ZN(n457) );
  INV_X1 U334 ( .A(KEYINPUT109), .ZN(n429) );
  XNOR2_X1 U335 ( .A(n338), .B(n337), .ZN(n342) );
  XNOR2_X1 U336 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U337 ( .A(n430), .B(n429), .ZN(n550) );
  XNOR2_X1 U338 ( .A(n461), .B(n460), .ZN(n462) );
  XOR2_X1 U339 ( .A(KEYINPUT36), .B(n384), .Z(n588) );
  XOR2_X1 U340 ( .A(n577), .B(KEYINPUT41), .Z(n563) );
  XNOR2_X1 U341 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U342 ( .A(n449), .B(G127GAT), .ZN(n450) );
  XNOR2_X1 U343 ( .A(n466), .B(n465), .ZN(G1351GAT) );
  XOR2_X1 U344 ( .A(G204GAT), .B(KEYINPUT83), .Z(n293) );
  XNOR2_X1 U345 ( .A(G218GAT), .B(KEYINPUT23), .ZN(n292) );
  XNOR2_X1 U346 ( .A(n293), .B(n292), .ZN(n308) );
  XOR2_X1 U347 ( .A(G211GAT), .B(KEYINPUT21), .Z(n295) );
  XNOR2_X1 U348 ( .A(G197GAT), .B(KEYINPUT82), .ZN(n294) );
  XNOR2_X1 U349 ( .A(n295), .B(n294), .ZN(n394) );
  XOR2_X1 U350 ( .A(G50GAT), .B(G162GAT), .Z(n352) );
  XOR2_X1 U351 ( .A(n394), .B(n352), .Z(n297) );
  NAND2_X1 U352 ( .A1(G228GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U353 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U354 ( .A(KEYINPUT24), .B(KEYINPUT81), .Z(n299) );
  XNOR2_X1 U355 ( .A(G22GAT), .B(KEYINPUT22), .ZN(n298) );
  XNOR2_X1 U356 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U357 ( .A(n301), .B(n300), .Z(n306) );
  XNOR2_X1 U358 ( .A(G106GAT), .B(G78GAT), .ZN(n302) );
  XNOR2_X1 U359 ( .A(n302), .B(G148GAT), .ZN(n334) );
  XOR2_X1 U360 ( .A(G155GAT), .B(KEYINPUT2), .Z(n304) );
  XNOR2_X1 U361 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n303) );
  XNOR2_X1 U362 ( .A(n304), .B(n303), .ZN(n421) );
  XNOR2_X1 U363 ( .A(n334), .B(n421), .ZN(n305) );
  XNOR2_X1 U364 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U365 ( .A(n308), .B(n307), .ZN(n474) );
  XOR2_X1 U366 ( .A(KEYINPUT28), .B(n474), .Z(n495) );
  XOR2_X1 U367 ( .A(G169GAT), .B(G8GAT), .Z(n401) );
  XOR2_X1 U368 ( .A(KEYINPUT68), .B(G1GAT), .Z(n310) );
  XNOR2_X1 U369 ( .A(G15GAT), .B(G22GAT), .ZN(n309) );
  XNOR2_X1 U370 ( .A(n310), .B(n309), .ZN(n376) );
  XOR2_X1 U371 ( .A(n401), .B(n376), .Z(n312) );
  XNOR2_X1 U372 ( .A(G36GAT), .B(G50GAT), .ZN(n311) );
  XNOR2_X1 U373 ( .A(n312), .B(n311), .ZN(n317) );
  XNOR2_X1 U374 ( .A(G29GAT), .B(KEYINPUT7), .ZN(n313) );
  XNOR2_X1 U375 ( .A(n313), .B(KEYINPUT8), .ZN(n354) );
  XOR2_X1 U376 ( .A(n354), .B(KEYINPUT66), .Z(n315) );
  NAND2_X1 U377 ( .A1(G229GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U378 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U379 ( .A(n317), .B(n316), .Z(n325) );
  XOR2_X1 U380 ( .A(G197GAT), .B(G141GAT), .Z(n319) );
  XNOR2_X1 U381 ( .A(G43GAT), .B(G113GAT), .ZN(n318) );
  XNOR2_X1 U382 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U383 ( .A(KEYINPUT30), .B(KEYINPUT65), .Z(n321) );
  XNOR2_X1 U384 ( .A(KEYINPUT29), .B(KEYINPUT67), .ZN(n320) );
  XNOR2_X1 U385 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U386 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U387 ( .A(n325), .B(n324), .ZN(n573) );
  INV_X1 U388 ( .A(G92GAT), .ZN(n326) );
  NAND2_X1 U389 ( .A1(G64GAT), .A2(n326), .ZN(n329) );
  INV_X1 U390 ( .A(G64GAT), .ZN(n327) );
  NAND2_X1 U391 ( .A1(n327), .A2(G92GAT), .ZN(n328) );
  NAND2_X1 U392 ( .A1(n329), .A2(n328), .ZN(n331) );
  XNOR2_X1 U393 ( .A(G176GAT), .B(G204GAT), .ZN(n330) );
  XNOR2_X1 U394 ( .A(n331), .B(n330), .ZN(n405) );
  XOR2_X1 U395 ( .A(G99GAT), .B(G85GAT), .Z(n358) );
  XNOR2_X1 U396 ( .A(n405), .B(n358), .ZN(n333) );
  AND2_X1 U397 ( .A1(G230GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U398 ( .A(n333), .B(n332), .ZN(n338) );
  XNOR2_X1 U399 ( .A(n334), .B(KEYINPUT31), .ZN(n336) );
  XOR2_X1 U400 ( .A(KEYINPUT71), .B(KEYINPUT70), .Z(n340) );
  XNOR2_X1 U401 ( .A(KEYINPUT69), .B(KEYINPUT33), .ZN(n339) );
  XNOR2_X1 U402 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U403 ( .A(n342), .B(n341), .ZN(n344) );
  XOR2_X1 U404 ( .A(G120GAT), .B(G71GAT), .Z(n433) );
  XOR2_X1 U405 ( .A(G57GAT), .B(KEYINPUT13), .Z(n372) );
  XOR2_X1 U406 ( .A(n433), .B(n372), .Z(n343) );
  XNOR2_X1 U407 ( .A(n344), .B(n343), .ZN(n577) );
  NAND2_X1 U408 ( .A1(n573), .A2(n563), .ZN(n345) );
  XNOR2_X1 U409 ( .A(KEYINPUT46), .B(n345), .ZN(n382) );
  XOR2_X1 U410 ( .A(KEYINPUT11), .B(KEYINPUT73), .Z(n347) );
  XNOR2_X1 U411 ( .A(KEYINPUT10), .B(KEYINPUT72), .ZN(n346) );
  XNOR2_X1 U412 ( .A(n347), .B(n346), .ZN(n362) );
  XNOR2_X1 U413 ( .A(G36GAT), .B(G190GAT), .ZN(n348) );
  XNOR2_X1 U414 ( .A(n348), .B(G218GAT), .ZN(n395) );
  NAND2_X1 U415 ( .A1(G232GAT), .A2(G233GAT), .ZN(n350) );
  INV_X1 U416 ( .A(KEYINPUT9), .ZN(n349) );
  XOR2_X1 U417 ( .A(n353), .B(n352), .Z(n357) );
  XOR2_X1 U418 ( .A(G43GAT), .B(G134GAT), .Z(n434) );
  XNOR2_X1 U419 ( .A(n354), .B(n434), .ZN(n355) );
  XOR2_X1 U420 ( .A(G106GAT), .B(n358), .Z(n359) );
  XNOR2_X1 U421 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U422 ( .A(n362), .B(n361), .ZN(n384) );
  XOR2_X1 U423 ( .A(G64GAT), .B(G211GAT), .Z(n364) );
  XNOR2_X1 U424 ( .A(G8GAT), .B(G155GAT), .ZN(n363) );
  XNOR2_X1 U425 ( .A(n364), .B(n363), .ZN(n368) );
  XOR2_X1 U426 ( .A(KEYINPUT76), .B(KEYINPUT12), .Z(n366) );
  XNOR2_X1 U427 ( .A(KEYINPUT14), .B(KEYINPUT15), .ZN(n365) );
  XNOR2_X1 U428 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U429 ( .A(n368), .B(n367), .ZN(n380) );
  XOR2_X1 U430 ( .A(G78GAT), .B(G71GAT), .Z(n370) );
  XNOR2_X1 U431 ( .A(G127GAT), .B(G183GAT), .ZN(n369) );
  XNOR2_X1 U432 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U433 ( .A(n372), .B(n371), .Z(n374) );
  NAND2_X1 U434 ( .A1(G231GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U435 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U436 ( .A(n375), .B(KEYINPUT75), .Z(n378) );
  XNOR2_X1 U437 ( .A(n376), .B(KEYINPUT74), .ZN(n377) );
  XNOR2_X1 U438 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U439 ( .A(n380), .B(n379), .ZN(n501) );
  INV_X1 U440 ( .A(n501), .ZN(n582) );
  NOR2_X1 U441 ( .A1(n384), .A2(n582), .ZN(n381) );
  AND2_X1 U442 ( .A1(n382), .A2(n381), .ZN(n383) );
  XNOR2_X1 U443 ( .A(n383), .B(KEYINPUT47), .ZN(n389) );
  NOR2_X1 U444 ( .A1(n501), .A2(n588), .ZN(n385) );
  XOR2_X1 U445 ( .A(KEYINPUT45), .B(n385), .Z(n386) );
  NOR2_X1 U446 ( .A1(n577), .A2(n386), .ZN(n387) );
  INV_X1 U447 ( .A(n573), .ZN(n518) );
  NAND2_X1 U448 ( .A1(n387), .A2(n518), .ZN(n388) );
  NAND2_X1 U449 ( .A1(n389), .A2(n388), .ZN(n391) );
  XNOR2_X1 U450 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n390) );
  XOR2_X1 U451 ( .A(G183GAT), .B(KEYINPUT17), .Z(n393) );
  XNOR2_X1 U452 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n392) );
  XNOR2_X1 U453 ( .A(n393), .B(n392), .ZN(n442) );
  XNOR2_X1 U454 ( .A(n442), .B(n394), .ZN(n399) );
  XOR2_X1 U455 ( .A(n395), .B(KEYINPUT90), .Z(n397) );
  NAND2_X1 U456 ( .A1(G226GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U457 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U458 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U459 ( .A(n400), .B(KEYINPUT89), .Z(n403) );
  XNOR2_X1 U460 ( .A(n401), .B(KEYINPUT74), .ZN(n402) );
  XNOR2_X1 U461 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U462 ( .A(n405), .B(n404), .ZN(n531) );
  XNOR2_X1 U463 ( .A(n531), .B(KEYINPUT27), .ZN(n476) );
  XOR2_X1 U464 ( .A(KEYINPUT85), .B(G57GAT), .Z(n407) );
  XNOR2_X1 U465 ( .A(G120GAT), .B(G148GAT), .ZN(n406) );
  XNOR2_X1 U466 ( .A(n407), .B(n406), .ZN(n411) );
  XOR2_X1 U467 ( .A(G85GAT), .B(G162GAT), .Z(n409) );
  XNOR2_X1 U468 ( .A(G29GAT), .B(G134GAT), .ZN(n408) );
  XNOR2_X1 U469 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U470 ( .A(n411), .B(n410), .ZN(n428) );
  XOR2_X1 U471 ( .A(KEYINPUT88), .B(KEYINPUT4), .Z(n413) );
  XNOR2_X1 U472 ( .A(KEYINPUT6), .B(KEYINPUT84), .ZN(n412) );
  XNOR2_X1 U473 ( .A(n413), .B(n412), .ZN(n417) );
  XOR2_X1 U474 ( .A(KEYINPUT1), .B(KEYINPUT86), .Z(n415) );
  XNOR2_X1 U475 ( .A(KEYINPUT5), .B(KEYINPUT87), .ZN(n414) );
  XNOR2_X1 U476 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U477 ( .A(n417), .B(n416), .Z(n426) );
  XOR2_X1 U478 ( .A(KEYINPUT0), .B(KEYINPUT78), .Z(n419) );
  XNOR2_X1 U479 ( .A(KEYINPUT77), .B(G127GAT), .ZN(n418) );
  XNOR2_X1 U480 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U481 ( .A(G113GAT), .B(n420), .Z(n445) );
  XOR2_X1 U482 ( .A(n421), .B(G1GAT), .Z(n423) );
  NAND2_X1 U483 ( .A1(G225GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U484 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U485 ( .A(n445), .B(n424), .ZN(n425) );
  XNOR2_X1 U486 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U487 ( .A(n428), .B(n427), .ZN(n481) );
  INV_X1 U488 ( .A(n481), .ZN(n529) );
  NOR2_X1 U489 ( .A1(n476), .A2(n529), .ZN(n468) );
  NAND2_X1 U490 ( .A1(n453), .A2(n468), .ZN(n430) );
  XOR2_X1 U491 ( .A(KEYINPUT79), .B(KEYINPUT20), .Z(n432) );
  XNOR2_X1 U492 ( .A(G169GAT), .B(G176GAT), .ZN(n431) );
  XNOR2_X1 U493 ( .A(n432), .B(n431), .ZN(n438) );
  INV_X1 U494 ( .A(G190GAT), .ZN(n463) );
  XOR2_X1 U495 ( .A(G99GAT), .B(G190GAT), .Z(n436) );
  XNOR2_X1 U496 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U497 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U498 ( .A(n438), .B(n437), .Z(n440) );
  NAND2_X1 U499 ( .A1(G227GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U500 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U501 ( .A(n441), .B(KEYINPUT80), .Z(n444) );
  XNOR2_X1 U502 ( .A(G15GAT), .B(n442), .ZN(n443) );
  XNOR2_X1 U503 ( .A(n444), .B(n443), .ZN(n446) );
  XNOR2_X1 U504 ( .A(n446), .B(n445), .ZN(n473) );
  INV_X1 U505 ( .A(n473), .ZN(n535) );
  NOR2_X1 U506 ( .A1(n550), .A2(n535), .ZN(n447) );
  XOR2_X1 U507 ( .A(KEYINPUT110), .B(n447), .Z(n448) );
  NAND2_X1 U508 ( .A1(n546), .A2(n582), .ZN(n451) );
  XOR2_X1 U509 ( .A(KEYINPUT50), .B(KEYINPUT111), .Z(n449) );
  XNOR2_X1 U510 ( .A(n451), .B(n450), .ZN(G1342GAT) );
  XOR2_X1 U511 ( .A(KEYINPUT116), .B(n531), .Z(n452) );
  NAND2_X1 U512 ( .A1(n453), .A2(n452), .ZN(n456) );
  XOR2_X1 U513 ( .A(KEYINPUT54), .B(KEYINPUT117), .Z(n454) );
  NOR2_X1 U514 ( .A1(n481), .A2(n457), .ZN(n570) );
  NAND2_X1 U515 ( .A1(n570), .A2(n474), .ZN(n461) );
  XOR2_X1 U516 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n459) );
  INV_X1 U517 ( .A(KEYINPUT55), .ZN(n458) );
  NOR2_X1 U518 ( .A1(n535), .A2(n462), .ZN(n568) );
  NAND2_X1 U519 ( .A1(n568), .A2(n384), .ZN(n466) );
  XOR2_X1 U520 ( .A(KEYINPUT58), .B(KEYINPUT122), .Z(n464) );
  NOR2_X1 U521 ( .A1(n577), .A2(n518), .ZN(n503) );
  NOR2_X1 U522 ( .A1(n473), .A2(n495), .ZN(n467) );
  NAND2_X1 U523 ( .A1(n468), .A2(n467), .ZN(n469) );
  XNOR2_X1 U524 ( .A(n469), .B(KEYINPUT91), .ZN(n483) );
  OR2_X1 U525 ( .A1(n531), .A2(n535), .ZN(n470) );
  XOR2_X1 U526 ( .A(KEYINPUT93), .B(n470), .Z(n471) );
  NAND2_X1 U527 ( .A1(n471), .A2(n474), .ZN(n472) );
  XNOR2_X1 U528 ( .A(KEYINPUT25), .B(n472), .ZN(n479) );
  NOR2_X1 U529 ( .A1(n474), .A2(n473), .ZN(n475) );
  XNOR2_X1 U530 ( .A(n475), .B(KEYINPUT26), .ZN(n571) );
  INV_X1 U531 ( .A(n571), .ZN(n549) );
  NOR2_X1 U532 ( .A1(n476), .A2(n549), .ZN(n477) );
  XNOR2_X1 U533 ( .A(n477), .B(KEYINPUT92), .ZN(n478) );
  NOR2_X1 U534 ( .A1(n479), .A2(n478), .ZN(n480) );
  NOR2_X1 U535 ( .A1(n481), .A2(n480), .ZN(n482) );
  NOR2_X1 U536 ( .A1(n483), .A2(n482), .ZN(n499) );
  NOR2_X1 U537 ( .A1(n501), .A2(n384), .ZN(n484) );
  XOR2_X1 U538 ( .A(KEYINPUT16), .B(n484), .Z(n485) );
  NOR2_X1 U539 ( .A1(n499), .A2(n485), .ZN(n519) );
  NAND2_X1 U540 ( .A1(n503), .A2(n519), .ZN(n496) );
  NOR2_X1 U541 ( .A1(n529), .A2(n496), .ZN(n487) );
  XNOR2_X1 U542 ( .A(KEYINPUT34), .B(KEYINPUT94), .ZN(n486) );
  XNOR2_X1 U543 ( .A(n487), .B(n486), .ZN(n488) );
  XOR2_X1 U544 ( .A(G1GAT), .B(n488), .Z(G1324GAT) );
  NOR2_X1 U545 ( .A1(n531), .A2(n496), .ZN(n490) );
  XNOR2_X1 U546 ( .A(G8GAT), .B(KEYINPUT95), .ZN(n489) );
  XNOR2_X1 U547 ( .A(n490), .B(n489), .ZN(G1325GAT) );
  NOR2_X1 U548 ( .A1(n496), .A2(n535), .ZN(n494) );
  XOR2_X1 U549 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n492) );
  XNOR2_X1 U550 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n491) );
  XNOR2_X1 U551 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U552 ( .A(n494), .B(n493), .ZN(G1326GAT) );
  INV_X1 U553 ( .A(n495), .ZN(n539) );
  NOR2_X1 U554 ( .A1(n539), .A2(n496), .ZN(n497) );
  XOR2_X1 U555 ( .A(KEYINPUT98), .B(n497), .Z(n498) );
  XNOR2_X1 U556 ( .A(G22GAT), .B(n498), .ZN(G1327GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT99), .B(KEYINPUT38), .Z(n505) );
  NOR2_X1 U558 ( .A1(n499), .A2(n588), .ZN(n500) );
  NAND2_X1 U559 ( .A1(n501), .A2(n500), .ZN(n502) );
  XNOR2_X1 U560 ( .A(KEYINPUT37), .B(n502), .ZN(n528) );
  NAND2_X1 U561 ( .A1(n503), .A2(n528), .ZN(n504) );
  XNOR2_X1 U562 ( .A(n505), .B(n504), .ZN(n513) );
  NOR2_X1 U563 ( .A1(n513), .A2(n529), .ZN(n507) );
  XNOR2_X1 U564 ( .A(KEYINPUT39), .B(KEYINPUT100), .ZN(n506) );
  XNOR2_X1 U565 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U566 ( .A(G29GAT), .B(n508), .ZN(G1328GAT) );
  NOR2_X1 U567 ( .A1(n513), .A2(n531), .ZN(n509) );
  XOR2_X1 U568 ( .A(G36GAT), .B(n509), .Z(G1329GAT) );
  XNOR2_X1 U569 ( .A(KEYINPUT40), .B(KEYINPUT101), .ZN(n511) );
  NOR2_X1 U570 ( .A1(n535), .A2(n513), .ZN(n510) );
  XNOR2_X1 U571 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U572 ( .A(G43GAT), .B(n512), .ZN(G1330GAT) );
  NOR2_X1 U573 ( .A1(n539), .A2(n513), .ZN(n514) );
  XOR2_X1 U574 ( .A(G50GAT), .B(n514), .Z(n515) );
  XNOR2_X1 U575 ( .A(KEYINPUT102), .B(n515), .ZN(G1331GAT) );
  XOR2_X1 U576 ( .A(KEYINPUT104), .B(KEYINPUT42), .Z(n517) );
  XNOR2_X1 U577 ( .A(G57GAT), .B(KEYINPUT103), .ZN(n516) );
  XNOR2_X1 U578 ( .A(n517), .B(n516), .ZN(n521) );
  AND2_X1 U579 ( .A1(n518), .A2(n563), .ZN(n527) );
  NAND2_X1 U580 ( .A1(n527), .A2(n519), .ZN(n524) );
  NOR2_X1 U581 ( .A1(n529), .A2(n524), .ZN(n520) );
  XOR2_X1 U582 ( .A(n521), .B(n520), .Z(G1332GAT) );
  NOR2_X1 U583 ( .A1(n531), .A2(n524), .ZN(n522) );
  XOR2_X1 U584 ( .A(G64GAT), .B(n522), .Z(G1333GAT) );
  NOR2_X1 U585 ( .A1(n535), .A2(n524), .ZN(n523) );
  XOR2_X1 U586 ( .A(G71GAT), .B(n523), .Z(G1334GAT) );
  NOR2_X1 U587 ( .A1(n539), .A2(n524), .ZN(n526) );
  XNOR2_X1 U588 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n525) );
  XNOR2_X1 U589 ( .A(n526), .B(n525), .ZN(G1335GAT) );
  NAND2_X1 U590 ( .A1(n528), .A2(n527), .ZN(n538) );
  NOR2_X1 U591 ( .A1(n529), .A2(n538), .ZN(n530) );
  XOR2_X1 U592 ( .A(G85GAT), .B(n530), .Z(G1336GAT) );
  NOR2_X1 U593 ( .A1(n531), .A2(n538), .ZN(n533) );
  XNOR2_X1 U594 ( .A(KEYINPUT105), .B(KEYINPUT106), .ZN(n532) );
  XNOR2_X1 U595 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U596 ( .A(G92GAT), .B(n534), .ZN(G1337GAT) );
  NOR2_X1 U597 ( .A1(n535), .A2(n538), .ZN(n537) );
  XNOR2_X1 U598 ( .A(G99GAT), .B(KEYINPUT107), .ZN(n536) );
  XNOR2_X1 U599 ( .A(n537), .B(n536), .ZN(G1338GAT) );
  NOR2_X1 U600 ( .A1(n539), .A2(n538), .ZN(n541) );
  XNOR2_X1 U601 ( .A(KEYINPUT44), .B(KEYINPUT108), .ZN(n540) );
  XNOR2_X1 U602 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U603 ( .A(G106GAT), .B(n542), .Z(G1339GAT) );
  NAND2_X1 U604 ( .A1(n546), .A2(n573), .ZN(n543) );
  XNOR2_X1 U605 ( .A(n543), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U606 ( .A(G120GAT), .B(KEYINPUT49), .Z(n545) );
  NAND2_X1 U607 ( .A1(n546), .A2(n563), .ZN(n544) );
  XNOR2_X1 U608 ( .A(n545), .B(n544), .ZN(G1341GAT) );
  XOR2_X1 U609 ( .A(G134GAT), .B(KEYINPUT51), .Z(n548) );
  NAND2_X1 U610 ( .A1(n546), .A2(n384), .ZN(n547) );
  XNOR2_X1 U611 ( .A(n548), .B(n547), .ZN(G1343GAT) );
  NOR2_X1 U612 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U613 ( .A(n551), .B(KEYINPUT112), .ZN(n560) );
  NAND2_X1 U614 ( .A1(n560), .A2(n573), .ZN(n552) );
  XNOR2_X1 U615 ( .A(n552), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT52), .B(KEYINPUT53), .Z(n554) );
  NAND2_X1 U617 ( .A1(n563), .A2(n560), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n554), .B(n553), .ZN(n556) );
  XOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT113), .Z(n555) );
  XNOR2_X1 U620 ( .A(n556), .B(n555), .ZN(G1345GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n558) );
  NAND2_X1 U622 ( .A1(n560), .A2(n582), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U624 ( .A(G155GAT), .B(n559), .ZN(G1346GAT) );
  NAND2_X1 U625 ( .A1(n560), .A2(n384), .ZN(n561) );
  XNOR2_X1 U626 ( .A(n561), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U627 ( .A1(n573), .A2(n568), .ZN(n562) );
  XNOR2_X1 U628 ( .A(G169GAT), .B(n562), .ZN(G1348GAT) );
  NAND2_X1 U629 ( .A1(n568), .A2(n563), .ZN(n565) );
  XOR2_X1 U630 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(n567) );
  XOR2_X1 U632 ( .A(G176GAT), .B(KEYINPUT56), .Z(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(G1349GAT) );
  NAND2_X1 U634 ( .A1(n582), .A2(n568), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n569), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n575) );
  NAND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n572), .B(KEYINPUT123), .ZN(n586) );
  NAND2_X1 U639 ( .A1(n586), .A2(n573), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(n576), .ZN(G1352GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n579) );
  NAND2_X1 U643 ( .A1(n586), .A2(n577), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n581) );
  XOR2_X1 U645 ( .A(G204GAT), .B(KEYINPUT124), .Z(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1353GAT) );
  NAND2_X1 U647 ( .A1(n582), .A2(n586), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n583), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U649 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n585) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n584) );
  XNOR2_X1 U651 ( .A(n585), .B(n584), .ZN(n590) );
  INV_X1 U652 ( .A(n586), .ZN(n587) );
  NOR2_X1 U653 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U654 ( .A(n590), .B(n589), .Z(G1355GAT) );
endmodule

