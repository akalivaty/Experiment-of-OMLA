//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 1 1 1 1 1 0 1 1 0 0 1 1 1 0 0 0 0 1 0 1 1 1 0 1 0 0 1 1 1 1 0 1 0 0 1 1 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:12 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(G110), .B(G140), .ZN(new_n192));
  INV_X1    g006(.A(G953), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G227), .ZN(new_n194));
  XOR2_X1   g008(.A(new_n192), .B(new_n194), .Z(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G128), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(KEYINPUT1), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G143), .ZN(new_n200));
  INV_X1    g014(.A(G143), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G146), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n198), .A2(new_n200), .A3(new_n202), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n197), .B1(new_n200), .B2(KEYINPUT1), .ZN(new_n204));
  XNOR2_X1  g018(.A(G143), .B(G146), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT10), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT75), .ZN(new_n210));
  INV_X1    g024(.A(G107), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT3), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n211), .B1(new_n212), .B2(G104), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(G104), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G104), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n216), .A2(KEYINPUT3), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n211), .A2(KEYINPUT71), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT71), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G107), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n217), .A2(new_n218), .A3(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G101), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n215), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(KEYINPUT72), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT72), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n215), .A2(new_n221), .A3(new_n225), .A4(new_n222), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(G101), .B1(new_n216), .B2(new_n211), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT71), .B(G107), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n228), .B1(new_n229), .B2(new_n216), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n210), .B1(new_n227), .B2(new_n231), .ZN(new_n232));
  AOI211_X1 g046(.A(KEYINPUT75), .B(new_n230), .C1(new_n224), .C2(new_n226), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n209), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n222), .B1(new_n215), .B2(new_n221), .ZN(new_n235));
  OR2_X1    g049(.A1(new_n235), .A2(KEYINPUT4), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n235), .B1(new_n224), .B2(new_n226), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT4), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n205), .A2(KEYINPUT0), .A3(G128), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT0), .B(G128), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n240), .B1(new_n205), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n239), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n205), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n200), .A2(KEYINPUT1), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n246), .A2(KEYINPUT74), .ZN(new_n247));
  OAI21_X1  g061(.A(G128), .B1(new_n246), .B2(KEYINPUT74), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n245), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  OR2_X1    g063(.A1(new_n203), .A2(KEYINPUT73), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n203), .A2(KEYINPUT73), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n252), .A2(new_n227), .A3(new_n231), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(new_n208), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n234), .A2(new_n244), .A3(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G131), .ZN(new_n256));
  AND2_X1   g070(.A1(KEYINPUT64), .A2(G134), .ZN(new_n257));
  NOR2_X1   g071(.A1(KEYINPUT64), .A2(G134), .ZN(new_n258));
  INV_X1    g072(.A(G137), .ZN(new_n259));
  NOR3_X1   g073(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(G134), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n261), .A2(G137), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT11), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT11), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n257), .A2(new_n258), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n264), .B1(new_n265), .B2(G137), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n256), .B1(new_n263), .B2(new_n266), .ZN(new_n267));
  OR2_X1    g081(.A1(KEYINPUT64), .A2(G134), .ZN(new_n268));
  NAND2_X1  g082(.A1(KEYINPUT64), .A2(G134), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n268), .A2(G137), .A3(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n262), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n264), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(KEYINPUT64), .B(G134), .ZN(new_n273));
  AOI21_X1  g087(.A(KEYINPUT11), .B1(new_n273), .B2(new_n259), .ZN(new_n274));
  NOR3_X1   g088(.A1(new_n272), .A2(new_n274), .A3(G131), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n267), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n255), .A2(new_n277), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n234), .A2(new_n244), .A3(new_n254), .A4(new_n276), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n196), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AND3_X1   g094(.A1(new_n252), .A2(new_n227), .A3(new_n231), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n232), .A2(new_n233), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n281), .B1(new_n282), .B2(new_n207), .ZN(new_n283));
  OAI21_X1  g097(.A(KEYINPUT12), .B1(new_n283), .B2(new_n276), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT12), .ZN(new_n285));
  NOR3_X1   g099(.A1(new_n232), .A2(new_n233), .A3(new_n206), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n285), .B(new_n277), .C1(new_n286), .C2(new_n281), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n284), .A2(new_n196), .A3(new_n279), .A4(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT76), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n280), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n227), .A2(new_n231), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT75), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n227), .A2(new_n210), .A3(new_n231), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n292), .A2(new_n293), .A3(new_n207), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(new_n253), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n285), .B1(new_n295), .B2(new_n277), .ZN(new_n296));
  AOI211_X1 g110(.A(KEYINPUT12), .B(new_n276), .C1(new_n294), .C2(new_n253), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n298), .A2(KEYINPUT76), .A3(new_n196), .A4(new_n279), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n290), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G469), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n300), .A2(new_n301), .A3(new_n190), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n301), .A2(new_n190), .ZN(new_n303));
  AND3_X1   g117(.A1(new_n278), .A2(new_n196), .A3(new_n279), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n284), .A2(new_n279), .A3(new_n287), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n304), .B1(new_n195), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n303), .B1(new_n306), .B2(G469), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n191), .B1(new_n302), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(G214), .B1(G237), .B2(G902), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G125), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n206), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n312), .B1(new_n242), .B2(new_n311), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n193), .A2(G224), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(KEYINPUT7), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n313), .B(new_n315), .ZN(new_n316));
  XNOR2_X1  g130(.A(G116), .B(G119), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT5), .ZN(new_n318));
  INV_X1    g132(.A(G116), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n319), .A2(G119), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n318), .B(G113), .C1(KEYINPUT5), .C2(new_n321), .ZN(new_n322));
  XOR2_X1   g136(.A(KEYINPUT2), .B(G113), .Z(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(new_n317), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n326), .B1(new_n232), .B2(new_n233), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n291), .A2(new_n325), .ZN(new_n328));
  AND2_X1   g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(G110), .B(G122), .ZN(new_n330));
  XOR2_X1   g144(.A(new_n330), .B(KEYINPUT8), .Z(new_n331));
  OAI211_X1 g145(.A(KEYINPUT78), .B(new_n316), .C1(new_n329), .C2(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT2), .B(G113), .ZN(new_n333));
  INV_X1    g147(.A(G119), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n334), .A2(G116), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n333), .B1(new_n320), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n324), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT65), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n337), .B(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n239), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n327), .A2(new_n340), .A3(new_n330), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT78), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n331), .B1(new_n327), .B2(new_n328), .ZN(new_n343));
  INV_X1    g157(.A(new_n316), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n332), .A2(new_n341), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n327), .A2(new_n340), .ZN(new_n347));
  INV_X1    g161(.A(new_n330), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(KEYINPUT6), .A3(new_n341), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n314), .B(KEYINPUT77), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n313), .B(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT6), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n347), .A2(new_n353), .A3(new_n348), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n350), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n346), .A2(new_n355), .A3(new_n190), .ZN(new_n356));
  OAI21_X1  g170(.A(G210), .B1(G237), .B2(G902), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n346), .A2(new_n355), .A3(new_n190), .A4(new_n357), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n310), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NOR2_X1   g175(.A1(G237), .A2(G953), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(G143), .A3(G214), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(G143), .B1(new_n362), .B2(G214), .ZN(new_n365));
  OAI21_X1  g179(.A(G131), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n365), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n367), .A2(new_n256), .A3(new_n363), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT17), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n366), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(KEYINPUT81), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT81), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n366), .A2(new_n368), .A3(new_n372), .A4(new_n369), .ZN(new_n373));
  OR2_X1    g187(.A1(new_n366), .A2(new_n369), .ZN(new_n374));
  NOR3_X1   g188(.A1(new_n311), .A2(KEYINPUT16), .A3(G140), .ZN(new_n375));
  XNOR2_X1  g189(.A(G125), .B(G140), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n375), .B1(new_n376), .B2(KEYINPUT16), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n377), .A2(G146), .ZN(new_n378));
  AOI211_X1 g192(.A(new_n199), .B(new_n375), .C1(KEYINPUT16), .C2(new_n376), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n371), .A2(new_n373), .A3(new_n374), .A4(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(G140), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G125), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n311), .A2(G140), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT69), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n376), .A2(KEYINPUT69), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(new_n388), .A3(new_n199), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n385), .A2(G146), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT18), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n367), .B(new_n363), .C1(new_n392), .C2(new_n256), .ZN(new_n393));
  OAI211_X1 g207(.A(KEYINPUT18), .B(G131), .C1(new_n364), .C2(new_n365), .ZN(new_n394));
  AND3_X1   g208(.A1(new_n391), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  XNOR2_X1  g210(.A(G113), .B(G122), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n397), .B(new_n216), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n381), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n398), .B1(new_n381), .B2(new_n396), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n190), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G475), .ZN(new_n403));
  AOI22_X1  g217(.A1(new_n366), .A2(new_n368), .B1(G146), .B2(new_n377), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT19), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n387), .A2(new_n388), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n385), .A2(KEYINPUT19), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n406), .A2(KEYINPUT79), .A3(new_n199), .A4(new_n407), .ZN(new_n408));
  AND2_X1   g222(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT79), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n406), .A2(new_n407), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n410), .B1(new_n411), .B2(G146), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n395), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(KEYINPUT80), .B1(new_n413), .B2(new_n398), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n412), .A2(new_n408), .A3(new_n404), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n396), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT80), .ZN(new_n417));
  INV_X1    g231(.A(new_n398), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n414), .A2(new_n419), .A3(new_n399), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT20), .ZN(new_n421));
  NOR2_X1   g235(.A1(G475), .A2(G902), .ZN(new_n422));
  AND3_X1   g236(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n421), .B1(new_n420), .B2(new_n422), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n403), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(KEYINPUT21), .B(G898), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n426), .B(KEYINPUT84), .ZN(new_n427));
  AOI211_X1 g241(.A(new_n190), .B(new_n193), .C1(G234), .C2(G237), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n193), .A2(G952), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n430), .B1(G234), .B2(G237), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(G478), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n435), .A2(KEYINPUT15), .ZN(new_n436));
  INV_X1    g250(.A(G217), .ZN(new_n437));
  NOR3_X1   g251(.A1(new_n188), .A2(new_n437), .A3(G953), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT82), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n439), .B1(new_n197), .B2(G143), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n201), .A2(KEYINPUT82), .A3(G128), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  AND2_X1   g256(.A1(KEYINPUT83), .A2(KEYINPUT13), .ZN(new_n443));
  NOR2_X1   g257(.A1(KEYINPUT83), .A2(KEYINPUT13), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n440), .B(new_n441), .C1(new_n444), .C2(new_n443), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n197), .A2(G143), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(G134), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n218), .A2(new_n220), .ZN(new_n451));
  INV_X1    g265(.A(G122), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(G116), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n319), .A2(G122), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n451), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g270(.A(G116), .B(G122), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n229), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  AOI22_X1  g273(.A1(new_n440), .A2(new_n441), .B1(new_n197), .B2(G143), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n265), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n450), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n452), .A2(G116), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n211), .B1(new_n463), .B2(KEYINPUT14), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT14), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n453), .A2(new_n454), .A3(new_n465), .ZN(new_n466));
  AOI22_X1  g280(.A1(new_n464), .A2(new_n466), .B1(new_n229), .B2(new_n457), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n442), .A2(new_n265), .A3(new_n448), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n265), .B1(new_n442), .B2(new_n448), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n438), .B1(new_n462), .B2(new_n470), .ZN(new_n471));
  AOI22_X1  g285(.A1(new_n442), .A2(new_n445), .B1(new_n197), .B2(G143), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n261), .B1(new_n472), .B2(new_n447), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n459), .A2(new_n461), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n470), .B(new_n438), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n436), .B1(new_n477), .B2(G902), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NOR3_X1   g293(.A1(new_n477), .A2(G902), .A3(new_n436), .ZN(new_n480));
  OR2_X1    g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NOR3_X1   g295(.A1(new_n425), .A2(new_n434), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n308), .A2(new_n361), .A3(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(G131), .B1(new_n272), .B2(new_n274), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n262), .B1(new_n265), .B2(G137), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n256), .B(new_n266), .C1(new_n485), .C2(new_n264), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n242), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(G137), .B1(new_n268), .B2(new_n269), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n259), .A2(G134), .ZN(new_n489));
  OAI21_X1  g303(.A(G131), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n206), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n275), .A2(new_n491), .ZN(new_n492));
  NOR3_X1   g306(.A1(new_n487), .A2(new_n492), .A3(KEYINPUT30), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT30), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n243), .B1(new_n267), .B2(new_n275), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n486), .A2(new_n206), .A3(new_n490), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n339), .B1(new_n493), .B2(new_n497), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n337), .B(KEYINPUT65), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n495), .A2(new_n499), .A3(new_n496), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n362), .A2(G210), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n501), .B(KEYINPUT27), .ZN(new_n502));
  XNOR2_X1  g316(.A(KEYINPUT26), .B(G101), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n502), .B(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n498), .A2(new_n500), .A3(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n504), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT28), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n339), .B1(new_n487), .B2(new_n492), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n507), .B1(new_n500), .B2(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n487), .A2(new_n492), .ZN(new_n510));
  AOI21_X1  g324(.A(KEYINPUT28), .B1(new_n510), .B2(new_n499), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n506), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT31), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n505), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(G472), .ZN(new_n515));
  NOR3_X1   g329(.A1(new_n339), .A2(new_n487), .A3(new_n492), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n495), .A2(new_n494), .A3(new_n496), .ZN(new_n517));
  OAI21_X1  g331(.A(KEYINPUT30), .B1(new_n487), .B2(new_n492), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n516), .B1(new_n519), .B2(new_n339), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(KEYINPUT31), .A3(new_n504), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n514), .A2(new_n515), .A3(new_n190), .A4(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT32), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT66), .ZN(new_n525));
  AOI211_X1 g339(.A(new_n506), .B(new_n516), .C1(new_n519), .C2(new_n339), .ZN(new_n526));
  AOI21_X1  g340(.A(G902), .B1(new_n526), .B2(KEYINPUT31), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n527), .A2(KEYINPUT32), .A3(new_n515), .A4(new_n514), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n524), .A2(new_n525), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n522), .A2(KEYINPUT66), .A3(new_n523), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NOR3_X1   g345(.A1(new_n509), .A2(new_n511), .A3(new_n506), .ZN(new_n532));
  AOI21_X1  g346(.A(G902), .B1(new_n532), .B2(KEYINPUT29), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n500), .A2(new_n508), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(KEYINPUT28), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n500), .A2(new_n507), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n535), .A2(KEYINPUT67), .A3(new_n536), .A4(new_n504), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT29), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n537), .B(new_n538), .C1(new_n504), .C2(new_n520), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n532), .A2(KEYINPUT67), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n533), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(G472), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n531), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n437), .B1(G234), .B2(new_n190), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n197), .A2(KEYINPUT23), .A3(G119), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n334), .A2(G128), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n334), .A2(G128), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n546), .B(new_n547), .C1(new_n548), .C2(KEYINPUT23), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(G110), .ZN(new_n550));
  XNOR2_X1  g364(.A(KEYINPUT24), .B(G110), .ZN(new_n551));
  OR3_X1    g365(.A1(new_n334), .A2(KEYINPUT68), .A3(G128), .ZN(new_n552));
  OAI21_X1  g366(.A(KEYINPUT68), .B1(new_n334), .B2(G128), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n552), .A2(new_n547), .A3(new_n553), .ZN(new_n554));
  OAI221_X1 g368(.A(new_n550), .B1(new_n551), .B2(new_n554), .C1(new_n378), .C2(new_n379), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n551), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n556), .B1(G110), .B2(new_n549), .ZN(new_n557));
  INV_X1    g371(.A(new_n379), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n557), .A2(new_n389), .A3(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(KEYINPUT22), .B(G137), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n193), .A2(G221), .A3(G234), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n560), .B(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n555), .A2(new_n559), .A3(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n562), .B1(new_n555), .B2(new_n559), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n566), .A2(KEYINPUT25), .A3(new_n190), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n555), .A2(new_n559), .ZN(new_n568));
  INV_X1    g382(.A(new_n562), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n570), .A2(new_n190), .A3(new_n563), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT25), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n545), .B1(new_n567), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n566), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n544), .A2(G902), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n543), .A2(KEYINPUT70), .A3(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT70), .ZN(new_n581));
  INV_X1    g395(.A(new_n540), .ZN(new_n582));
  INV_X1    g396(.A(new_n520), .ZN(new_n583));
  AOI21_X1  g397(.A(KEYINPUT29), .B1(new_n583), .B2(new_n506), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n582), .A2(new_n584), .A3(new_n537), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n515), .B1(new_n585), .B2(new_n533), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n586), .B1(new_n529), .B2(new_n530), .ZN(new_n587));
  INV_X1    g401(.A(new_n579), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n581), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n483), .B1(new_n580), .B2(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(new_n222), .ZN(G3));
  NAND2_X1  g405(.A1(new_n527), .A2(new_n514), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(G472), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n522), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n594), .A2(new_n588), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n308), .A2(new_n595), .ZN(new_n596));
  XOR2_X1   g410(.A(new_n596), .B(KEYINPUT85), .Z(new_n597));
  AND2_X1   g411(.A1(KEYINPUT86), .A2(KEYINPUT33), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n599), .B1(new_n471), .B2(new_n476), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n470), .B1(new_n473), .B2(new_n474), .ZN(new_n601));
  INV_X1    g415(.A(new_n438), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(KEYINPUT86), .A2(KEYINPUT33), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n603), .B(new_n475), .C1(new_n604), .C2(new_n598), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n435), .A2(G902), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n600), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT87), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n600), .A2(new_n605), .A3(KEYINPUT87), .A4(new_n606), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n435), .B1(new_n477), .B2(G902), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g426(.A(KEYINPUT88), .B1(new_n609), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n607), .A2(new_n608), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT88), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n614), .A2(new_n615), .A3(new_n610), .A4(new_n611), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n425), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  AND3_X1   g433(.A1(new_n361), .A2(new_n433), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n597), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT34), .B(G104), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G6));
  NAND2_X1  g437(.A1(new_n420), .A2(new_n422), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(KEYINPUT20), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT89), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n423), .A2(KEYINPUT89), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT91), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n481), .A2(new_n403), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n433), .B(KEYINPUT90), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n631), .A2(new_n632), .A3(new_n634), .A4(new_n635), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n634), .A2(new_n629), .A3(new_n628), .A4(new_n635), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(KEYINPUT91), .ZN(new_n638));
  AND3_X1   g452(.A1(new_n636), .A2(new_n361), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n597), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT35), .B(G107), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G9));
  NOR2_X1   g456(.A1(new_n569), .A2(KEYINPUT36), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n568), .B(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n645), .A2(new_n577), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n574), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(KEYINPUT92), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT92), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n649), .B1(new_n574), .B2(new_n646), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n651), .A2(new_n594), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n308), .A2(new_n652), .A3(new_n361), .A4(new_n482), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT37), .B(G110), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G12));
  AOI21_X1  g469(.A(new_n651), .B1(new_n531), .B2(new_n542), .ZN(new_n656));
  XNOR2_X1  g470(.A(KEYINPUT93), .B(G900), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n431), .B1(new_n428), .B2(new_n657), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n630), .A2(new_n633), .A3(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n656), .A2(new_n308), .A3(new_n361), .A4(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G128), .ZN(G30));
  XOR2_X1   g475(.A(new_n658), .B(KEYINPUT39), .Z(new_n662));
  NAND2_X1  g476(.A1(new_n308), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(new_n663), .B(KEYINPUT40), .Z(new_n664));
  NAND2_X1  g478(.A1(new_n359), .A2(new_n360), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT38), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n359), .A2(KEYINPUT38), .A3(new_n360), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n520), .A2(new_n506), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n190), .B1(new_n534), .B2(new_n504), .ZN(new_n671));
  OAI21_X1  g485(.A(G472), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n531), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n481), .A2(new_n309), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n625), .A2(new_n627), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n674), .B1(new_n675), .B2(new_n403), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n648), .A2(new_n650), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n669), .A2(new_n673), .A3(new_n679), .ZN(new_n680));
  OR2_X1    g494(.A1(new_n680), .A2(KEYINPUT94), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(KEYINPUT94), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n664), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G143), .ZN(G45));
  INV_X1    g498(.A(new_n658), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n617), .A2(new_n425), .A3(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n656), .A2(new_n308), .A3(new_n361), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G146), .ZN(G48));
  NAND2_X1  g503(.A1(new_n300), .A2(new_n190), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(G469), .ZN(new_n691));
  INV_X1    g505(.A(new_n191), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n691), .A2(new_n692), .A3(new_n302), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(KEYINPUT95), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n587), .A2(new_n588), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT95), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n691), .A2(new_n696), .A3(new_n692), .A4(new_n302), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n694), .A2(new_n695), .A3(new_n620), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(KEYINPUT41), .B(G113), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G15));
  NAND4_X1  g514(.A1(new_n639), .A2(new_n694), .A3(new_n695), .A4(new_n697), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G116), .ZN(G18));
  AND4_X1   g516(.A1(new_n692), .A2(new_n691), .A3(new_n302), .A4(new_n361), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n703), .A2(new_n482), .A3(new_n656), .ZN(new_n704));
  XNOR2_X1  g518(.A(KEYINPUT96), .B(G119), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G21));
  AND4_X1   g520(.A1(new_n665), .A2(new_n595), .A3(new_n635), .A4(new_n676), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n707), .A2(new_n694), .A3(new_n697), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT97), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n707), .A2(new_n694), .A3(KEYINPUT97), .A4(new_n697), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G122), .ZN(G24));
  AND3_X1   g527(.A1(new_n691), .A2(new_n692), .A3(new_n302), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n651), .A2(new_n686), .A3(new_n594), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n714), .A2(new_n361), .A3(new_n715), .ZN(new_n716));
  XOR2_X1   g530(.A(KEYINPUT98), .B(G125), .Z(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G27));
  INV_X1    g532(.A(KEYINPUT99), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n305), .A2(new_n719), .A3(new_n195), .ZN(new_n720));
  INV_X1    g534(.A(new_n304), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n719), .B1(new_n305), .B2(new_n195), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n303), .B1(new_n724), .B2(G469), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n191), .B1(new_n725), .B2(new_n302), .ZN(new_n726));
  AND3_X1   g540(.A1(new_n359), .A2(new_n309), .A3(new_n360), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n695), .A2(new_n726), .A3(new_n687), .A4(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT42), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT101), .ZN(new_n731));
  INV_X1    g545(.A(new_n723), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n732), .A2(new_n721), .A3(new_n720), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n301), .B1(new_n733), .B2(new_n190), .ZN(new_n734));
  INV_X1    g548(.A(new_n302), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n727), .B(new_n692), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n514), .A2(new_n190), .A3(new_n521), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT100), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n737), .A2(new_n738), .A3(KEYINPUT32), .A4(new_n515), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n528), .A2(KEYINPUT100), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n739), .A2(new_n542), .A3(new_n524), .A4(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n686), .A2(new_n729), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n741), .A2(new_n742), .A3(new_n579), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n731), .B1(new_n736), .B2(new_n743), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n741), .A2(new_n742), .A3(new_n579), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n745), .A2(KEYINPUT101), .A3(new_n727), .A4(new_n726), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n730), .A2(new_n744), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G131), .ZN(G33));
  NAND4_X1  g562(.A1(new_n695), .A2(new_n726), .A3(new_n659), .A4(new_n727), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT102), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n736), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n752), .A2(KEYINPUT102), .A3(new_n695), .A4(new_n659), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G134), .ZN(G36));
  NAND2_X1  g569(.A1(new_n724), .A2(KEYINPUT45), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n306), .A2(KEYINPUT45), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n757), .A2(new_n301), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(new_n303), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT46), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n735), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n303), .B1(new_n756), .B2(new_n758), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(KEYINPUT46), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n191), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT43), .ZN(new_n767));
  AND4_X1   g581(.A1(new_n767), .A2(new_n617), .A3(new_n675), .A4(new_n403), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n425), .A2(KEYINPUT103), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT103), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n675), .A2(new_n770), .A3(new_n403), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n769), .A2(new_n771), .A3(new_n617), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n768), .B1(KEYINPUT43), .B2(new_n772), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n594), .A2(new_n678), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n773), .A2(KEYINPUT44), .A3(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n727), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n773), .A2(new_n774), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT44), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n766), .A2(new_n662), .A3(new_n775), .A4(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(KEYINPUT104), .B(G137), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n780), .B(new_n781), .ZN(G39));
  INV_X1    g596(.A(new_n765), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n302), .B1(new_n764), .B2(KEYINPUT46), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n692), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n692), .B(new_n786), .C1(new_n783), .C2(new_n784), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NOR4_X1   g604(.A1(new_n543), .A2(new_n776), .A3(new_n579), .A4(new_n686), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G140), .ZN(G42));
  AND2_X1   g607(.A1(new_n691), .A2(new_n302), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(KEYINPUT49), .ZN(new_n795));
  NOR4_X1   g609(.A1(new_n669), .A2(new_n191), .A3(new_n310), .A4(new_n772), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n673), .A2(new_n588), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT54), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n701), .A2(new_n698), .A3(new_n704), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n634), .A2(new_n675), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n617), .A2(new_n425), .A3(KEYINPUT106), .ZN(new_n802));
  AOI21_X1  g616(.A(KEYINPUT106), .B1(new_n617), .B2(new_n425), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n801), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n635), .ZN(new_n805));
  AOI211_X1 g619(.A(new_n310), .B(new_n805), .C1(new_n359), .C2(new_n360), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n804), .A2(new_n308), .A3(new_n806), .A4(new_n595), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(new_n653), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n483), .ZN(new_n810));
  AOI21_X1  g624(.A(KEYINPUT70), .B1(new_n543), .B2(new_n579), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n587), .A2(new_n581), .A3(new_n588), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT107), .B1(new_n809), .B2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT107), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n590), .A2(new_n808), .A3(new_n815), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n712), .B(new_n800), .C1(new_n814), .C2(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n665), .A2(new_n647), .A3(new_n685), .A4(new_n676), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n726), .A2(new_n673), .A3(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n660), .A2(new_n688), .A3(new_n716), .A4(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(KEYINPUT109), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n308), .A2(new_n361), .A3(new_n659), .ZN(new_n823));
  AOI22_X1  g637(.A1(new_n823), .A2(new_n656), .B1(new_n703), .B2(new_n715), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT109), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n824), .A2(new_n825), .A3(new_n688), .A4(new_n820), .ZN(new_n826));
  AOI21_X1  g640(.A(KEYINPUT52), .B1(new_n822), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n481), .A2(new_n658), .ZN(new_n828));
  AND4_X1   g642(.A1(new_n403), .A2(new_n631), .A3(new_n678), .A4(new_n828), .ZN(new_n829));
  AND4_X1   g643(.A1(new_n308), .A2(new_n829), .A3(new_n543), .A4(new_n727), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n752), .A2(KEYINPUT108), .A3(new_n715), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT108), .ZN(new_n832));
  INV_X1    g646(.A(new_n715), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n832), .B1(new_n736), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n830), .B1(new_n831), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n747), .A2(new_n835), .A3(new_n754), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n817), .A2(new_n827), .A3(new_n836), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n821), .A2(KEYINPUT52), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(KEYINPUT53), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT110), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n822), .A2(new_n826), .A3(KEYINPUT52), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n837), .A2(KEYINPUT53), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n840), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  OR2_X1    g658(.A1(new_n843), .A2(new_n841), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n799), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT115), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n309), .B1(new_n667), .B2(new_n668), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n594), .A2(new_n432), .A3(new_n588), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n714), .A2(new_n848), .A3(new_n773), .A4(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT113), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n772), .A2(KEYINPUT43), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n617), .A2(new_n767), .A3(new_n675), .A4(new_n403), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n853), .A2(new_n854), .A3(new_n849), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n855), .A2(KEYINPUT113), .A3(new_n714), .A4(new_n848), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT114), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT50), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n852), .A2(new_n856), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  OR2_X1    g673(.A1(new_n850), .A2(new_n858), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(KEYINPUT50), .B1(new_n850), .B2(new_n851), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n857), .B1(new_n862), .B2(new_n856), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n847), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n862), .A2(new_n856), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(KEYINPUT114), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n866), .A2(KEYINPUT115), .A3(new_n859), .A4(new_n860), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n693), .A2(new_n776), .A3(new_n432), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n868), .A2(new_n797), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n617), .A2(new_n425), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n868), .A2(new_n652), .A3(new_n773), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n794), .A2(new_n191), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(KEYINPUT112), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n788), .A2(new_n789), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n855), .A2(new_n727), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT111), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n877), .B(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n873), .B1(new_n876), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n864), .A2(new_n867), .A3(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT51), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n741), .A2(new_n579), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n868), .A2(new_n884), .A3(new_n773), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(KEYINPUT48), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n869), .A2(new_n619), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n855), .A2(new_n703), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n430), .B(KEYINPUT116), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n886), .A2(new_n887), .A3(new_n888), .A4(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n871), .A2(KEYINPUT51), .A3(new_n872), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n788), .A2(new_n789), .A3(new_n874), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n891), .B1(new_n892), .B2(new_n879), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n866), .A2(new_n859), .A3(new_n860), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n890), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n883), .A2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT117), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n883), .A2(new_n895), .A3(KEYINPUT117), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT53), .B1(new_n837), .B2(new_n842), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n701), .A2(new_n698), .A3(new_n704), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n902), .B1(new_n710), .B2(new_n711), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n746), .A2(new_n744), .ZN(new_n904));
  AOI22_X1  g718(.A1(new_n904), .A2(new_n730), .B1(new_n753), .B2(new_n751), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n809), .A2(new_n813), .A3(KEYINPUT107), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n815), .B1(new_n590), .B2(new_n808), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n903), .A2(new_n905), .A3(new_n908), .A4(new_n835), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT53), .ZN(new_n910));
  NOR4_X1   g724(.A1(new_n909), .A2(new_n910), .A3(new_n827), .A4(new_n838), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n901), .A2(new_n911), .A3(KEYINPUT54), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n846), .A2(new_n900), .A3(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(G952), .A2(G953), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n798), .B1(new_n913), .B2(new_n914), .ZN(G75));
  NOR2_X1   g729(.A1(new_n193), .A2(G952), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n817), .A2(new_n836), .ZN(new_n918));
  INV_X1    g732(.A(new_n827), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n918), .A2(new_n842), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n910), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n837), .A2(KEYINPUT53), .A3(new_n839), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n190), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(KEYINPUT56), .B1(new_n923), .B2(G210), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n350), .A2(new_n354), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(new_n352), .ZN(new_n926));
  XNOR2_X1  g740(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n926), .B(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n917), .B1(new_n924), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(G902), .B1(new_n901), .B2(new_n911), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(KEYINPUT119), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT119), .ZN(new_n932));
  OAI211_X1 g746(.A(new_n932), .B(G902), .C1(new_n901), .C2(new_n911), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n931), .A2(new_n358), .A3(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT56), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n928), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n929), .B1(new_n934), .B2(new_n936), .ZN(G51));
  XNOR2_X1  g751(.A(new_n303), .B(KEYINPUT57), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n799), .B1(new_n921), .B2(new_n922), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n938), .B1(new_n912), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(new_n300), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n931), .A2(new_n756), .A3(new_n758), .A4(new_n933), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n916), .B1(new_n941), .B2(new_n942), .ZN(G54));
  AND2_X1   g757(.A1(KEYINPUT58), .A2(G475), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n931), .A2(new_n933), .A3(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n420), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n931), .A2(new_n420), .A3(new_n933), .A4(new_n944), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n947), .A2(new_n917), .A3(new_n948), .ZN(G60));
  NAND2_X1  g763(.A1(new_n600), .A2(new_n605), .ZN(new_n950));
  NAND2_X1  g764(.A1(G478), .A2(G902), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(KEYINPUT59), .Z(new_n952));
  NOR2_X1   g766(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n953), .B1(new_n912), .B2(new_n939), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n917), .ZN(new_n955));
  INV_X1    g769(.A(new_n952), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n956), .B1(new_n846), .B2(new_n912), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n955), .B1(new_n957), .B2(new_n950), .ZN(G63));
  NAND2_X1  g772(.A1(KEYINPUT121), .A2(KEYINPUT61), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT121), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT61), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(G217), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT120), .Z(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT60), .Z(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n966), .B1(new_n921), .B2(new_n922), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n917), .B1(new_n967), .B2(new_n566), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n965), .B1(new_n901), .B2(new_n911), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n969), .A2(new_n645), .ZN(new_n970));
  OAI211_X1 g784(.A(new_n959), .B(new_n962), .C1(new_n968), .C2(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n916), .B1(new_n969), .B2(new_n575), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n967), .A2(new_n644), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n972), .A2(new_n973), .A3(new_n960), .A4(new_n961), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n971), .A2(new_n974), .ZN(G66));
  INV_X1    g789(.A(G224), .ZN(new_n976));
  OAI21_X1  g790(.A(G953), .B1(new_n427), .B2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n817), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n977), .B1(new_n978), .B2(G953), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n925), .B1(G898), .B2(new_n193), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n979), .B(new_n980), .ZN(G69));
  AOI21_X1  g795(.A(new_n193), .B1(G227), .B2(G900), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT127), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n982), .A2(new_n983), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT125), .ZN(new_n986));
  OAI211_X1 g800(.A(new_n692), .B(new_n662), .C1(new_n783), .C2(new_n784), .ZN(new_n987));
  INV_X1    g801(.A(new_n665), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n988), .A2(new_n677), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n884), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n986), .B1(new_n987), .B2(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(new_n990), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n766), .A2(KEYINPUT125), .A3(new_n662), .A4(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  AND3_X1   g808(.A1(new_n792), .A2(new_n994), .A3(new_n905), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT124), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n779), .A2(new_n775), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n997), .A2(new_n987), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n824), .A2(new_n688), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n996), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(new_n999), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n780), .A2(KEYINPUT124), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(G953), .B1(new_n995), .B2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n193), .A2(G900), .ZN(new_n1005));
  OAI21_X1  g819(.A(KEYINPUT126), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT126), .ZN(new_n1007));
  INV_X1    g821(.A(new_n1005), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n792), .A2(new_n994), .A3(new_n905), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1009), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1010));
  OAI211_X1 g824(.A(new_n1007), .B(new_n1008), .C1(new_n1010), .C2(G953), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n411), .B(KEYINPUT122), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n519), .B(new_n1012), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1006), .A2(new_n1011), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n804), .A2(new_n727), .ZN(new_n1015));
  AOI211_X1 g829(.A(new_n663), .B(new_n1015), .C1(new_n580), .C2(new_n589), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n998), .A2(new_n1016), .ZN(new_n1017));
  AND3_X1   g831(.A1(new_n683), .A2(KEYINPUT62), .A3(new_n1001), .ZN(new_n1018));
  AOI21_X1  g832(.A(KEYINPUT62), .B1(new_n683), .B2(new_n1001), .ZN(new_n1019));
  OAI211_X1 g833(.A(new_n792), .B(new_n1017), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1020), .A2(new_n193), .ZN(new_n1021));
  XOR2_X1   g835(.A(new_n1013), .B(KEYINPUT123), .Z(new_n1022));
  NAND2_X1  g836(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  AOI211_X1 g837(.A(new_n984), .B(new_n985), .C1(new_n1014), .C2(new_n1023), .ZN(new_n1024));
  AND4_X1   g838(.A1(new_n983), .A2(new_n1014), .A3(new_n982), .A4(new_n1023), .ZN(new_n1025));
  NOR2_X1   g839(.A1(new_n1024), .A2(new_n1025), .ZN(G72));
  NAND2_X1  g840(.A1(G472), .A2(G902), .ZN(new_n1027));
  XOR2_X1   g841(.A(new_n1027), .B(KEYINPUT63), .Z(new_n1028));
  OAI21_X1  g842(.A(new_n1028), .B1(new_n1020), .B2(new_n817), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1029), .A2(new_n670), .ZN(new_n1030));
  INV_X1    g844(.A(new_n1028), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1031), .B1(new_n1010), .B2(new_n978), .ZN(new_n1032));
  NOR2_X1   g846(.A1(new_n583), .A2(new_n504), .ZN(new_n1033));
  INV_X1    g847(.A(new_n1033), .ZN(new_n1034));
  OAI211_X1 g848(.A(new_n1030), .B(new_n917), .C1(new_n1032), .C2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n844), .A2(new_n845), .ZN(new_n1036));
  NOR3_X1   g850(.A1(new_n1033), .A2(new_n670), .A3(new_n1031), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n1035), .B1(new_n1036), .B2(new_n1037), .ZN(G57));
endmodule


