//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 1 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 1 0 1 1 0 0 0 1 0 0 1 1 1 1 1 0 0 0 1 1 0 0 0 0 1 1 1 1 0 0 0 0 0 0 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n797, new_n798, new_n799,
    new_n801, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n973, new_n974, new_n975, new_n976,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1014,
    new_n1015;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G64gat), .B(G92gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n202), .B(new_n203), .Z(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT65), .B(KEYINPUT25), .ZN(new_n206));
  AND3_X1   g005(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n207));
  AOI21_X1  g006(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209));
  NOR3_X1   g008(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  AND2_X1   g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211));
  INV_X1    g010(.A(G169gat), .ZN(new_n212));
  INV_X1    g011(.A(G176gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT23), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n211), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n215), .A2(G176gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n212), .A2(KEYINPUT66), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT66), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(G169gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n217), .A2(new_n218), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n216), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT67), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n210), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n216), .A2(new_n221), .A3(KEYINPUT67), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n206), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT68), .ZN(new_n227));
  NAND2_X1  g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228));
  AOI22_X1  g027(.A1(new_n217), .A2(new_n212), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n214), .A2(new_n215), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n211), .A2(KEYINPUT68), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n229), .A2(KEYINPUT25), .A3(new_n230), .A4(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(G183gat), .A2(G190gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT69), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT24), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(KEYINPUT69), .A2(G183gat), .A3(G190gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT70), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT70), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n235), .A2(new_n239), .A3(new_n236), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  AND2_X1   g040(.A1(KEYINPUT71), .A2(G190gat), .ZN(new_n242));
  NOR2_X1   g041(.A1(KEYINPUT71), .A2(G190gat), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(G183gat), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n207), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n232), .B1(new_n241), .B2(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(KEYINPUT72), .B1(new_n226), .B2(new_n247), .ZN(new_n248));
  AND3_X1   g047(.A1(new_n235), .A2(new_n239), .A3(new_n236), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n239), .B1(new_n235), .B2(new_n236), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n246), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n232), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT72), .ZN(new_n254));
  AND3_X1   g053(.A1(new_n216), .A2(new_n221), .A3(KEYINPUT67), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT67), .B1(new_n216), .B2(new_n221), .ZN(new_n256));
  NOR3_X1   g055(.A1(new_n255), .A2(new_n256), .A3(new_n210), .ZN(new_n257));
  OAI211_X1 g056(.A(new_n253), .B(new_n254), .C1(new_n257), .C2(new_n206), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT74), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT26), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n259), .A2(new_n260), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n261), .B1(new_n262), .B2(new_n214), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n259), .A2(new_n260), .A3(new_n212), .A4(new_n213), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n263), .A2(new_n228), .A3(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT27), .B(G183gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n244), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(KEYINPUT28), .ZN(new_n268));
  OR3_X1    g067(.A1(new_n245), .A2(KEYINPUT73), .A3(KEYINPUT27), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT28), .ZN(new_n270));
  OAI21_X1  g069(.A(KEYINPUT27), .B1(new_n245), .B2(KEYINPUT73), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n269), .A2(new_n244), .A3(new_n270), .A4(new_n271), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n265), .A2(new_n268), .A3(new_n233), .A4(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT75), .ZN(new_n274));
  AOI22_X1  g073(.A1(new_n267), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT75), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n275), .A2(new_n276), .A3(new_n265), .A4(new_n272), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n248), .A2(new_n258), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(G226gat), .A2(G233gat), .ZN(new_n280));
  XOR2_X1   g079(.A(new_n280), .B(KEYINPUT81), .Z(new_n281));
  NAND2_X1  g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n281), .ZN(new_n283));
  INV_X1    g082(.A(new_n273), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n222), .A2(new_n223), .ZN(new_n285));
  INV_X1    g084(.A(new_n210), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(new_n225), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n206), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n284), .B1(new_n289), .B2(new_n253), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n283), .B1(new_n290), .B2(KEYINPUT29), .ZN(new_n291));
  NAND2_X1  g090(.A1(G211gat), .A2(G218gat), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT22), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AND2_X1   g093(.A1(KEYINPUT79), .A2(G197gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(KEYINPUT79), .A2(G197gat), .ZN(new_n296));
  INV_X1    g095(.A(G204gat), .ZN(new_n297));
  NOR3_X1   g096(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT79), .ZN(new_n299));
  INV_X1    g098(.A(G197gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(KEYINPUT79), .A2(G197gat), .ZN(new_n302));
  AOI21_X1  g101(.A(G204gat), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n294), .B1(new_n298), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(G211gat), .ZN(new_n305));
  INV_X1    g104(.A(G218gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT80), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n307), .A2(new_n308), .A3(new_n292), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n304), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n297), .B1(new_n295), .B2(new_n296), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n301), .A2(G204gat), .A3(new_n302), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n314), .A2(new_n309), .A3(new_n294), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  AND3_X1   g115(.A1(new_n282), .A2(new_n291), .A3(new_n316), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n281), .A2(KEYINPUT29), .ZN(new_n318));
  AOI221_X4 g117(.A(new_n316), .B1(new_n290), .B2(new_n281), .C1(new_n279), .C2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n205), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n282), .A2(new_n291), .A3(new_n316), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n279), .A2(new_n318), .ZN(new_n322));
  AND3_X1   g121(.A1(new_n314), .A2(new_n309), .A3(new_n294), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n309), .B1(new_n314), .B2(new_n294), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n290), .A2(new_n281), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n322), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n321), .A2(new_n327), .A3(new_n204), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n320), .A2(KEYINPUT30), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n321), .A2(new_n327), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT30), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n331), .A2(new_n332), .A3(new_n204), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT78), .ZN(new_n334));
  AND2_X1   g133(.A1(G113gat), .A2(G120gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(G113gat), .A2(G120gat), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n334), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(G113gat), .ZN(new_n338));
  INV_X1    g137(.A(G120gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(G113gat), .A2(G120gat), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n340), .A2(KEYINPUT78), .A3(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT1), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n337), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(KEYINPUT76), .B(G134gat), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT77), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(new_n346), .A3(G127gat), .ZN(new_n347));
  INV_X1    g146(.A(G134gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT76), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT76), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(G134gat), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n349), .A2(new_n351), .A3(G127gat), .ZN(new_n352));
  INV_X1    g151(.A(G127gat), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n346), .B1(new_n353), .B2(G134gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n344), .A2(new_n347), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(KEYINPUT1), .B1(new_n353), .B2(G134gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n348), .A2(G127gat), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n357), .A2(new_n340), .A3(new_n341), .A4(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  AND2_X1   g159(.A1(G155gat), .A2(G162gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(G155gat), .A2(G162gat), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(G141gat), .B(G148gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(KEYINPUT82), .B(KEYINPUT2), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(G141gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(G148gat), .ZN(new_n368));
  INV_X1    g167(.A(G148gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(G141gat), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n368), .A2(new_n370), .A3(KEYINPUT83), .ZN(new_n371));
  OR3_X1    g170(.A1(new_n369), .A2(KEYINPUT83), .A3(G141gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(G155gat), .B(G162gat), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(G155gat), .A2(G162gat), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT84), .ZN(new_n376));
  AND3_X1   g175(.A1(new_n375), .A2(new_n376), .A3(KEYINPUT2), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n376), .B1(new_n375), .B2(KEYINPUT2), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n366), .B1(new_n374), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n360), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT86), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT2), .ZN(new_n383));
  OAI21_X1  g182(.A(KEYINPUT84), .B1(new_n361), .B2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n375), .A2(new_n376), .A3(KEYINPUT2), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n386), .A2(new_n371), .A3(new_n373), .A4(new_n372), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n356), .A2(new_n387), .A3(new_n366), .A4(new_n359), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n381), .A2(new_n382), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(G225gat), .A2(G233gat), .ZN(new_n390));
  XOR2_X1   g189(.A(new_n390), .B(KEYINPUT85), .Z(new_n391));
  NAND3_X1  g190(.A1(new_n360), .A2(KEYINPUT86), .A3(new_n380), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n389), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT4), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n388), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT3), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT3), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n366), .B(new_n397), .C1(new_n374), .C2(new_n379), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n396), .A2(new_n360), .A3(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n380), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n400), .A2(KEYINPUT4), .A3(new_n356), .A4(new_n359), .ZN(new_n401));
  INV_X1    g200(.A(new_n391), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n395), .A2(new_n399), .A3(new_n401), .A4(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n393), .A2(KEYINPUT5), .A3(new_n403), .ZN(new_n404));
  AND2_X1   g203(.A1(new_n395), .A2(new_n401), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT5), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n405), .A2(new_n406), .A3(new_n402), .A4(new_n399), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(G1gat), .B(G29gat), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT0), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(G57gat), .B(G85gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n411), .B(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n408), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT6), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n393), .A2(KEYINPUT5), .A3(new_n403), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n413), .B1(new_n403), .B2(KEYINPUT5), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n415), .B(new_n416), .C1(new_n417), .C2(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n408), .A2(KEYINPUT6), .A3(new_n414), .ZN(new_n420));
  AOI22_X1  g219(.A1(new_n329), .A2(new_n333), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  XNOR2_X1  g220(.A(KEYINPUT31), .B(G50gat), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(G228gat), .A2(G233gat), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT29), .B1(new_n311), .B2(new_n315), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n380), .B1(new_n426), .B2(KEYINPUT3), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT29), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n398), .A2(new_n428), .ZN(new_n429));
  AND3_X1   g228(.A1(new_n325), .A2(new_n429), .A3(KEYINPUT88), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT88), .B1(new_n325), .B2(new_n429), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n425), .B(new_n427), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(G22gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n424), .B(KEYINPUT87), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n316), .B1(new_n428), .B2(new_n398), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n307), .A2(new_n292), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n304), .A2(new_n436), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n314), .A2(KEYINPUT22), .A3(new_n292), .A4(new_n307), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n437), .A2(new_n428), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n400), .B1(new_n439), .B2(new_n397), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n434), .B1(new_n435), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n432), .A2(new_n433), .A3(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n433), .B1(new_n432), .B2(new_n441), .ZN(new_n444));
  XNOR2_X1  g243(.A(G78gat), .B(G106gat), .ZN(new_n445));
  NOR3_X1   g244(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n445), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n432), .A2(new_n441), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(G22gat), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n447), .B1(new_n449), .B2(new_n442), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n423), .B1(new_n446), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n445), .B1(new_n443), .B2(new_n444), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n449), .A2(new_n442), .A3(new_n447), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n452), .A2(new_n453), .A3(new_n422), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n360), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n279), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n248), .A2(new_n258), .A3(new_n278), .A4(new_n360), .ZN(new_n458));
  NAND2_X1  g257(.A1(G227gat), .A2(G233gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n459), .B(KEYINPUT64), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n457), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT32), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT33), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  XOR2_X1   g263(.A(G15gat), .B(G43gat), .Z(new_n465));
  XNOR2_X1  g264(.A(G71gat), .B(G99gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n465), .B(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n462), .A2(new_n464), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n457), .A2(new_n458), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n460), .A2(KEYINPUT34), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n459), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT34), .ZN(new_n473));
  INV_X1    g272(.A(new_n467), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n461), .B(KEYINPUT32), .C1(new_n463), .C2(new_n474), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n468), .A2(new_n471), .A3(new_n473), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n468), .A2(new_n475), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n473), .A2(new_n471), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n421), .A2(new_n455), .A3(new_n476), .A4(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT35), .ZN(new_n481));
  INV_X1    g280(.A(new_n476), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n468), .A2(new_n475), .B1(new_n471), .B2(new_n473), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n329), .A2(new_n333), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n416), .B1(new_n417), .B2(new_n418), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n413), .B(KEYINPUT89), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n487), .B1(new_n404), .B2(new_n407), .ZN(new_n488));
  OR2_X1    g287(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(KEYINPUT35), .B1(new_n489), .B2(new_n420), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n484), .A2(new_n485), .A3(new_n455), .A4(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n481), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT36), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n493), .B1(new_n482), .B2(new_n483), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n479), .A2(KEYINPUT36), .A3(new_n476), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(KEYINPUT93), .B(KEYINPUT37), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n205), .B1(new_n330), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT37), .ZN(new_n501));
  AOI22_X1  g300(.A1(new_n279), .A2(new_n318), .B1(new_n281), .B2(new_n290), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n501), .B1(new_n502), .B2(new_n316), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n282), .A2(new_n291), .A3(new_n325), .ZN(new_n504));
  AOI21_X1  g303(.A(KEYINPUT38), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n500), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n501), .B1(new_n321), .B2(new_n327), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT38), .B1(new_n499), .B2(new_n507), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n420), .B(new_n328), .C1(new_n486), .C2(new_n488), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n506), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n395), .A2(new_n399), .A3(new_n401), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(new_n391), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n391), .B1(new_n389), .B2(new_n392), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT39), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n514), .B1(new_n517), .B2(KEYINPUT91), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT91), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n519), .B1(new_n515), .B2(new_n516), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n512), .A2(new_n516), .A3(new_n391), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(new_n487), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT90), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n521), .A2(KEYINPUT90), .A3(new_n487), .ZN(new_n525));
  AOI22_X1  g324(.A1(new_n518), .A2(new_n520), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g325(.A1(KEYINPUT92), .A2(KEYINPUT40), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n488), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n517), .A2(KEYINPUT91), .ZN(new_n530));
  AND3_X1   g329(.A1(new_n530), .A2(new_n520), .A3(new_n513), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n524), .A2(new_n525), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n527), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n529), .A2(new_n533), .A3(new_n333), .A4(new_n329), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n511), .A2(new_n534), .A3(new_n455), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n421), .A2(new_n455), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n496), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n492), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT104), .ZN(new_n540));
  XOR2_X1   g339(.A(G57gat), .B(G64gat), .Z(new_n541));
  INV_X1    g340(.A(KEYINPUT9), .ZN(new_n542));
  INV_X1    g341(.A(G71gat), .ZN(new_n543));
  INV_X1    g342(.A(G78gat), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n541), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(G71gat), .B(G78gat), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n541), .A2(new_n547), .A3(new_n545), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT21), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(G231gat), .A2(G233gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(G127gat), .B(G155gat), .Z(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(KEYINPUT20), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n555), .B(new_n557), .ZN(new_n558));
  XOR2_X1   g357(.A(G183gat), .B(G211gat), .Z(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  OR2_X1    g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n558), .A2(new_n560), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT101), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n551), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n549), .A2(KEYINPUT101), .A3(new_n550), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT21), .ZN(new_n568));
  INV_X1    g367(.A(G1gat), .ZN(new_n569));
  XOR2_X1   g368(.A(G15gat), .B(G22gat), .Z(new_n570));
  INV_X1    g369(.A(KEYINPUT97), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(G15gat), .B(G22gat), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n573), .A2(KEYINPUT97), .A3(G1gat), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n572), .B(new_n574), .C1(KEYINPUT16), .C2(new_n570), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT98), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n576), .B1(new_n573), .B2(G1gat), .ZN(new_n577));
  INV_X1    g376(.A(G8gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n575), .B(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n568), .A2(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(KEYINPUT100), .B(KEYINPUT19), .Z(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n563), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n561), .A2(new_n584), .A3(new_n562), .ZN(new_n587));
  AND2_X1   g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g387(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT95), .ZN(new_n591));
  OR2_X1    g390(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n591), .B1(new_n592), .B2(G36gat), .ZN(new_n593));
  NOR3_X1   g392(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(KEYINPUT95), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n590), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G43gat), .B(G50gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(KEYINPUT15), .ZN(new_n599));
  NAND2_X1  g398(.A1(G29gat), .A2(G36gat), .ZN(new_n600));
  AND2_X1   g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(G43gat), .B(G50gat), .Z(new_n602));
  INV_X1    g401(.A(KEYINPUT15), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n597), .A2(KEYINPUT96), .A3(new_n601), .A4(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT96), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n604), .A2(new_n600), .A3(new_n599), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n606), .B1(new_n607), .B2(new_n596), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n599), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n600), .B1(new_n590), .B2(new_n594), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT17), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI22_X1  g414(.A1(new_n605), .A2(new_n608), .B1(new_n611), .B2(new_n610), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(KEYINPUT17), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT8), .ZN(new_n618));
  NAND2_X1  g417(.A1(G99gat), .A2(G106gat), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n618), .B1(new_n619), .B2(KEYINPUT103), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n620), .B1(KEYINPUT103), .B2(new_n619), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT7), .ZN(new_n622));
  INV_X1    g421(.A(G85gat), .ZN(new_n623));
  NOR3_X1   g422(.A1(new_n622), .A2(new_n623), .A3(G92gat), .ZN(new_n624));
  OAI21_X1  g423(.A(G92gat), .B1(KEYINPUT7), .B2(G85gat), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n625), .B1(KEYINPUT7), .B2(G85gat), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n621), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(G99gat), .B(G106gat), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  OAI211_X1 g429(.A(new_n621), .B(new_n628), .C1(new_n624), .C2(new_n626), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n615), .A2(new_n617), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(G232gat), .A2(G233gat), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n634), .B(KEYINPUT102), .Z(new_n635));
  INV_X1    g434(.A(KEYINPUT41), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n632), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n637), .B1(new_n613), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n633), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g439(.A(G190gat), .B(G218gat), .Z(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n635), .A2(new_n636), .ZN(new_n643));
  XOR2_X1   g442(.A(G134gat), .B(G162gat), .Z(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n641), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n633), .A2(new_n646), .A3(new_n639), .ZN(new_n647));
  AND3_X1   g446(.A1(new_n642), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n645), .B1(new_n642), .B2(new_n647), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n540), .B1(new_n588), .B2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n650), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n586), .A2(new_n587), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n652), .A2(new_n653), .A3(KEYINPUT104), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT108), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n549), .A2(new_n550), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n628), .A2(KEYINPUT105), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n656), .A2(new_n631), .A3(new_n630), .A4(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n549), .A2(new_n550), .A3(new_n657), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n632), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT10), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n658), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n567), .A2(KEYINPUT10), .A3(new_n638), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(G230gat), .A2(G233gat), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n665), .B(KEYINPUT106), .Z(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n658), .A2(new_n660), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(new_n666), .ZN(new_n670));
  XNOR2_X1  g469(.A(G120gat), .B(G148gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT107), .ZN(new_n672));
  XNOR2_X1  g471(.A(G176gat), .B(G204gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n668), .A2(new_n670), .A3(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n674), .B1(new_n668), .B2(new_n670), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n655), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n677), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n679), .A2(KEYINPUT108), .A3(new_n675), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n651), .A2(new_n654), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n575), .B(new_n579), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n684), .B1(new_n613), .B2(new_n614), .ZN(new_n685));
  AOI22_X1  g484(.A1(new_n685), .A2(new_n617), .B1(new_n613), .B2(new_n684), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT99), .ZN(new_n687));
  NAND2_X1  g486(.A1(G229gat), .A2(G233gat), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n686), .A2(new_n687), .A3(KEYINPUT18), .A4(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n613), .A2(new_n684), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n581), .B1(new_n616), .B2(KEYINPUT17), .ZN(new_n691));
  AND3_X1   g490(.A1(new_n609), .A2(KEYINPUT17), .A3(new_n612), .ZN(new_n692));
  OAI211_X1 g491(.A(new_n688), .B(new_n690), .C1(new_n691), .C2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT18), .ZN(new_n694));
  OAI21_X1  g493(.A(KEYINPUT99), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n689), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(G113gat), .B(G141gat), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(new_n300), .ZN(new_n698));
  XNOR2_X1  g497(.A(KEYINPUT11), .B(G169gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(KEYINPUT94), .B(KEYINPUT12), .ZN(new_n701));
  XOR2_X1   g500(.A(new_n700), .B(new_n701), .Z(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n581), .A2(new_n616), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n690), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n688), .B(KEYINPUT13), .Z(new_n706));
  AOI22_X1  g505(.A1(new_n693), .A2(new_n694), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  AND3_X1   g506(.A1(new_n696), .A2(new_n703), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n703), .B1(new_n696), .B2(new_n707), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n683), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n539), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n419), .A2(new_n420), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(KEYINPUT109), .B(G1gat), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(G1324gat));
  INV_X1    g515(.A(new_n712), .ZN(new_n717));
  INV_X1    g516(.A(new_n485), .ZN(new_n718));
  XOR2_X1   g517(.A(KEYINPUT16), .B(G8gat), .Z(new_n719));
  NAND3_X1  g518(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT110), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n720), .A2(new_n721), .A3(KEYINPUT42), .ZN(new_n722));
  AOI21_X1  g521(.A(KEYINPUT42), .B1(new_n720), .B2(new_n721), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT111), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n717), .A2(new_n718), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n724), .B1(new_n725), .B2(G8gat), .ZN(new_n726));
  AOI211_X1 g525(.A(KEYINPUT111), .B(new_n578), .C1(new_n717), .C2(new_n718), .ZN(new_n727));
  OAI22_X1  g526(.A1(new_n722), .A2(new_n723), .B1(new_n726), .B2(new_n727), .ZN(G1325gat));
  INV_X1    g527(.A(new_n484), .ZN(new_n729));
  OR3_X1    g528(.A1(new_n712), .A2(G15gat), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(G15gat), .B1(new_n712), .B2(new_n496), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(G1326gat));
  NOR2_X1   g531(.A1(new_n712), .A2(new_n455), .ZN(new_n733));
  XOR2_X1   g532(.A(KEYINPUT43), .B(G22gat), .Z(new_n734));
  XNOR2_X1  g533(.A(new_n733), .B(new_n734), .ZN(G1327gat));
  AOI21_X1  g534(.A(new_n652), .B1(new_n492), .B2(new_n538), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n710), .A2(new_n653), .A3(new_n681), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  OR2_X1    g537(.A1(new_n713), .A2(G29gat), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(KEYINPUT112), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT112), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n738), .A2(new_n743), .A3(new_n740), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT45), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT44), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n509), .B1(new_n500), .B2(new_n505), .ZN(new_n749));
  AOI22_X1  g548(.A1(new_n749), .A2(new_n508), .B1(new_n454), .B2(new_n451), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n536), .B1(new_n750), .B2(new_n534), .ZN(new_n751));
  AOI22_X1  g550(.A1(new_n751), .A2(new_n496), .B1(new_n481), .B2(new_n491), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n748), .B1(new_n752), .B2(new_n652), .ZN(new_n753));
  AND3_X1   g552(.A1(new_n496), .A2(new_n535), .A3(new_n537), .ZN(new_n754));
  AND4_X1   g553(.A1(new_n476), .A2(new_n455), .A3(new_n479), .A4(new_n485), .ZN(new_n755));
  AOI22_X1  g554(.A1(new_n755), .A2(new_n490), .B1(new_n480), .B2(KEYINPUT35), .ZN(new_n756));
  OAI211_X1 g555(.A(KEYINPUT44), .B(new_n650), .C1(new_n754), .C2(new_n756), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n737), .ZN(new_n759));
  OAI21_X1  g558(.A(G29gat), .B1(new_n759), .B2(new_n713), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n742), .A2(KEYINPUT45), .A3(new_n744), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n747), .A2(new_n760), .A3(new_n761), .ZN(G1328gat));
  INV_X1    g561(.A(G36gat), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n738), .A2(new_n763), .A3(new_n718), .ZN(new_n764));
  XOR2_X1   g563(.A(new_n764), .B(KEYINPUT46), .Z(new_n765));
  OAI21_X1  g564(.A(G36gat), .B1(new_n759), .B2(new_n485), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(G1329gat));
  INV_X1    g566(.A(new_n496), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n753), .A2(new_n768), .A3(new_n737), .A4(new_n757), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(G43gat), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n729), .A2(G43gat), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n736), .A2(new_n737), .A3(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT47), .B1(new_n774), .B2(KEYINPUT113), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n772), .B1(new_n769), .B2(G43gat), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT113), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT47), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n775), .A2(new_n779), .ZN(G1330gat));
  INV_X1    g579(.A(new_n455), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n781), .A2(G50gat), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n753), .A2(new_n737), .A3(new_n757), .A4(new_n782), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n738), .A2(new_n781), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n783), .B1(new_n784), .B2(G50gat), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(KEYINPUT48), .ZN(G1331gat));
  AND4_X1   g585(.A1(new_n710), .A2(new_n651), .A3(new_n654), .A4(new_n681), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n539), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n788), .A2(new_n713), .ZN(new_n789));
  XOR2_X1   g588(.A(KEYINPUT114), .B(G57gat), .Z(new_n790));
  XNOR2_X1  g589(.A(new_n789), .B(new_n790), .ZN(G1332gat));
  NOR2_X1   g590(.A1(new_n788), .A2(new_n485), .ZN(new_n792));
  NOR2_X1   g591(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n793));
  AND2_X1   g592(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n792), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n795), .B1(new_n792), .B2(new_n793), .ZN(G1333gat));
  OAI21_X1  g595(.A(G71gat), .B1(new_n788), .B2(new_n496), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n484), .A2(new_n543), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n797), .B1(new_n788), .B2(new_n798), .ZN(new_n799));
  XOR2_X1   g598(.A(new_n799), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g599(.A1(new_n788), .A2(new_n455), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(new_n544), .ZN(G1335gat));
  NOR3_X1   g601(.A1(new_n682), .A2(G85gat), .A3(new_n713), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n696), .A2(new_n707), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n702), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n696), .A2(new_n703), .A3(new_n707), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n807), .A2(new_n653), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n809), .B1(new_n736), .B2(KEYINPUT115), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n811), .B1(new_n752), .B2(new_n652), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n810), .A2(KEYINPUT51), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(KEYINPUT51), .B1(new_n810), .B2(new_n812), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n803), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(new_n713), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n809), .A2(new_n682), .ZN(new_n817));
  AND3_X1   g616(.A1(new_n758), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n815), .B1(new_n818), .B2(new_n623), .ZN(G1336gat));
  NOR3_X1   g618(.A1(new_n682), .A2(new_n485), .A3(G92gat), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT51), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n539), .A2(KEYINPUT115), .A3(new_n650), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(new_n808), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n736), .A2(KEYINPUT115), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n822), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n810), .A2(KEYINPUT51), .A3(new_n812), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n821), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n753), .A2(new_n718), .A3(new_n757), .A4(new_n817), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(G92gat), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(KEYINPUT52), .B1(new_n828), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n820), .B1(new_n813), .B2(new_n814), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT52), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n833), .A2(new_n834), .A3(new_n830), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n832), .A2(new_n835), .ZN(G1337gat));
  XOR2_X1   g635(.A(KEYINPUT117), .B(G99gat), .Z(new_n837));
  NOR3_X1   g636(.A1(new_n729), .A2(new_n682), .A3(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n838), .B1(new_n813), .B2(new_n814), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n753), .A2(new_n768), .A3(new_n757), .A4(new_n817), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(KEYINPUT116), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n837), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n840), .A2(KEYINPUT116), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n839), .B1(new_n842), .B2(new_n843), .ZN(G1338gat));
  NOR3_X1   g643(.A1(new_n455), .A2(new_n682), .A3(G106gat), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n846), .B1(new_n826), .B2(new_n827), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n753), .A2(new_n781), .A3(new_n757), .A4(new_n817), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(G106gat), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(KEYINPUT53), .B1(new_n847), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n845), .B1(new_n813), .B2(new_n814), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT53), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n852), .A2(new_n853), .A3(new_n849), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n851), .A2(new_n854), .ZN(G1339gat));
  NAND4_X1  g654(.A1(new_n651), .A2(new_n710), .A3(new_n654), .A4(new_n682), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n686), .A2(new_n688), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n705), .A2(new_n706), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n700), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n650), .A2(new_n806), .A3(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT118), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n662), .A2(new_n663), .A3(new_n666), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n668), .A2(KEYINPUT54), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n666), .B1(new_n662), .B2(new_n663), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n674), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n863), .A2(KEYINPUT55), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n675), .ZN(new_n868));
  AOI21_X1  g667(.A(KEYINPUT55), .B1(new_n863), .B2(new_n866), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n861), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n863), .A2(new_n866), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT55), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n873), .A2(KEYINPUT118), .A3(new_n675), .A4(new_n867), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n860), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n681), .A2(new_n806), .A3(new_n859), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n877), .B1(new_n710), .B2(new_n875), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n876), .B1(new_n878), .B2(new_n652), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n856), .B1(new_n879), .B2(new_n653), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n880), .A2(new_n816), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(new_n755), .A3(new_n807), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(new_n338), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n882), .A2(new_n338), .ZN(new_n885));
  OAI21_X1  g684(.A(KEYINPUT119), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(new_n885), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT119), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n887), .A2(new_n883), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n886), .A2(new_n889), .ZN(G1340gat));
  NAND2_X1  g689(.A1(new_n881), .A2(new_n755), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n891), .A2(new_n682), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n892), .B(new_n339), .ZN(G1341gat));
  NOR2_X1   g692(.A1(new_n891), .A2(new_n588), .ZN(new_n894));
  NOR2_X1   g693(.A1(KEYINPUT120), .A2(G127gat), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n894), .B(new_n895), .ZN(G1342gat));
  NOR2_X1   g695(.A1(new_n729), .A2(new_n781), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n718), .A2(new_n652), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n881), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(G134gat), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n881), .A2(new_n345), .A3(new_n897), .A4(new_n898), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT121), .ZN(new_n902));
  AND3_X1   g701(.A1(new_n901), .A2(new_n902), .A3(KEYINPUT56), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n902), .B1(new_n901), .B2(KEYINPUT56), .ZN(new_n904));
  OAI221_X1 g703(.A(new_n900), .B1(KEYINPUT56), .B2(new_n901), .C1(new_n903), .C2(new_n904), .ZN(G1343gat));
  NOR3_X1   g704(.A1(new_n768), .A2(new_n713), .A3(new_n718), .ZN(new_n906));
  AOI21_X1  g705(.A(KEYINPUT57), .B1(new_n880), .B2(new_n781), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT57), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n455), .A2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n873), .A2(new_n675), .A3(new_n867), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n911), .B1(new_n805), .B2(new_n806), .ZN(new_n912));
  AND3_X1   g711(.A1(new_n681), .A2(new_n806), .A3(new_n859), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n652), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n588), .B1(new_n915), .B2(new_n876), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n910), .B1(new_n916), .B2(new_n856), .ZN(new_n917));
  OAI211_X1 g716(.A(new_n807), .B(new_n906), .C1(new_n907), .C2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(G141gat), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT58), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n768), .A2(new_n713), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n880), .A2(new_n781), .A3(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT122), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n710), .A2(G141gat), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n880), .A2(KEYINPUT122), .A3(new_n781), .A4(new_n921), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n924), .A2(new_n485), .A3(new_n925), .A4(new_n926), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n919), .A2(new_n920), .A3(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(new_n922), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n710), .A2(new_n718), .A3(G141gat), .ZN(new_n930));
  AOI22_X1  g729(.A1(new_n918), .A2(G141gat), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n928), .B1(new_n931), .B2(new_n920), .ZN(G1344gat));
  NAND2_X1  g731(.A1(new_n906), .A2(new_n681), .ZN(new_n933));
  INV_X1    g732(.A(new_n856), .ZN(new_n934));
  OR2_X1    g733(.A1(new_n860), .A2(new_n911), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n653), .B1(new_n914), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n781), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(new_n908), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n880), .A2(new_n909), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n933), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g739(.A(KEYINPUT59), .B1(new_n940), .B2(new_n369), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n369), .A2(KEYINPUT59), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n906), .B1(new_n907), .B2(new_n917), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n942), .B1(new_n943), .B2(new_n682), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n682), .A2(G148gat), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n924), .A2(new_n485), .A3(new_n926), .A4(new_n946), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n947), .A2(KEYINPUT123), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n947), .A2(KEYINPUT123), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n945), .B1(new_n948), .B2(new_n949), .ZN(G1345gat));
  OAI21_X1  g749(.A(G155gat), .B1(new_n943), .B2(new_n588), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n588), .A2(G155gat), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n924), .A2(new_n485), .A3(new_n926), .A4(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n951), .A2(new_n953), .ZN(G1346gat));
  OAI211_X1 g753(.A(new_n650), .B(new_n906), .C1(new_n907), .C2(new_n917), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(G162gat), .ZN(new_n956));
  INV_X1    g755(.A(G162gat), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n924), .A2(new_n957), .A3(new_n898), .A4(new_n926), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT124), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n956), .A2(KEYINPUT124), .A3(new_n958), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(G1347gat));
  NOR2_X1   g762(.A1(new_n816), .A2(new_n485), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n880), .A2(new_n897), .A3(new_n964), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n965), .A2(new_n710), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n966), .A2(new_n218), .A3(new_n220), .ZN(new_n967));
  OR2_X1    g766(.A1(new_n967), .A2(KEYINPUT125), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(KEYINPUT125), .ZN(new_n969));
  OAI211_X1 g768(.A(new_n968), .B(new_n969), .C1(new_n212), .C2(new_n966), .ZN(G1348gat));
  NOR2_X1   g769(.A1(new_n965), .A2(new_n682), .ZN(new_n971));
  XNOR2_X1  g770(.A(new_n971), .B(new_n213), .ZN(G1349gat));
  OAI21_X1  g771(.A(new_n245), .B1(new_n965), .B2(new_n588), .ZN(new_n973));
  OR2_X1    g772(.A1(new_n965), .A2(new_n588), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n973), .B1(new_n974), .B2(new_n266), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT60), .ZN(new_n976));
  XNOR2_X1  g775(.A(new_n975), .B(new_n976), .ZN(G1350gat));
  INV_X1    g776(.A(KEYINPUT61), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n965), .A2(new_n652), .ZN(new_n979));
  INV_X1    g778(.A(G190gat), .ZN(new_n980));
  OAI211_X1 g779(.A(KEYINPUT126), .B(new_n978), .C1(new_n979), .C2(new_n980), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n979), .A2(new_n244), .ZN(new_n982));
  OAI21_X1  g781(.A(KEYINPUT126), .B1(new_n979), .B2(new_n980), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n983), .A2(KEYINPUT61), .ZN(new_n984));
  NOR3_X1   g783(.A1(new_n979), .A2(KEYINPUT126), .A3(new_n980), .ZN(new_n985));
  OAI211_X1 g784(.A(new_n981), .B(new_n982), .C1(new_n984), .C2(new_n985), .ZN(G1351gat));
  AND2_X1   g785(.A1(new_n880), .A2(new_n781), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n496), .A2(new_n964), .ZN(new_n988));
  INV_X1    g787(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n990), .A2(KEYINPUT127), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT127), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n987), .A2(new_n992), .A3(new_n989), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n991), .A2(new_n807), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g793(.A(new_n988), .B1(new_n938), .B2(new_n939), .ZN(new_n995));
  NOR2_X1   g794(.A1(new_n710), .A2(new_n300), .ZN(new_n996));
  AOI22_X1  g795(.A1(new_n994), .A2(new_n300), .B1(new_n995), .B2(new_n996), .ZN(G1352gat));
  INV_X1    g796(.A(new_n995), .ZN(new_n998));
  OAI21_X1  g797(.A(G204gat), .B1(new_n998), .B2(new_n682), .ZN(new_n999));
  NAND4_X1  g798(.A1(new_n987), .A2(new_n297), .A3(new_n681), .A4(new_n989), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n1000), .A2(KEYINPUT62), .ZN(new_n1001));
  OR2_X1    g800(.A1(new_n1000), .A2(KEYINPUT62), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n999), .A2(new_n1001), .A3(new_n1002), .ZN(G1353gat));
  AND2_X1   g802(.A1(new_n914), .A2(new_n935), .ZN(new_n1004));
  OAI21_X1  g803(.A(new_n856), .B1(new_n1004), .B2(new_n653), .ZN(new_n1005));
  AOI21_X1  g804(.A(KEYINPUT57), .B1(new_n1005), .B2(new_n781), .ZN(new_n1006));
  INV_X1    g805(.A(new_n939), .ZN(new_n1007));
  OAI211_X1 g806(.A(new_n653), .B(new_n989), .C1(new_n1006), .C2(new_n1007), .ZN(new_n1008));
  AND3_X1   g807(.A1(new_n1008), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1009));
  AOI21_X1  g808(.A(KEYINPUT63), .B1(new_n1008), .B2(G211gat), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n991), .A2(new_n993), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n653), .A2(new_n305), .ZN(new_n1012));
  OAI22_X1  g811(.A1(new_n1009), .A2(new_n1010), .B1(new_n1011), .B2(new_n1012), .ZN(G1354gat));
  OAI21_X1  g812(.A(G218gat), .B1(new_n998), .B2(new_n652), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n650), .A2(new_n306), .ZN(new_n1015));
  OAI21_X1  g814(.A(new_n1014), .B1(new_n1011), .B2(new_n1015), .ZN(G1355gat));
endmodule


