//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0 0 1 1 1 1 0 0 0 0 0 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1 0 0 0 1 0 1 0 1 1 1 1 0 0 1 1 1 0 0 1 1 0 0 1 1 0 0 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:51 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1278,
    new_n1279, new_n1281, new_n1282, new_n1283, new_n1284, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1340, new_n1341,
    new_n1342, new_n1343;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G58), .ZN(new_n216));
  INV_X1    g0016(.A(G68), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G50), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n220), .B1(new_n217), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n225));
  INV_X1    g0025(.A(G232), .ZN(new_n226));
  INV_X1    g0026(.A(G97), .ZN(new_n227));
  INV_X1    g0027(.A(G257), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n225), .B1(new_n216), .B2(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n209), .B1(new_n224), .B2(new_n229), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n212), .B1(new_n215), .B2(new_n219), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(new_n226), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT2), .B(G226), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n241), .B(new_n242), .Z(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  INV_X1    g0047(.A(KEYINPUT3), .ZN(new_n248));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  AOI21_X1  g0051(.A(G1698), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G222), .ZN(new_n253));
  INV_X1    g0053(.A(G77), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n250), .A2(new_n251), .ZN(new_n255));
  INV_X1    g0055(.A(G223), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(G1698), .ZN(new_n257));
  OAI221_X1 g0057(.A(new_n253), .B1(new_n254), .B2(new_n255), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G41), .ZN(new_n261));
  INV_X1    g0061(.A(G45), .ZN(new_n262));
  AOI21_X1  g0062(.A(G1), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G33), .A2(G41), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n264), .A2(G1), .A3(G13), .ZN(new_n265));
  AND3_X1   g0065(.A1(new_n263), .A2(new_n265), .A3(G274), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n259), .A2(new_n263), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n266), .B1(G226), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n260), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G190), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT10), .ZN(new_n271));
  OAI22_X1  g0071(.A1(new_n269), .A2(new_n270), .B1(KEYINPUT68), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G200), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n273), .B1(new_n260), .B2(new_n268), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT9), .ZN(new_n276));
  NAND3_X1  g0076(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n213), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT8), .B(G58), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT64), .ZN(new_n281));
  OR3_X1    g0081(.A1(new_n216), .A2(KEYINPUT64), .A3(KEYINPUT8), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(KEYINPUT65), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT65), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n281), .A2(new_n285), .A3(new_n282), .ZN(new_n286));
  NAND4_X1  g0086(.A1(new_n284), .A2(new_n207), .A3(G33), .A4(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(KEYINPUT66), .B1(new_n203), .B2(G20), .ZN(new_n288));
  AND3_X1   g0088(.A1(new_n203), .A2(KEYINPUT66), .A3(G20), .ZN(new_n289));
  NOR2_X1   g0089(.A1(G20), .A2(G33), .ZN(new_n290));
  AOI211_X1 g0090(.A(new_n288), .B(new_n289), .C1(G150), .C2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n279), .B1(new_n287), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n202), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n279), .B1(G1), .B2(new_n207), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n295), .B1(new_n296), .B2(new_n202), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n276), .B1(new_n292), .B2(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n292), .A2(new_n297), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(KEYINPUT9), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n275), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n301), .A2(KEYINPUT68), .A3(new_n271), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n271), .A2(KEYINPUT68), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n275), .A2(new_n300), .A3(new_n303), .A4(new_n298), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G169), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n269), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n307), .B1(G179), .B2(new_n269), .ZN(new_n308));
  OR2_X1    g0108(.A1(new_n308), .A2(new_n299), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n305), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT14), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n312), .A2(KEYINPUT70), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(G33), .A2(G97), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n226), .A2(G1698), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n316), .B1(G226), .B2(G1698), .ZN(new_n317));
  AND2_X1   g0117(.A1(KEYINPUT3), .A2(G33), .ZN(new_n318));
  NOR2_X1   g0118(.A1(KEYINPUT3), .A2(G33), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n315), .B1(new_n317), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n266), .B1(new_n321), .B2(new_n259), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT13), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT69), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n324), .B1(new_n259), .B2(new_n263), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n265), .A2(KEYINPUT69), .A3(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n325), .A2(G238), .A3(new_n327), .ZN(new_n328));
  AND3_X1   g0128(.A1(new_n322), .A2(new_n323), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n323), .B1(new_n322), .B2(new_n328), .ZN(new_n330));
  OAI211_X1 g0130(.A(G169), .B(new_n314), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n263), .A2(new_n265), .A3(G274), .ZN(new_n332));
  NOR2_X1   g0132(.A1(G226), .A2(G1698), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n333), .B1(new_n226), .B2(G1698), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n334), .A2(new_n255), .B1(G33), .B2(G97), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n332), .B1(new_n335), .B2(new_n265), .ZN(new_n336));
  AND3_X1   g0136(.A1(new_n325), .A2(G238), .A3(new_n327), .ZN(new_n337));
  OAI21_X1  g0137(.A(KEYINPUT13), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n322), .A2(new_n323), .A3(new_n328), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n338), .A2(G179), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n331), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n338), .A2(new_n339), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n314), .B1(new_n342), .B2(G169), .ZN(new_n343));
  OAI21_X1  g0143(.A(KEYINPUT71), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(G169), .B1(new_n329), .B2(new_n330), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n313), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT71), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n346), .A2(new_n347), .A3(new_n340), .A4(new_n331), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n217), .A2(G20), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n207), .A2(G33), .ZN(new_n351));
  INV_X1    g0151(.A(new_n290), .ZN(new_n352));
  OAI221_X1 g0152(.A(new_n350), .B1(new_n351), .B2(new_n254), .C1(new_n352), .C2(new_n202), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n278), .ZN(new_n354));
  XNOR2_X1  g0154(.A(new_n354), .B(KEYINPUT11), .ZN(new_n355));
  INV_X1    g0155(.A(G13), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n356), .A2(G1), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n357), .A2(KEYINPUT67), .A3(G20), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT67), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n293), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n279), .ZN(new_n362));
  OAI21_X1  g0162(.A(G68), .B1(new_n207), .B2(G1), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n355), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n357), .ZN(new_n365));
  NOR3_X1   g0165(.A1(new_n365), .A2(KEYINPUT12), .A3(new_n350), .ZN(new_n366));
  AND2_X1   g0166(.A1(new_n358), .A2(new_n360), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n217), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n366), .B1(new_n368), .B2(KEYINPUT12), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n364), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n349), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n342), .A2(G200), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n338), .A2(G190), .A3(new_n339), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n370), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n252), .A2(G232), .ZN(new_n376));
  INV_X1    g0176(.A(G107), .ZN(new_n377));
  OAI221_X1 g0177(.A(new_n376), .B1(new_n377), .B2(new_n255), .C1(new_n221), .C2(new_n257), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n259), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n266), .B1(G244), .B2(new_n267), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(new_n306), .ZN(new_n382));
  OAI22_X1  g0182(.A1(new_n280), .A2(new_n352), .B1(new_n207), .B2(new_n254), .ZN(new_n383));
  XNOR2_X1  g0183(.A(KEYINPUT15), .B(G87), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n384), .A2(new_n351), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n278), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(G77), .B1(new_n207), .B2(G1), .ZN(new_n387));
  OAI221_X1 g0187(.A(new_n386), .B1(G77), .B2(new_n361), .C1(new_n362), .C2(new_n387), .ZN(new_n388));
  AND2_X1   g0188(.A1(new_n382), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(G179), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n379), .A2(new_n390), .A3(new_n380), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n388), .B1(new_n381), .B2(G200), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n393), .B1(new_n270), .B2(new_n381), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n311), .A2(new_n372), .A3(new_n375), .A4(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT75), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT73), .ZN(new_n398));
  NOR2_X1   g0198(.A1(G223), .A2(G1698), .ZN(new_n399));
  INV_X1    g0199(.A(G226), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n399), .B1(new_n400), .B2(G1698), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n401), .A2(new_n255), .B1(G33), .B2(G87), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n398), .B1(new_n402), .B2(new_n265), .ZN(new_n403));
  INV_X1    g0203(.A(G1698), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n256), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n400), .A2(G1698), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n405), .B(new_n406), .C1(new_n318), .C2(new_n319), .ZN(new_n407));
  NAND2_X1  g0207(.A1(G33), .A2(G87), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n265), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(KEYINPUT73), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n403), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n265), .A2(G232), .A3(new_n326), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n332), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(KEYINPUT74), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT74), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n332), .A2(new_n412), .A3(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n414), .A2(new_n390), .A3(new_n416), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n411), .A2(new_n417), .ZN(new_n418));
  AND3_X1   g0218(.A1(new_n332), .A2(new_n412), .A3(new_n415), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n415), .B1(new_n332), .B2(new_n412), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n409), .ZN(new_n422));
  AOI21_X1  g0222(.A(G169), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n397), .B1(new_n418), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n414), .A2(new_n422), .A3(new_n416), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(new_n306), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n426), .B(KEYINPUT75), .C1(new_n411), .C2(new_n417), .ZN(new_n427));
  AND3_X1   g0227(.A1(new_n281), .A2(new_n285), .A3(new_n282), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n285), .B1(new_n281), .B2(new_n282), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n293), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n284), .A2(new_n286), .A3(new_n296), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n250), .A2(new_n207), .A3(new_n251), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT7), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n250), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n251), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n435), .A2(KEYINPUT72), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT72), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n433), .A2(new_n438), .A3(new_n434), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n437), .A2(G68), .A3(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n216), .A2(new_n217), .ZN(new_n441));
  OAI21_X1  g0241(.A(G20), .B1(new_n441), .B2(new_n201), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n290), .A2(G159), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(KEYINPUT16), .B1(new_n440), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(KEYINPUT7), .B1(new_n320), .B2(new_n207), .ZN(new_n447));
  INV_X1    g0247(.A(new_n436), .ZN(new_n448));
  OAI21_X1  g0248(.A(G68), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n449), .A2(KEYINPUT16), .A3(new_n445), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n278), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n432), .B1(new_n446), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n424), .A2(new_n427), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT18), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT18), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n424), .A2(new_n427), .A3(new_n452), .A4(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  AND2_X1   g0257(.A1(new_n430), .A2(new_n431), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n440), .A2(new_n445), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT16), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n435), .A2(new_n436), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n444), .B1(new_n462), .B2(G68), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n279), .B1(new_n463), .B2(KEYINPUT16), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n458), .B1(new_n461), .B2(new_n464), .ZN(new_n465));
  NOR3_X1   g0265(.A1(new_n419), .A2(new_n420), .A3(new_n409), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n414), .A2(new_n270), .A3(new_n416), .ZN(new_n467));
  OAI22_X1  g0267(.A1(G200), .A2(new_n466), .B1(new_n411), .B2(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(KEYINPUT17), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  AND2_X1   g0269(.A1(new_n403), .A2(new_n410), .ZN(new_n470));
  INV_X1    g0270(.A(new_n467), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n470), .A2(new_n471), .B1(new_n425), .B2(new_n273), .ZN(new_n472));
  OAI21_X1  g0272(.A(KEYINPUT76), .B1(new_n452), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n461), .A2(new_n464), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT76), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n474), .A2(new_n475), .A3(new_n432), .A4(new_n468), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n469), .B1(new_n477), .B2(KEYINPUT17), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NOR3_X1   g0279(.A1(new_n396), .A2(new_n457), .A3(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(G274), .ZN(new_n481));
  INV_X1    g0281(.A(new_n213), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n481), .B1(new_n482), .B2(new_n264), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n262), .A2(G1), .ZN(new_n484));
  XNOR2_X1  g0284(.A(KEYINPUT5), .B(G41), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n484), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n265), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n486), .B1(new_n488), .B2(new_n228), .ZN(new_n489));
  AND2_X1   g0289(.A1(KEYINPUT4), .A2(G244), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n252), .A2(new_n490), .B1(G33), .B2(G283), .ZN(new_n491));
  OAI211_X1 g0291(.A(G244), .B(new_n404), .C1(new_n318), .C2(new_n319), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI211_X1 g0294(.A(G250), .B(G1698), .C1(new_n318), .C2(new_n319), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(KEYINPUT79), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT79), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n255), .A2(new_n497), .A3(G250), .A4(G1698), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n491), .A2(new_n494), .A3(new_n496), .A4(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n489), .B1(new_n499), .B2(new_n259), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n390), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n252), .A2(new_n490), .ZN(new_n502));
  NAND2_X1  g0302(.A1(G33), .A2(G283), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n494), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n496), .A2(new_n498), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n259), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n489), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n306), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n290), .A2(G77), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT77), .ZN(new_n511));
  XNOR2_X1  g0311(.A(new_n510), .B(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT6), .ZN(new_n513));
  NOR3_X1   g0313(.A1(new_n513), .A2(new_n227), .A3(G107), .ZN(new_n514));
  XNOR2_X1  g0314(.A(G97), .B(G107), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n514), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n512), .B1(new_n207), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n437), .A2(G107), .A3(new_n439), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n517), .B1(new_n518), .B2(KEYINPUT78), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT78), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n437), .A2(new_n520), .A3(G107), .A4(new_n439), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n279), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n294), .A2(new_n227), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n279), .B(new_n293), .C1(G1), .C2(new_n249), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n523), .B1(new_n524), .B2(new_n227), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n501), .B(new_n509), .C1(new_n522), .C2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n519), .A2(new_n521), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n278), .ZN(new_n528));
  INV_X1    g0328(.A(new_n525), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n506), .A2(new_n270), .A3(new_n507), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(G200), .B2(new_n500), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n528), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(G20), .B1(new_n250), .B2(new_n251), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(G68), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT19), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n207), .B1(new_n315), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n222), .A2(new_n227), .A3(new_n377), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n207), .A2(G33), .A3(G97), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n539), .A2(KEYINPUT81), .A3(new_n535), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(KEYINPUT81), .B1(new_n539), .B2(new_n535), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n534), .B(new_n538), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n278), .ZN(new_n544));
  INV_X1    g0344(.A(new_n384), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n361), .A2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n544), .A2(KEYINPUT82), .A3(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT82), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n539), .A2(new_n535), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT81), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n540), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n533), .A2(G68), .B1(new_n536), .B2(new_n537), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n279), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n549), .B1(new_n555), .B2(new_n546), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n548), .A2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(new_n524), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n545), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT80), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n561), .B1(new_n262), .B2(G1), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n206), .A2(KEYINPUT80), .A3(G45), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n265), .A2(new_n562), .A3(G250), .A4(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n265), .A2(G274), .ZN(new_n565));
  INV_X1    g0365(.A(new_n484), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  OAI211_X1 g0367(.A(G244), .B(G1698), .C1(new_n318), .C2(new_n319), .ZN(new_n568));
  OAI211_X1 g0368(.A(G238), .B(new_n404), .C1(new_n318), .C2(new_n319), .ZN(new_n569));
  INV_X1    g0369(.A(G116), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n568), .B(new_n569), .C1(new_n249), .C2(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n567), .B1(new_n259), .B2(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n572), .A2(G169), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n573), .B1(new_n390), .B2(new_n572), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n560), .A2(new_n574), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n548), .A2(new_n556), .B1(G87), .B2(new_n558), .ZN(new_n576));
  AOI21_X1  g0376(.A(KEYINPUT83), .B1(new_n572), .B2(G190), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n571), .A2(new_n259), .ZN(new_n578));
  INV_X1    g0378(.A(new_n567), .ZN(new_n579));
  AND4_X1   g0379(.A1(KEYINPUT83), .A2(new_n578), .A3(new_n579), .A4(G190), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n578), .A2(new_n579), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(G200), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n576), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  AND4_X1   g0384(.A1(new_n526), .A2(new_n532), .A3(new_n575), .A4(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n503), .B(new_n207), .C1(G33), .C2(new_n227), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(KEYINPUT85), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n249), .A2(G97), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT85), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n588), .A2(new_n589), .A3(new_n207), .A4(new_n503), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n570), .A2(G20), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n587), .A2(new_n278), .A3(new_n590), .A4(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT20), .ZN(new_n593));
  XNOR2_X1  g0393(.A(new_n592), .B(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n570), .B1(new_n206), .B2(G33), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  OAI22_X1  g0396(.A1(new_n362), .A2(new_n596), .B1(G116), .B2(new_n361), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n255), .A2(G257), .A3(new_n404), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(KEYINPUT84), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT84), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n252), .A2(new_n602), .A3(G257), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n320), .A2(G303), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n255), .A2(G264), .A3(G1698), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n601), .A2(new_n603), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n259), .ZN(new_n607));
  INV_X1    g0407(.A(G270), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n486), .B1(new_n488), .B2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n599), .A2(G169), .A3(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT21), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n609), .B1(new_n606), .B2(new_n259), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n599), .A2(G179), .A3(new_n615), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n599), .A2(new_n611), .A3(KEYINPUT21), .A4(G169), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n615), .A2(G190), .ZN(new_n618));
  XNOR2_X1  g0418(.A(new_n592), .B(KEYINPUT20), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n619), .A2(new_n597), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n618), .B(new_n620), .C1(new_n273), .C2(new_n615), .ZN(new_n621));
  AND4_X1   g0421(.A1(new_n614), .A2(new_n616), .A3(new_n617), .A4(new_n621), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n207), .B(G87), .C1(new_n318), .C2(new_n319), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(KEYINPUT22), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT22), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n255), .A2(new_n625), .A3(new_n207), .A4(G87), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT24), .ZN(new_n628));
  NOR3_X1   g0428(.A1(new_n249), .A2(new_n570), .A3(G20), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT23), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(new_n207), .B2(G107), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n377), .A2(KEYINPUT23), .A3(G20), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n629), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n627), .A2(new_n628), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n628), .B1(new_n627), .B2(new_n633), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n278), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n294), .A2(new_n377), .ZN(new_n637));
  XNOR2_X1  g0437(.A(new_n637), .B(KEYINPUT25), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n638), .B1(G107), .B2(new_n558), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n487), .A2(G264), .A3(new_n265), .ZN(new_n641));
  NOR2_X1   g0441(.A1(G250), .A2(G1698), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n642), .B1(new_n228), .B2(G1698), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n643), .A2(new_n255), .B1(G33), .B2(G294), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n641), .B(new_n486), .C1(new_n644), .C2(new_n265), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n306), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n643), .A2(new_n255), .ZN(new_n647));
  NAND2_X1  g0447(.A1(G33), .A2(G294), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n259), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n650), .A2(new_n390), .A3(new_n486), .A4(new_n641), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n646), .A2(new_n651), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n640), .A2(KEYINPUT86), .A3(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(KEYINPUT86), .B1(new_n640), .B2(new_n652), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n645), .A2(G200), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n655), .B1(new_n270), .B2(new_n645), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n640), .A2(new_n656), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n653), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  AND4_X1   g0458(.A1(new_n480), .A2(new_n585), .A3(new_n622), .A4(new_n658), .ZN(G372));
  INV_X1    g0459(.A(KEYINPUT26), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n583), .A2(KEYINPUT87), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT87), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n582), .A2(new_n662), .A3(G200), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n576), .A2(new_n581), .A3(new_n661), .A4(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n575), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n660), .B1(new_n665), .B2(new_n526), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT88), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n528), .A2(new_n529), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n509), .A2(new_n501), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n575), .A2(new_n584), .A3(new_n669), .A4(new_n670), .ZN(new_n671));
  XOR2_X1   g0471(.A(KEYINPUT89), .B(KEYINPUT26), .Z(new_n672));
  OR2_X1    g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  OAI211_X1 g0473(.A(KEYINPUT88), .B(new_n660), .C1(new_n665), .C2(new_n526), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n668), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n575), .ZN(new_n676));
  OAI211_X1 g0476(.A(new_n664), .B(new_n575), .C1(new_n640), .C2(new_n656), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n532), .A2(new_n526), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AND3_X1   g0479(.A1(new_n614), .A2(new_n616), .A3(new_n617), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n640), .A2(new_n652), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n676), .B1(new_n679), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n675), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n480), .A2(new_n684), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n454), .A2(new_n456), .ZN(new_n686));
  INV_X1    g0486(.A(new_n392), .ZN(new_n687));
  AOI22_X1  g0487(.A1(new_n349), .A2(new_n371), .B1(new_n687), .B2(new_n375), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n686), .B1(new_n688), .B2(new_n479), .ZN(new_n689));
  OR2_X1    g0489(.A1(new_n689), .A2(KEYINPUT90), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n305), .B1(new_n689), .B2(KEYINPUT90), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n310), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n685), .A2(new_n692), .ZN(G369));
  INV_X1    g0493(.A(new_n680), .ZN(new_n694));
  OR3_X1    g0494(.A1(new_n365), .A2(KEYINPUT27), .A3(G20), .ZN(new_n695));
  OAI21_X1  g0495(.A(KEYINPUT27), .B1(new_n365), .B2(G20), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(G213), .A3(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(G343), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n620), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n694), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n622), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n702), .B1(new_n703), .B2(new_n701), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(G330), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n640), .A2(new_n699), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n658), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n681), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(new_n699), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n706), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n680), .A2(new_n699), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n658), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(new_n681), .B2(new_n699), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n712), .A2(new_n716), .ZN(G399));
  INV_X1    g0517(.A(new_n210), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(G41), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(new_n206), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n537), .A2(G116), .ZN(new_n721));
  INV_X1    g0521(.A(new_n219), .ZN(new_n722));
  AOI22_X1  g0522(.A1(new_n720), .A2(new_n721), .B1(new_n722), .B2(new_n719), .ZN(new_n723));
  XOR2_X1   g0523(.A(new_n723), .B(KEYINPUT28), .Z(new_n724));
  XNOR2_X1  g0524(.A(new_n678), .B(KEYINPUT93), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n653), .A2(new_n654), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n677), .B1(new_n680), .B2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n676), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n671), .A2(new_n672), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(KEYINPUT92), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT92), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n671), .A2(new_n731), .A3(new_n672), .ZN(new_n732));
  OR3_X1    g0532(.A1(new_n665), .A2(new_n660), .A3(new_n526), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n730), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n699), .B1(new_n728), .B2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT29), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n585), .A2(new_n622), .A3(new_n658), .A4(new_n700), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n615), .A2(G179), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n259), .B1(new_n484), .B2(new_n485), .ZN(new_n741));
  AOI22_X1  g0541(.A1(new_n649), .A2(new_n259), .B1(new_n741), .B2(G264), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n506), .A2(new_n507), .A3(new_n572), .A4(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(KEYINPUT91), .B1(new_n740), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(KEYINPUT30), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT30), .ZN(new_n746));
  OAI211_X1 g0546(.A(KEYINPUT91), .B(new_n746), .C1(new_n740), .C2(new_n743), .ZN(new_n747));
  AND2_X1   g0547(.A1(new_n645), .A2(new_n390), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n611), .A2(new_n508), .A3(new_n748), .A4(new_n582), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n745), .A2(new_n747), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(new_n699), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT31), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n750), .A2(KEYINPUT31), .A3(new_n699), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n739), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G330), .ZN(new_n756));
  AOI211_X1 g0556(.A(KEYINPUT29), .B(new_n699), .C1(new_n675), .C2(new_n683), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n738), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n724), .B1(new_n760), .B2(G1), .ZN(G364));
  NOR2_X1   g0561(.A1(new_n356), .A2(G20), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n762), .B(KEYINPUT94), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G45), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n720), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n706), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n767), .B1(G330), .B2(new_n704), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n210), .A2(new_n255), .ZN(new_n769));
  INV_X1    g0569(.A(G355), .ZN(new_n770));
  OAI22_X1  g0570(.A1(new_n769), .A2(new_n770), .B1(G116), .B2(new_n210), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n718), .A2(new_n255), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n773), .B1(new_n262), .B2(new_n722), .ZN(new_n774));
  OR2_X1    g0574(.A1(new_n243), .A2(new_n262), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n771), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G13), .A2(G33), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G20), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n213), .B1(G20), .B2(new_n306), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n776), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n765), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n207), .A2(new_n390), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR3_X1   g0586(.A1(new_n786), .A2(G190), .A3(new_n273), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n217), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n785), .A2(new_n270), .A3(new_n273), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n785), .A2(G190), .A3(new_n273), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n255), .B1(new_n790), .B2(new_n254), .C1(new_n216), .C2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n207), .A2(G179), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n793), .A2(new_n270), .A3(G200), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n377), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n793), .A2(G190), .A3(G200), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n222), .ZN(new_n797));
  NOR4_X1   g0597(.A1(new_n789), .A2(new_n792), .A3(new_n795), .A4(new_n797), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n785), .A2(G190), .A3(G200), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n799), .A2(KEYINPUT95), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n799), .A2(KEYINPUT95), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(G179), .A2(G200), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n207), .B1(new_n804), .B2(G190), .ZN(new_n805));
  AND2_X1   g0605(.A1(new_n805), .A2(KEYINPUT97), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n805), .A2(KEYINPUT97), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n803), .A2(G50), .B1(new_n809), .B2(G97), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n804), .A2(G20), .A3(new_n270), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT96), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n811), .A2(new_n812), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(G159), .ZN(new_n816));
  OAI21_X1  g0616(.A(KEYINPUT32), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  OR3_X1    g0617(.A1(new_n815), .A2(KEYINPUT32), .A3(new_n816), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n798), .A2(new_n810), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT98), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n802), .B(new_n820), .ZN(new_n821));
  AND2_X1   g0621(.A1(new_n821), .A2(G326), .ZN(new_n822));
  INV_X1    g0622(.A(G311), .ZN(new_n823));
  INV_X1    g0623(.A(G322), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n320), .B1(new_n790), .B2(new_n823), .C1(new_n824), .C2(new_n791), .ZN(new_n825));
  INV_X1    g0625(.A(new_n815), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n825), .B1(G329), .B2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(G283), .ZN(new_n828));
  INV_X1    g0628(.A(G303), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n794), .A2(new_n828), .B1(new_n796), .B2(new_n829), .ZN(new_n830));
  XNOR2_X1  g0630(.A(KEYINPUT33), .B(G317), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n830), .B1(new_n787), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(G294), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n827), .B(new_n832), .C1(new_n833), .C2(new_n808), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n819), .B1(new_n822), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n835), .A2(KEYINPUT99), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(KEYINPUT99), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(new_n780), .ZN(new_n838));
  INV_X1    g0638(.A(new_n779), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n784), .B1(new_n836), .B2(new_n838), .C1(new_n704), .C2(new_n839), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n768), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(G396));
  AOI21_X1  g0642(.A(new_n699), .B1(new_n675), .B2(new_n683), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n388), .A2(new_n699), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n395), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT101), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(new_n392), .B2(new_n700), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n389), .A2(KEYINPUT101), .A3(new_n391), .A4(new_n699), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n845), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n843), .B(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n766), .B1(new_n851), .B2(new_n756), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n756), .B2(new_n851), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n320), .B1(new_n826), .B2(G132), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(KEYINPUT100), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n794), .A2(new_n217), .ZN(new_n858));
  INV_X1    g0658(.A(new_n796), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n858), .B1(G50), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n860), .B1(new_n216), .B2(new_n808), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n855), .A2(KEYINPUT100), .ZN(new_n862));
  NOR3_X1   g0662(.A1(new_n857), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n791), .ZN(new_n865));
  INV_X1    g0665(.A(new_n790), .ZN(new_n866));
  AOI22_X1  g0666(.A1(G143), .A2(new_n865), .B1(new_n866), .B2(G159), .ZN(new_n867));
  INV_X1    g0667(.A(G150), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n867), .B1(new_n868), .B2(new_n788), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n869), .B1(G137), .B2(new_n803), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n870), .B(KEYINPUT34), .ZN(new_n871));
  OAI221_X1 g0671(.A(new_n320), .B1(new_n790), .B2(new_n570), .C1(new_n833), .C2(new_n791), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(G311), .B2(new_n826), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n794), .A2(new_n222), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n874), .B1(new_n787), .B2(G283), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n873), .B(new_n875), .C1(new_n377), .C2(new_n796), .ZN(new_n876));
  OAI22_X1  g0676(.A1(new_n802), .A2(new_n829), .B1(new_n808), .B2(new_n227), .ZN(new_n877));
  OAI22_X1  g0677(.A1(new_n864), .A2(new_n871), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n780), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n780), .A2(new_n777), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n765), .B1(new_n254), .B2(new_n880), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n879), .B(new_n881), .C1(new_n850), .C2(new_n778), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n853), .A2(new_n882), .ZN(G384));
  NOR2_X1   g0683(.A1(new_n763), .A2(new_n206), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n371), .A2(new_n699), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n372), .A2(new_n375), .A3(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n375), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n371), .B(new_n699), .C1(new_n349), .C2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  AND3_X1   g0689(.A1(new_n889), .A2(new_n755), .A3(new_n850), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT38), .ZN(new_n891));
  INV_X1    g0691(.A(new_n697), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n449), .A2(new_n445), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT103), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT16), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n463), .A2(KEYINPUT103), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n451), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n892), .B1(new_n897), .B2(new_n458), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(new_n686), .B2(new_n478), .ZN(new_n899));
  INV_X1    g0699(.A(new_n477), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT37), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n452), .A2(new_n892), .ZN(new_n902));
  AND3_X1   g0702(.A1(new_n453), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n424), .B(new_n427), .C1(new_n897), .C2(new_n458), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n904), .A2(new_n473), .A3(new_n476), .A4(new_n898), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n900), .A2(new_n903), .B1(new_n905), .B2(KEYINPUT37), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n891), .B1(new_n899), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n903), .A2(new_n900), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n895), .A2(new_n896), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n458), .B1(new_n909), .B2(new_n464), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n424), .A2(new_n427), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n910), .B1(new_n911), .B2(new_n697), .ZN(new_n912));
  OAI21_X1  g0712(.A(KEYINPUT37), .B1(new_n912), .B2(new_n477), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n908), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT17), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n915), .B1(new_n473), .B2(new_n476), .ZN(new_n916));
  NOR3_X1   g0716(.A1(new_n457), .A2(new_n916), .A3(new_n469), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n914), .B(KEYINPUT38), .C1(new_n917), .C2(new_n898), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n907), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT40), .B1(new_n890), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n902), .B1(new_n686), .B2(new_n478), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n453), .B(new_n902), .C1(new_n452), .C2(new_n472), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n903), .A2(new_n900), .B1(new_n922), .B2(KEYINPUT37), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n891), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n924), .A2(new_n918), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n889), .A2(new_n755), .A3(KEYINPUT40), .A4(new_n850), .ZN(new_n926));
  OAI21_X1  g0726(.A(KEYINPUT104), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n924), .A2(new_n918), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT104), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n890), .A2(new_n928), .A3(new_n929), .A4(KEYINPUT40), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n920), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  XOR2_X1   g0731(.A(new_n931), .B(KEYINPUT105), .Z(new_n932));
  NAND2_X1  g0732(.A1(new_n480), .A2(new_n755), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n932), .A2(new_n933), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n934), .A2(G330), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n843), .A2(new_n850), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n392), .A2(new_n699), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n940), .A2(new_n919), .A3(new_n889), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT39), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n928), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n372), .A2(new_n699), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n907), .A2(new_n918), .A3(KEYINPUT39), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n457), .A2(new_n697), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n941), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n480), .B1(new_n737), .B2(new_n757), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n692), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n948), .B(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n884), .B1(new_n936), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n951), .B2(new_n936), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT35), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n516), .A2(new_n954), .ZN(new_n955));
  AOI211_X1 g0755(.A(new_n570), .B(new_n215), .C1(new_n516), .C2(new_n954), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n955), .B1(new_n957), .B2(KEYINPUT102), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(KEYINPUT102), .B2(new_n957), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT36), .ZN(new_n960));
  NOR3_X1   g0760(.A1(new_n219), .A2(new_n254), .A3(new_n441), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n217), .A2(G50), .ZN(new_n962));
  OAI211_X1 g0762(.A(G1), .B(new_n356), .C1(new_n961), .C2(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n953), .A2(new_n960), .A3(new_n963), .ZN(G367));
  OAI221_X1 g0764(.A(new_n781), .B1(new_n210), .B2(new_n384), .C1(new_n773), .C2(new_n239), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n766), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT46), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n796), .B2(new_n570), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n859), .A2(KEYINPUT46), .A3(G116), .ZN(new_n969));
  INV_X1    g0769(.A(G317), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n968), .B(new_n969), .C1(new_n815), .C2(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n794), .A2(new_n227), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n320), .B1(new_n790), .B2(new_n828), .C1(new_n829), .C2(new_n791), .ZN(new_n973));
  AOI211_X1 g0773(.A(new_n972), .B(new_n973), .C1(G294), .C2(new_n787), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n377), .B2(new_n808), .ZN(new_n975));
  AOI211_X1 g0775(.A(new_n971), .B(new_n975), .C1(G311), .C2(new_n821), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n808), .A2(new_n217), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n788), .A2(new_n816), .B1(new_n216), .B2(new_n796), .ZN(new_n978));
  INV_X1    g0778(.A(new_n794), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n978), .B1(G77), .B2(new_n979), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n255), .B1(new_n790), .B2(new_n202), .C1(new_n868), .C2(new_n791), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(G137), .B2(new_n826), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n977), .B(new_n983), .C1(G143), .C2(new_n821), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n976), .A2(new_n984), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n985), .B(KEYINPUT47), .Z(new_n986));
  AOI21_X1  g0786(.A(new_n966), .B1(new_n986), .B2(new_n780), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n576), .A2(new_n700), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n676), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(new_n665), .B2(new_n988), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT106), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n779), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n987), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n764), .A2(G1), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT45), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n669), .A2(new_n699), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n725), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n669), .A2(new_n670), .A3(new_n699), .ZN(new_n998));
  AND2_X1   g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n995), .B1(new_n999), .B2(new_n715), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n997), .A2(new_n998), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n716), .A2(new_n1001), .A3(KEYINPUT45), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n999), .A2(KEYINPUT44), .A3(new_n715), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT44), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n716), .B2(new_n1001), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1003), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n712), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1008), .B(new_n1009), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n708), .B(new_n710), .C1(new_n680), .C2(new_n699), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT108), .ZN(new_n1012));
  AND2_X1   g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n714), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(new_n706), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1016), .A2(new_n759), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  NOR3_X1   g0818(.A1(new_n1010), .A2(new_n1018), .A3(KEYINPUT109), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT109), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1008), .B(new_n712), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1020), .B1(new_n1021), .B2(new_n1017), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n760), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n719), .B(KEYINPUT41), .Z(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n994), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1001), .A2(new_n658), .A3(new_n713), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n1027), .A2(KEYINPUT42), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT107), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n526), .B1(new_n997), .B2(new_n726), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n1027), .A2(KEYINPUT42), .B1(new_n1030), .B2(new_n700), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT43), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n991), .A2(new_n1033), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n991), .A2(new_n1033), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1032), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n712), .A2(new_n999), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1029), .A2(new_n1033), .A3(new_n991), .A4(new_n1031), .ZN(new_n1038));
  AND3_X1   g0838(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1037), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n993), .B1(new_n1026), .B2(new_n1042), .ZN(G387));
  INV_X1    g0843(.A(new_n994), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n1016), .A2(new_n1044), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n769), .A2(new_n721), .B1(G107), .B2(new_n210), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n236), .A2(new_n262), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n721), .ZN(new_n1048));
  AOI211_X1 g0848(.A(G45), .B(new_n1048), .C1(G68), .C2(G77), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n280), .A2(G50), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT50), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n773), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1046), .B1(new_n1047), .B2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n766), .B1(new_n1053), .B2(new_n782), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n428), .A2(new_n429), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n1055), .A2(new_n787), .B1(G68), .B2(new_n866), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT110), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n815), .A2(new_n868), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n796), .A2(new_n254), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n255), .B1(new_n791), .B2(new_n202), .ZN(new_n1060));
  NOR4_X1   g0860(.A1(new_n1058), .A2(new_n972), .A3(new_n1059), .A4(new_n1060), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n803), .A2(G159), .B1(new_n809), .B2(new_n545), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1057), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n809), .A2(G283), .B1(G294), .B2(new_n859), .ZN(new_n1064));
  XOR2_X1   g0864(.A(KEYINPUT111), .B(G322), .Z(new_n1065));
  NAND2_X1  g0865(.A1(new_n821), .A2(new_n1065), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n791), .A2(new_n970), .B1(new_n790), .B2(new_n829), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(G311), .B2(new_n787), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT112), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT48), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1064), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  XOR2_X1   g0873(.A(new_n1073), .B(KEYINPUT113), .Z(new_n1074));
  NAND2_X1  g0874(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1074), .A2(KEYINPUT49), .A3(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n320), .B1(new_n794), .B2(new_n570), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(new_n826), .B2(G326), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(KEYINPUT49), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1063), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1054), .B1(new_n1081), .B2(new_n780), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT114), .ZN(new_n1083));
  OR2_X1    g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n711), .A2(new_n839), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1045), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1016), .A2(new_n759), .ZN(new_n1088));
  XOR2_X1   g0888(.A(new_n719), .B(KEYINPUT115), .Z(new_n1089));
  NAND3_X1  g0889(.A1(new_n1018), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1087), .A2(new_n1090), .ZN(G393));
  AOI211_X1 g0891(.A(new_n255), .B(new_n795), .C1(G294), .C2(new_n866), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n826), .A2(new_n1065), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n787), .A2(G303), .B1(G283), .B2(new_n859), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1092), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n802), .A2(new_n970), .B1(new_n823), .B2(new_n791), .ZN(new_n1096));
  XOR2_X1   g0896(.A(new_n1096), .B(KEYINPUT52), .Z(new_n1097));
  AOI211_X1 g0897(.A(new_n1095), .B(new_n1097), .C1(G116), .C2(new_n809), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n803), .A2(G150), .B1(G159), .B2(new_n865), .ZN(new_n1099));
  XOR2_X1   g0899(.A(KEYINPUT116), .B(KEYINPUT51), .Z(new_n1100));
  AND2_X1   g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n809), .A2(G77), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n826), .A2(G143), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n255), .B1(new_n790), .B2(new_n280), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1105), .A2(new_n874), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n787), .A2(G50), .B1(G68), .B2(new_n859), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1103), .A2(new_n1104), .A3(new_n1106), .A4(new_n1107), .ZN(new_n1108));
  NOR3_X1   g0908(.A1(new_n1101), .A2(new_n1102), .A3(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n780), .B1(new_n1098), .B2(new_n1109), .ZN(new_n1110));
  AND2_X1   g0910(.A1(new_n772), .A2(new_n246), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n781), .B1(new_n227), .B2(new_n210), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1110), .B(new_n766), .C1(new_n1111), .C2(new_n1112), .ZN(new_n1113));
  XOR2_X1   g0913(.A(new_n1113), .B(KEYINPUT117), .Z(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n1001), .B2(new_n839), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n1010), .B2(new_n1044), .ZN(new_n1116));
  OAI21_X1  g0916(.A(KEYINPUT109), .B1(new_n1010), .B2(new_n1018), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1021), .A2(new_n1020), .A3(new_n1017), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1089), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(new_n1010), .B2(new_n1018), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1116), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(G390));
  INV_X1    g0923(.A(new_n944), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n938), .B1(new_n843), .B2(new_n850), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n889), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1124), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n943), .A2(new_n945), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n755), .A2(G330), .A3(new_n850), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1130), .A2(new_n1126), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(KEYINPUT118), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT118), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1133), .B1(new_n1130), .B2(new_n1126), .ZN(new_n1134));
  AND2_X1   g0934(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n925), .A2(new_n944), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n938), .B1(new_n735), .B2(new_n850), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1136), .B1(new_n1137), .B2(new_n1126), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1129), .A2(new_n1135), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1131), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n395), .A2(new_n844), .B1(new_n847), .B2(new_n848), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n699), .B(new_n1141), .C1(new_n728), .C2(new_n734), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n889), .B1(new_n1142), .B2(new_n938), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n1127), .A2(new_n1128), .B1(new_n1143), .B2(new_n1136), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1139), .B(new_n994), .C1(new_n1140), .C2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT119), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1145), .B(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1139), .B1(new_n1140), .B2(new_n1144), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n480), .A2(G330), .A3(new_n755), .ZN(new_n1149));
  AND3_X1   g0949(.A1(new_n949), .A2(new_n692), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1130), .A2(new_n1126), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1132), .A2(new_n1137), .A3(new_n1134), .A4(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1151), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n940), .B1(new_n1153), .B2(new_n1131), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1150), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1148), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1129), .A2(new_n1138), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n1131), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1159), .A2(new_n1139), .A3(new_n1150), .A4(new_n1155), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1157), .A2(new_n1160), .A3(new_n1089), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n880), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n766), .B1(new_n1055), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n803), .A2(G128), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n809), .A2(G159), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(KEYINPUT54), .B(G143), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n255), .B1(new_n790), .B2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(G132), .B2(new_n865), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n787), .A2(G137), .B1(G50), .B2(new_n979), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1164), .A2(new_n1165), .A3(new_n1168), .A4(new_n1169), .ZN(new_n1170));
  OR3_X1    g0970(.A1(new_n796), .A2(KEYINPUT53), .A3(new_n868), .ZN(new_n1171));
  OAI21_X1  g0971(.A(KEYINPUT53), .B1(new_n796), .B2(new_n868), .ZN(new_n1172));
  INV_X1    g0972(.A(G125), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1171), .B(new_n1172), .C1(new_n815), .C2(new_n1173), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n797), .B(new_n858), .C1(G107), .C2(new_n787), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n320), .B1(new_n790), .B2(new_n227), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(G116), .B2(new_n865), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1175), .B(new_n1177), .C1(new_n833), .C2(new_n815), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1103), .B1(new_n828), .B2(new_n802), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n1170), .A2(new_n1174), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1163), .B1(new_n1180), .B2(new_n780), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1128), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1181), .B1(new_n1182), .B2(new_n778), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1147), .A2(new_n1161), .A3(new_n1183), .ZN(G378));
  NAND2_X1  g0984(.A1(new_n927), .A2(new_n930), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n920), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT121), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n892), .B1(new_n292), .B2(new_n297), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n305), .B2(new_n310), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n302), .A2(new_n304), .A3(new_n309), .A4(new_n1188), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1192));
  AND3_X1   g0992(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1192), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1187), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1192), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1198), .A2(KEYINPUT121), .A3(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1195), .A2(new_n1200), .ZN(new_n1201));
  AND4_X1   g1001(.A1(G330), .A2(new_n1185), .A3(new_n1186), .A4(new_n1201), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(new_n931), .B2(G330), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n948), .B1(new_n1202), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n930), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n926), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n929), .B1(new_n1208), .B2(new_n928), .ZN(new_n1209));
  OAI211_X1 g1009(.A(G330), .B(new_n1186), .C1(new_n1207), .C2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(new_n1203), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n948), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n931), .A2(G330), .A3(new_n1201), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1206), .A2(KEYINPUT122), .A3(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1150), .B1(new_n1148), .B2(new_n1156), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT122), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1217), .B(new_n948), .C1(new_n1202), .C2(new_n1205), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1215), .A2(new_n1216), .A3(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT57), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1220), .B1(new_n1160), .B2(new_n1150), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1206), .A2(new_n1214), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1120), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1221), .A2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1215), .A2(new_n994), .A3(new_n1218), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n766), .B1(G50), .B2(new_n1162), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n255), .A2(G41), .ZN(new_n1228));
  AOI211_X1 g1028(.A(G50), .B(new_n1228), .C1(new_n249), .C2(new_n261), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n1228), .B1(new_n791), .B2(new_n377), .C1(new_n384), .C2(new_n790), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(G283), .B2(new_n826), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n794), .A2(new_n216), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n1059), .B(new_n1232), .C1(G97), .C2(new_n787), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1231), .A2(new_n1233), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n977), .B(new_n1234), .C1(G116), .C2(new_n803), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1229), .B1(new_n1235), .B2(KEYINPUT58), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n865), .A2(G128), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n866), .A2(G137), .ZN(new_n1238));
  INV_X1    g1038(.A(G132), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1237), .B(new_n1238), .C1(new_n788), .C2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1166), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1240), .B1(new_n859), .B2(new_n1241), .ZN(new_n1242));
  OAI221_X1 g1042(.A(new_n1242), .B1(new_n1173), .B2(new_n802), .C1(new_n868), .C2(new_n808), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(new_n1243), .B(KEYINPUT120), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1245), .A2(KEYINPUT59), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n826), .A2(G124), .ZN(new_n1247));
  AOI211_X1 g1047(.A(G33), .B(G41), .C1(new_n979), .C2(G159), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT59), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1247), .B(new_n1248), .C1(new_n1244), .C2(new_n1249), .ZN(new_n1250));
  OAI221_X1 g1050(.A(new_n1236), .B1(KEYINPUT58), .B2(new_n1235), .C1(new_n1246), .C2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1227), .B1(new_n1251), .B2(new_n780), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(new_n1201), .B2(new_n778), .ZN(new_n1253));
  AND2_X1   g1053(.A1(new_n1226), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1225), .A2(new_n1254), .ZN(G375));
  NAND2_X1  g1055(.A1(new_n1126), .A2(new_n777), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n766), .B1(G68), .B2(new_n1162), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT123), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n255), .B1(new_n979), .B2(G77), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n803), .A2(G294), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  OAI221_X1 g1060(.A(new_n1260), .B1(new_n1258), .B2(new_n1259), .C1(new_n384), .C2(new_n808), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n791), .A2(new_n828), .B1(new_n790), .B2(new_n377), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1262), .B1(G116), .B2(new_n787), .ZN(new_n1263));
  OAI221_X1 g1063(.A(new_n1263), .B1(new_n227), .B2(new_n796), .C1(new_n829), .C2(new_n815), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n826), .A2(G128), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n859), .A2(G159), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1232), .B1(new_n787), .B2(new_n1241), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n255), .B1(new_n790), .B2(new_n868), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1268), .B1(G137), .B2(new_n865), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1265), .A2(new_n1266), .A3(new_n1267), .A4(new_n1269), .ZN(new_n1270));
  OAI22_X1  g1070(.A1(new_n802), .A2(new_n1239), .B1(new_n808), .B2(new_n202), .ZN(new_n1271));
  OAI22_X1  g1071(.A1(new_n1261), .A2(new_n1264), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1257), .B1(new_n1272), .B2(new_n780), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(new_n1155), .A2(new_n994), .B1(new_n1256), .B2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1156), .A2(new_n1025), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1150), .A2(new_n1155), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1274), .B1(new_n1275), .B2(new_n1276), .ZN(G381));
  NAND3_X1  g1077(.A1(new_n1087), .A2(new_n841), .A3(new_n1090), .ZN(new_n1278));
  OR4_X1    g1078(.A1(G384), .A2(new_n1278), .A3(G390), .A4(G381), .ZN(new_n1279));
  OR4_X1    g1079(.A1(G387), .A2(new_n1279), .A3(G378), .A4(G375), .ZN(G407));
  INV_X1    g1080(.A(G378), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n698), .A2(G213), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(new_n1282), .B(KEYINPUT124), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1281), .A2(new_n1283), .ZN(new_n1284));
  OAI211_X1 g1084(.A(G407), .B(G213), .C1(G375), .C2(new_n1284), .ZN(G409));
  NAND2_X1  g1085(.A1(G393), .A2(G396), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n1278), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n759), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1044), .B1(new_n1288), .B2(new_n1024), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1041), .ZN(new_n1290));
  AOI21_X1  g1090(.A(G390), .B1(new_n1290), .B2(new_n993), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n993), .ZN(new_n1292));
  AOI211_X1 g1092(.A(new_n1292), .B(new_n1122), .C1(new_n1289), .C2(new_n1041), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1287), .B1(new_n1291), .B2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(G387), .A2(new_n1122), .ZN(new_n1295));
  AND2_X1   g1095(.A1(new_n1286), .A2(new_n1278), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1290), .A2(new_n993), .A3(G390), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1295), .A2(new_n1296), .A3(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1294), .A2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT63), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1225), .A2(G378), .A3(new_n1254), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT125), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1223), .A2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1206), .A2(KEYINPUT125), .A3(new_n1214), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1303), .A2(new_n994), .A3(new_n1304), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1215), .A2(new_n1216), .A3(new_n1025), .A4(new_n1218), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1305), .A2(new_n1253), .A3(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(new_n1281), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1301), .A2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1283), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1276), .A2(KEYINPUT60), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT60), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1312), .B1(new_n1150), .B2(new_n1155), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1311), .A2(new_n1089), .A3(new_n1156), .A4(new_n1313), .ZN(new_n1314));
  AND3_X1   g1114(.A1(new_n1314), .A2(G384), .A3(new_n1274), .ZN(new_n1315));
  AOI21_X1  g1115(.A(G384), .B1(new_n1314), .B2(new_n1274), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1309), .A2(new_n1310), .A3(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1299), .B1(new_n1300), .B2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1283), .A2(G2897), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1321), .ZN(new_n1322));
  XNOR2_X1  g1122(.A(new_n1317), .B(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(KEYINPUT61), .B1(new_n1320), .B2(new_n1323), .ZN(new_n1324));
  OAI211_X1 g1124(.A(new_n1319), .B(new_n1324), .C1(new_n1300), .C2(new_n1318), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1283), .B1(new_n1301), .B2(new_n1308), .ZN(new_n1326));
  AND3_X1   g1126(.A1(new_n1326), .A2(KEYINPUT62), .A3(new_n1317), .ZN(new_n1327));
  AOI21_X1  g1127(.A(KEYINPUT62), .B1(new_n1326), .B2(new_n1317), .ZN(new_n1328));
  OAI211_X1 g1128(.A(new_n1324), .B(KEYINPUT126), .C1(new_n1327), .C2(new_n1328), .ZN(new_n1329));
  AND3_X1   g1129(.A1(new_n1294), .A2(new_n1298), .A3(KEYINPUT127), .ZN(new_n1330));
  AOI21_X1  g1130(.A(KEYINPUT127), .B1(new_n1294), .B2(new_n1298), .ZN(new_n1331));
  NOR2_X1   g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1329), .A2(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT62), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1318), .A2(new_n1334), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1326), .A2(KEYINPUT62), .A3(new_n1317), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  AOI21_X1  g1137(.A(KEYINPUT126), .B1(new_n1337), .B2(new_n1324), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1325), .B1(new_n1333), .B2(new_n1338), .ZN(G405));
  NAND2_X1  g1139(.A1(G375), .A2(new_n1281), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1340), .A2(new_n1301), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1317), .ZN(new_n1342));
  XNOR2_X1  g1142(.A(new_n1341), .B(new_n1342), .ZN(new_n1343));
  XOR2_X1   g1143(.A(new_n1343), .B(new_n1299), .Z(G402));
endmodule


