//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 1 1 0 0 0 0 1 0 1 1 1 0 1 1 0 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 0 1 1 1 0 1 1 1 1 0 1 0 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:33 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G128), .ZN(new_n191));
  AOI21_X1  g005(.A(KEYINPUT73), .B1(new_n191), .B2(G119), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT23), .ZN(new_n193));
  OR2_X1    g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n193), .ZN(new_n195));
  INV_X1    g009(.A(G119), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G128), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n194), .A2(new_n195), .A3(new_n197), .ZN(new_n198));
  XNOR2_X1  g012(.A(G119), .B(G128), .ZN(new_n199));
  XOR2_X1   g013(.A(KEYINPUT24), .B(G110), .Z(new_n200));
  OAI22_X1  g014(.A1(new_n198), .A2(G110), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G125), .ZN(new_n202));
  NOR3_X1   g016(.A1(new_n202), .A2(KEYINPUT16), .A3(G140), .ZN(new_n203));
  XNOR2_X1  g017(.A(G125), .B(G140), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(KEYINPUT16), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G146), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n204), .A2(new_n207), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n201), .A2(new_n206), .A3(new_n208), .ZN(new_n209));
  AOI22_X1  g023(.A1(new_n198), .A2(G110), .B1(new_n199), .B2(new_n200), .ZN(new_n210));
  XNOR2_X1  g024(.A(new_n205), .B(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT22), .B(G137), .ZN(new_n214));
  INV_X1    g028(.A(G953), .ZN(new_n215));
  AND3_X1   g029(.A1(new_n215), .A2(G221), .A3(G234), .ZN(new_n216));
  XOR2_X1   g030(.A(new_n214), .B(new_n216), .Z(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n213), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n209), .A2(new_n212), .A3(new_n217), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(new_n188), .A3(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT25), .ZN(new_n222));
  OR2_X1    g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n222), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n190), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n219), .A2(new_n220), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n189), .A2(G902), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n225), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(G472), .A2(G902), .ZN(new_n232));
  NOR2_X1   g046(.A1(G237), .A2(G953), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G210), .ZN(new_n234));
  XNOR2_X1  g048(.A(new_n234), .B(KEYINPUT27), .ZN(new_n235));
  XNOR2_X1  g049(.A(KEYINPUT26), .B(G101), .ZN(new_n236));
  XNOR2_X1  g050(.A(new_n235), .B(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT11), .ZN(new_n239));
  INV_X1    g053(.A(G134), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n239), .B1(new_n240), .B2(G137), .ZN(new_n241));
  INV_X1    g055(.A(G137), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n242), .A2(KEYINPUT11), .A3(G134), .ZN(new_n243));
  INV_X1    g057(.A(G131), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n240), .A2(G137), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n241), .A2(new_n243), .A3(new_n244), .A4(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G143), .ZN(new_n247));
  OAI21_X1  g061(.A(KEYINPUT1), .B1(new_n247), .B2(G146), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n247), .A2(G146), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n207), .A2(G143), .ZN(new_n250));
  OAI211_X1 g064(.A(G128), .B(new_n248), .C1(new_n249), .C2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n207), .A2(G143), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n247), .A2(G146), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n252), .B(new_n253), .C1(KEYINPUT1), .C2(new_n191), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n240), .A2(G137), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n242), .A2(G134), .ZN(new_n256));
  OAI21_X1  g070(.A(G131), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  AND3_X1   g071(.A1(new_n251), .A2(new_n254), .A3(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n241), .A2(new_n243), .A3(new_n245), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G131), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(new_n246), .ZN(new_n261));
  AND2_X1   g075(.A1(KEYINPUT0), .A2(G128), .ZN(new_n262));
  AND3_X1   g076(.A1(new_n252), .A2(new_n253), .A3(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n262), .B1(new_n252), .B2(new_n253), .ZN(new_n264));
  OAI21_X1  g078(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  NOR3_X1   g080(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n263), .B1(new_n264), .B2(new_n268), .ZN(new_n269));
  AOI22_X1  g083(.A1(new_n246), .A2(new_n258), .B1(new_n261), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G116), .ZN(new_n271));
  OAI21_X1  g085(.A(KEYINPUT65), .B1(new_n271), .B2(G119), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT65), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n273), .A2(new_n196), .A3(G116), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g089(.A(KEYINPUT66), .B(G116), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G119), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g092(.A(KEYINPUT2), .B(G113), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n279), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n281), .B1(new_n275), .B2(new_n277), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n238), .B1(new_n270), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT67), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n258), .A2(new_n285), .A3(new_n246), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n261), .A2(new_n269), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n251), .A2(new_n246), .A3(new_n257), .A4(new_n254), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(KEYINPUT67), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n283), .A2(new_n286), .A3(new_n287), .A4(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n287), .A2(new_n288), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n272), .A2(new_n274), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n292), .B1(G119), .B2(new_n276), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n281), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n278), .A2(new_n279), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n291), .A2(KEYINPUT68), .A3(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n284), .A2(new_n290), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT28), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT69), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n270), .A2(new_n283), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT28), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n299), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n298), .A2(KEYINPUT69), .A3(KEYINPUT28), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n237), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT30), .ZN(new_n308));
  AND3_X1   g122(.A1(new_n287), .A2(new_n308), .A3(new_n288), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n286), .A2(new_n287), .A3(new_n289), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n309), .B1(KEYINPUT30), .B2(new_n310), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n237), .B(new_n290), .C1(new_n311), .C2(new_n283), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(KEYINPUT31), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n260), .A2(new_n246), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n268), .A2(new_n264), .ZN(new_n315));
  INV_X1    g129(.A(new_n263), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  OAI22_X1  g131(.A1(new_n314), .A2(new_n317), .B1(KEYINPUT67), .B2(new_n288), .ZN(new_n318));
  INV_X1    g132(.A(new_n289), .ZN(new_n319));
  OAI21_X1  g133(.A(KEYINPUT30), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n309), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n296), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT31), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n323), .A2(new_n324), .A3(new_n237), .A4(new_n290), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n313), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n232), .B1(new_n307), .B2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT70), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT32), .ZN(new_n330));
  OAI211_X1 g144(.A(KEYINPUT70), .B(new_n232), .C1(new_n307), .C2(new_n326), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n232), .ZN(new_n333));
  INV_X1    g147(.A(new_n326), .ZN(new_n334));
  INV_X1    g148(.A(new_n237), .ZN(new_n335));
  AND3_X1   g149(.A1(new_n298), .A2(KEYINPUT69), .A3(KEYINPUT28), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n303), .B1(new_n298), .B2(KEYINPUT28), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n335), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n333), .B1(new_n334), .B2(new_n338), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n318), .A2(new_n319), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT71), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(new_n341), .A3(new_n283), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n290), .A2(KEYINPUT71), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n310), .A2(new_n296), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(KEYINPUT28), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n301), .A2(new_n302), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n346), .A2(KEYINPUT29), .A3(new_n237), .A4(new_n347), .ZN(new_n348));
  NOR3_X1   g162(.A1(new_n336), .A2(new_n337), .A3(new_n335), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT29), .ZN(new_n350));
  INV_X1    g164(.A(new_n290), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n351), .B1(new_n322), .B2(new_n296), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n350), .B1(new_n352), .B2(new_n237), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n348), .B(new_n188), .C1(new_n349), .C2(new_n353), .ZN(new_n354));
  AOI22_X1  g168(.A1(new_n339), .A2(KEYINPUT32), .B1(new_n354), .B2(G472), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n332), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT72), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n332), .A2(new_n355), .A3(KEYINPUT72), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n231), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(G469), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n215), .A2(G227), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n362), .B(KEYINPUT74), .ZN(new_n363));
  XNOR2_X1  g177(.A(G110), .B(G140), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n363), .B(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT79), .ZN(new_n367));
  NAND2_X1  g181(.A1(KEYINPUT75), .A2(G104), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(KEYINPUT3), .A2(G107), .ZN(new_n370));
  NOR2_X1   g184(.A1(KEYINPUT75), .A2(G104), .ZN(new_n371));
  NOR3_X1   g185(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT3), .ZN(new_n373));
  INV_X1    g187(.A(G107), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(new_n374), .A3(G104), .ZN(new_n375));
  NAND2_X1  g189(.A1(KEYINPUT3), .A2(G107), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(KEYINPUT76), .B1(new_n372), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT4), .ZN(new_n379));
  AND2_X1   g193(.A1(KEYINPUT3), .A2(G107), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n380), .B1(G104), .B2(new_n370), .ZN(new_n381));
  OR2_X1    g195(.A1(KEYINPUT75), .A2(G104), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n373), .A2(new_n374), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n382), .A2(new_n383), .A3(new_n368), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT76), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n381), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n378), .A2(new_n379), .A3(G101), .A4(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(KEYINPUT77), .ZN(new_n388));
  INV_X1    g202(.A(G101), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n381), .A2(new_n384), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n389), .B1(new_n390), .B2(KEYINPUT76), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT77), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n391), .A2(new_n392), .A3(new_n379), .A4(new_n386), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n388), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n378), .A2(G101), .A3(new_n386), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n381), .A2(new_n384), .A3(new_n389), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n396), .A2(KEYINPUT4), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n317), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  AND2_X1   g212(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n382), .A2(new_n374), .A3(new_n368), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n389), .B1(G104), .B2(G107), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n396), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n251), .A2(new_n254), .ZN(new_n404));
  NOR3_X1   g218(.A1(new_n403), .A2(KEYINPUT10), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(KEYINPUT78), .ZN(new_n406));
  INV_X1    g220(.A(new_n404), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT78), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n396), .A2(new_n408), .A3(new_n402), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n406), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n405), .B1(new_n410), .B2(KEYINPUT10), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n367), .B1(new_n399), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n410), .A2(KEYINPUT10), .ZN(new_n413));
  INV_X1    g227(.A(new_n405), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n394), .A2(new_n398), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n415), .A2(KEYINPUT79), .A3(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n412), .A2(new_n261), .A3(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n415), .A2(new_n314), .A3(new_n416), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n366), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n403), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n421), .A2(new_n407), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n403), .A2(new_n404), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n261), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT12), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  OAI211_X1 g240(.A(KEYINPUT12), .B(new_n261), .C1(new_n422), .C2(new_n423), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AND3_X1   g242(.A1(new_n419), .A2(new_n428), .A3(new_n366), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n361), .B(new_n188), .C1(new_n420), .C2(new_n429), .ZN(new_n430));
  AOI22_X1  g244(.A1(new_n413), .A2(new_n414), .B1(new_n394), .B2(new_n398), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n365), .B1(new_n431), .B2(new_n314), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n261), .B1(new_n431), .B2(KEYINPUT79), .ZN(new_n433));
  INV_X1    g247(.A(new_n417), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n419), .A2(new_n428), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n365), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n435), .A2(G469), .A3(new_n437), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n361), .A2(new_n188), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n430), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(G221), .ZN(new_n442));
  XNOR2_X1  g256(.A(KEYINPUT9), .B(G234), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n442), .B1(new_n444), .B2(new_n188), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n441), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(G214), .B1(G237), .B2(G902), .ZN(new_n448));
  XNOR2_X1  g262(.A(G110), .B(G122), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT80), .ZN(new_n451));
  AOI22_X1  g265(.A1(new_n395), .A2(new_n397), .B1(new_n294), .B2(new_n295), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n394), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n293), .A2(KEYINPUT5), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n196), .A2(G116), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n454), .B(G113), .C1(KEYINPUT5), .C2(new_n455), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n456), .A2(new_n294), .A3(new_n406), .A4(new_n409), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n451), .B1(new_n394), .B2(new_n452), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n450), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n394), .A2(new_n452), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(KEYINPUT80), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n462), .A2(new_n449), .A3(new_n457), .A4(new_n453), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n460), .A2(KEYINPUT6), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n269), .A2(G125), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n465), .B1(G125), .B2(new_n404), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n215), .A2(G224), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n467), .B(KEYINPUT81), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n466), .B(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT6), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n470), .B(new_n450), .C1(new_n458), .C2(new_n459), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n464), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n467), .A2(KEYINPUT7), .ZN(new_n473));
  XOR2_X1   g287(.A(new_n466), .B(new_n473), .Z(new_n474));
  NAND3_X1  g288(.A1(new_n456), .A2(new_n294), .A3(new_n403), .ZN(new_n475));
  XOR2_X1   g289(.A(new_n449), .B(KEYINPUT8), .Z(new_n476));
  NAND2_X1  g290(.A1(new_n456), .A2(new_n294), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n476), .B1(new_n477), .B2(new_n421), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n474), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(G902), .B1(new_n479), .B2(new_n463), .ZN(new_n480));
  OAI21_X1  g294(.A(G210), .B1(G237), .B2(G902), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n472), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n481), .B1(new_n472), .B2(new_n480), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n448), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n447), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT86), .ZN(new_n486));
  AOI21_X1  g300(.A(G143), .B1(new_n233), .B2(G214), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n233), .A2(G143), .A3(G214), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n490), .A2(KEYINPUT18), .A3(G131), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n204), .B(new_n207), .ZN(new_n492));
  NAND2_X1  g306(.A1(KEYINPUT18), .A2(G131), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n488), .A2(new_n489), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n491), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n205), .B(new_n207), .ZN(new_n497));
  INV_X1    g311(.A(new_n489), .ZN(new_n498));
  OAI21_X1  g312(.A(G131), .B1(new_n498), .B2(new_n487), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n488), .A2(new_n244), .A3(new_n489), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT85), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT17), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n499), .A2(new_n500), .A3(new_n501), .A4(new_n502), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n497), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(KEYINPUT84), .B1(new_n499), .B2(new_n502), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT84), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n490), .A2(new_n506), .A3(KEYINPUT17), .A4(G131), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n499), .A2(new_n500), .A3(new_n502), .ZN(new_n508));
  AOI22_X1  g322(.A1(new_n505), .A2(new_n507), .B1(new_n508), .B2(KEYINPUT85), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n496), .B1(new_n504), .B2(new_n509), .ZN(new_n510));
  XNOR2_X1  g324(.A(G113), .B(G122), .ZN(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT83), .B(G104), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n511), .B(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n486), .B1(new_n510), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n505), .A2(new_n507), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n508), .A2(KEYINPUT85), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n515), .A2(new_n516), .A3(new_n497), .A4(new_n503), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n517), .A2(new_n495), .A3(new_n513), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n518), .A2(KEYINPUT86), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n499), .A2(new_n500), .ZN(new_n520));
  XOR2_X1   g334(.A(new_n204), .B(KEYINPUT19), .Z(new_n521));
  OAI211_X1 g335(.A(new_n520), .B(new_n206), .C1(new_n521), .C2(G146), .ZN(new_n522));
  AND2_X1   g336(.A1(new_n522), .A2(new_n495), .ZN(new_n523));
  OAI22_X1  g337(.A1(new_n514), .A2(new_n519), .B1(new_n523), .B2(new_n513), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT20), .ZN(new_n525));
  NOR2_X1   g339(.A1(G475), .A2(G902), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  XOR2_X1   g341(.A(KEYINPUT82), .B(KEYINPUT20), .Z(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n523), .A2(new_n513), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n510), .A2(new_n486), .A3(new_n513), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n518), .A2(KEYINPUT86), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n526), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n529), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n527), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n514), .A2(new_n519), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT88), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n538), .B1(new_n510), .B2(new_n513), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n517), .A2(new_n495), .ZN(new_n540));
  INV_X1    g354(.A(new_n513), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n540), .A2(KEYINPUT88), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n188), .B1(new_n537), .B2(new_n543), .ZN(new_n544));
  XOR2_X1   g358(.A(KEYINPUT87), .B(G475), .Z(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n536), .A2(new_n546), .ZN(new_n547));
  NOR3_X1   g361(.A1(new_n443), .A2(new_n187), .A3(G953), .ZN(new_n548));
  XNOR2_X1  g362(.A(G128), .B(G143), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n549), .B(new_n240), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n276), .A2(G122), .ZN(new_n551));
  OR2_X1    g365(.A1(new_n271), .A2(G122), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(new_n374), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT14), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n551), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT90), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n374), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n557), .B(KEYINPUT90), .C1(KEYINPUT14), .C2(new_n551), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n554), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT89), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT13), .ZN(new_n565));
  AOI22_X1  g379(.A1(new_n564), .A2(new_n565), .B1(new_n191), .B2(G143), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n566), .B1(new_n564), .B2(new_n565), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(G134), .ZN(new_n568));
  INV_X1    g382(.A(new_n549), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n567), .A2(G134), .A3(new_n549), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n551), .A2(new_n552), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(G107), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n553), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n548), .B1(new_n563), .B2(new_n576), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n572), .A2(new_n575), .ZN(new_n578));
  INV_X1    g392(.A(new_n548), .ZN(new_n579));
  NOR3_X1   g393(.A1(new_n578), .A2(new_n562), .A3(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n188), .B1(new_n577), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(G478), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n582), .A2(KEYINPUT15), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  OAI221_X1 g398(.A(new_n188), .B1(KEYINPUT15), .B2(new_n582), .C1(new_n577), .C2(new_n580), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(G952), .ZN(new_n587));
  AOI211_X1 g401(.A(G953), .B(new_n587), .C1(G234), .C2(G237), .ZN(new_n588));
  XNOR2_X1  g402(.A(KEYINPUT21), .B(G898), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(KEYINPUT91), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  AOI211_X1 g405(.A(new_n188), .B(new_n215), .C1(G234), .C2(G237), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n588), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NOR3_X1   g407(.A1(new_n547), .A2(new_n586), .A3(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n360), .A2(new_n485), .A3(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(G101), .ZN(G3));
  OAI21_X1  g410(.A(new_n188), .B1(new_n307), .B2(new_n326), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(G472), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n329), .A2(new_n598), .A3(new_n331), .A4(new_n230), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n447), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(KEYINPUT92), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n472), .A2(new_n480), .ZN(new_n602));
  INV_X1    g416(.A(new_n481), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n472), .A2(new_n480), .A3(new_n481), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n593), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n606), .A2(new_n448), .A3(new_n607), .ZN(new_n608));
  OR2_X1    g422(.A1(new_n577), .A2(new_n580), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT33), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n582), .A2(G902), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n581), .ZN(new_n614));
  XOR2_X1   g428(.A(KEYINPUT93), .B(G478), .Z(new_n615));
  OAI22_X1  g429(.A1(new_n611), .A2(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n547), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n608), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n601), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT34), .B(G104), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G6));
  AND2_X1   g435(.A1(new_n546), .A2(new_n586), .ZN(new_n622));
  OR4_X1    g436(.A1(KEYINPUT94), .A2(new_n533), .A3(new_n529), .A4(new_n534), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n524), .A2(new_n528), .A3(new_n526), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n624), .A2(new_n535), .A3(KEYINPUT94), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n622), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n608), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n601), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT35), .B(G107), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G9));
  AND3_X1   g444(.A1(new_n329), .A2(new_n598), .A3(new_n331), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n218), .A2(KEYINPUT36), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n213), .B(new_n632), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n633), .A2(new_n227), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n225), .A2(new_n634), .ZN(new_n635));
  NOR4_X1   g449(.A1(new_n547), .A2(new_n635), .A3(new_n586), .A4(new_n593), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n485), .A2(new_n631), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(KEYINPUT37), .B(G110), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(KEYINPUT95), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n637), .B(new_n639), .ZN(G12));
  NOR2_X1   g454(.A1(new_n447), .A2(new_n635), .ZN(new_n641));
  INV_X1    g455(.A(G900), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n592), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n588), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n622), .A2(new_n623), .A3(new_n625), .A4(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n646), .A2(new_n484), .ZN(new_n647));
  AND3_X1   g461(.A1(new_n332), .A2(new_n355), .A3(KEYINPUT72), .ZN(new_n648));
  AOI21_X1  g462(.A(KEYINPUT72), .B1(new_n332), .B2(new_n355), .ZN(new_n649));
  OAI211_X1 g463(.A(new_n641), .B(new_n647), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(G128), .ZN(G30));
  OR2_X1    g465(.A1(new_n352), .A2(new_n335), .ZN(new_n652));
  OAI211_X1 g466(.A(new_n652), .B(new_n188), .C1(new_n237), .C2(new_n345), .ZN(new_n653));
  AOI22_X1  g467(.A1(new_n339), .A2(KEYINPUT32), .B1(G472), .B2(new_n653), .ZN(new_n654));
  AND3_X1   g468(.A1(new_n332), .A2(new_n654), .A3(KEYINPUT96), .ZN(new_n655));
  AOI21_X1  g469(.A(KEYINPUT96), .B1(new_n332), .B2(new_n654), .ZN(new_n656));
  OR2_X1    g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n606), .B(KEYINPUT38), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n586), .A2(new_n448), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n659), .B1(new_n536), .B2(new_n546), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n657), .A2(new_n635), .A3(new_n658), .A4(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n645), .B(KEYINPUT39), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n441), .A2(new_n446), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT40), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(new_n247), .ZN(G45));
  NAND3_X1  g480(.A1(new_n616), .A2(new_n547), .A3(new_n645), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n484), .A2(new_n667), .ZN(new_n668));
  OAI211_X1 g482(.A(new_n641), .B(new_n668), .C1(new_n648), .C2(new_n649), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT97), .B(G146), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G48));
  OAI21_X1  g485(.A(new_n419), .B1(new_n433), .B2(new_n434), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n429), .B1(new_n672), .B2(new_n365), .ZN(new_n673));
  OAI21_X1  g487(.A(G469), .B1(new_n673), .B2(G902), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n674), .A2(new_n446), .A3(new_n430), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT98), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n674), .A2(KEYINPUT98), .A3(new_n446), .A4(new_n430), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT99), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n677), .A2(KEYINPUT99), .A3(new_n678), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n360), .A2(new_n618), .A3(new_n681), .A4(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(KEYINPUT41), .B(G113), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G15));
  NAND4_X1  g499(.A1(new_n360), .A2(new_n627), .A3(new_n681), .A4(new_n682), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G116), .ZN(G18));
  NAND2_X1  g501(.A1(new_n358), .A2(new_n359), .ZN(new_n688));
  INV_X1    g502(.A(new_n448), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n689), .B1(new_n604), .B2(new_n605), .ZN(new_n690));
  AND3_X1   g504(.A1(new_n677), .A2(new_n690), .A3(new_n678), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n688), .A2(new_n691), .A3(new_n636), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G119), .ZN(G21));
  AOI21_X1  g507(.A(new_n237), .B1(new_n346), .B2(new_n347), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n232), .B1(new_n694), .B2(new_n326), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT100), .ZN(new_n696));
  AND3_X1   g510(.A1(new_n597), .A2(new_n696), .A3(G472), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n696), .B1(new_n597), .B2(G472), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n230), .B(new_n695), .C1(new_n697), .C2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n606), .A2(new_n660), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n699), .A2(new_n700), .A3(new_n593), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n681), .A2(new_n701), .A3(new_n682), .ZN(new_n702));
  XNOR2_X1  g516(.A(KEYINPUT101), .B(G122), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G24));
  INV_X1    g518(.A(new_n635), .ZN(new_n705));
  OAI211_X1 g519(.A(new_n705), .B(new_n695), .C1(new_n697), .C2(new_n698), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n706), .A2(new_n667), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n691), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G125), .ZN(G27));
  NOR2_X1   g523(.A1(new_n482), .A2(new_n483), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n445), .A2(new_n689), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT102), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n438), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n435), .A2(KEYINPUT102), .A3(G469), .A4(new_n437), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n716), .A2(KEYINPUT103), .A3(new_n430), .A4(new_n440), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n430), .A2(new_n714), .A3(new_n440), .A4(new_n715), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT103), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n712), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n667), .A2(KEYINPUT42), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n688), .A2(new_n721), .A3(new_n230), .A4(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n711), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n606), .A2(new_n724), .ZN(new_n725));
  AND2_X1   g539(.A1(new_n718), .A2(new_n719), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n718), .A2(new_n719), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n355), .B1(KEYINPUT32), .B2(new_n339), .ZN(new_n729));
  INV_X1    g543(.A(new_n667), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n729), .A2(new_n230), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g545(.A(KEYINPUT42), .B1(new_n728), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n723), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(new_n244), .ZN(G33));
  INV_X1    g548(.A(new_n646), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n360), .A2(new_n735), .A3(new_n721), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G134), .ZN(G36));
  AND2_X1   g551(.A1(new_n536), .A2(new_n546), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n616), .ZN(new_n739));
  XOR2_X1   g553(.A(new_n739), .B(KEYINPUT43), .Z(new_n740));
  INV_X1    g554(.A(new_n631), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n740), .A2(new_n741), .A3(new_n705), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT44), .ZN(new_n743));
  OR2_X1    g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n435), .A2(new_n437), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT45), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n435), .A2(KEYINPUT45), .A3(new_n437), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n747), .A2(G469), .A3(new_n748), .ZN(new_n749));
  AOI21_X1  g563(.A(KEYINPUT46), .B1(new_n749), .B2(new_n440), .ZN(new_n750));
  INV_X1    g564(.A(new_n430), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n749), .A2(KEYINPUT46), .A3(new_n440), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n445), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n754), .A2(new_n662), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n742), .A2(new_n743), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n710), .A2(new_n448), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n744), .A2(new_n755), .A3(new_n756), .A4(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(KEYINPUT104), .B(G137), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n759), .B(new_n760), .ZN(G39));
  NAND2_X1  g575(.A1(KEYINPUT105), .A2(KEYINPUT47), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n754), .A2(new_n762), .ZN(new_n763));
  XOR2_X1   g577(.A(KEYINPUT105), .B(KEYINPUT47), .Z(new_n764));
  OAI21_X1  g578(.A(new_n763), .B1(new_n754), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n758), .A2(new_n231), .A3(new_n730), .ZN(new_n766));
  OR2_X1    g580(.A1(new_n766), .A2(new_n688), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  XOR2_X1   g582(.A(new_n768), .B(KEYINPUT106), .Z(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G140), .ZN(G42));
  NAND2_X1  g584(.A1(new_n587), .A2(new_n215), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(KEYINPUT117), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT51), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n740), .A2(new_n588), .ZN(new_n774));
  INV_X1    g588(.A(new_n699), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n658), .A2(new_n679), .A3(new_n448), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  XOR2_X1   g592(.A(new_n778), .B(KEYINPUT50), .Z(new_n779));
  NOR2_X1   g593(.A1(new_n679), .A2(new_n757), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n774), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n781), .A2(new_n706), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(KEYINPUT115), .ZN(new_n783));
  INV_X1    g597(.A(new_n780), .ZN(new_n784));
  NOR4_X1   g598(.A1(new_n784), .A2(new_n657), .A3(new_n231), .A4(new_n644), .ZN(new_n785));
  INV_X1    g599(.A(new_n616), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n785), .A2(new_n738), .A3(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n779), .A2(new_n783), .A3(new_n787), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n776), .A2(new_n758), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n674), .A2(new_n430), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n790), .A2(KEYINPUT114), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(KEYINPUT114), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n791), .A2(new_n445), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n765), .A2(new_n793), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n789), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n773), .B1(new_n788), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n729), .A2(new_n230), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n781), .A2(new_n797), .ZN(new_n798));
  XOR2_X1   g612(.A(new_n798), .B(KEYINPUT48), .Z(new_n799));
  NAND3_X1  g613(.A1(new_n785), .A2(new_n547), .A3(new_n616), .ZN(new_n800));
  AOI211_X1 g614(.A(new_n587), .B(G953), .C1(new_n776), .C2(new_n691), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n788), .A2(new_n773), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT116), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n789), .B1(new_n794), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n805), .B1(new_n804), .B2(new_n794), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n796), .B(new_n802), .C1(new_n803), .C2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n645), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n808), .A2(new_n445), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n606), .A2(new_n635), .A3(new_n660), .A4(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n717), .A2(new_n720), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n811), .B(new_n812), .C1(new_n656), .C2(new_n655), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n708), .A2(new_n813), .A3(new_n650), .A4(new_n669), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT52), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n708), .A2(new_n650), .A3(new_n669), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n813), .A2(KEYINPUT52), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT111), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n708), .A2(new_n650), .A3(new_n669), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n813), .A2(KEYINPUT52), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT111), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n816), .B1(new_n819), .B2(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n683), .A2(new_n686), .A3(new_n692), .A4(new_n702), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(KEYINPUT112), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n702), .A2(new_n692), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT112), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n827), .A2(new_n828), .A3(new_n683), .A4(new_n686), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n536), .A2(new_n546), .A3(new_n586), .A4(new_n607), .ZN(new_n831));
  OAI21_X1  g645(.A(KEYINPUT109), .B1(new_n484), .B2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT109), .ZN(new_n833));
  INV_X1    g647(.A(new_n831), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n690), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n600), .A2(new_n832), .A3(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n836), .A2(new_n637), .A3(KEYINPUT110), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n723), .A2(new_n732), .A3(KEYINPUT53), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n230), .B1(new_n648), .B2(new_n649), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n839), .A2(new_n728), .A3(new_n646), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n721), .A2(new_n707), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n586), .A2(new_n808), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n623), .A2(new_n625), .A3(new_n546), .A4(new_n842), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n606), .A2(new_n843), .A3(new_n689), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n641), .B(new_n844), .C1(new_n648), .C2(new_n649), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n841), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n840), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n618), .A2(new_n600), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n485), .A2(new_n594), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n848), .B1(new_n839), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(KEYINPUT110), .B1(new_n836), .B2(new_n637), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AND4_X1   g666(.A1(new_n837), .A2(new_n838), .A3(new_n847), .A4(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n824), .A2(new_n830), .A3(new_n853), .A4(KEYINPUT113), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n817), .A2(new_n818), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n816), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n836), .A2(new_n637), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT110), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n859), .A2(new_n595), .A3(new_n837), .A4(new_n848), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n825), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n736), .A2(new_n841), .A3(new_n845), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n863), .A2(new_n733), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n856), .A2(new_n861), .A3(new_n862), .A4(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT53), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n854), .A2(new_n867), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n838), .A2(new_n847), .A3(new_n852), .A4(new_n837), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n869), .B1(new_n826), .B2(new_n829), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT113), .B1(new_n870), .B2(new_n824), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT54), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n861), .A2(new_n862), .ZN(new_n875));
  NOR4_X1   g689(.A1(new_n875), .A2(KEYINPUT53), .A3(new_n733), .A4(new_n863), .ZN(new_n876));
  AOI22_X1  g690(.A1(new_n876), .A2(new_n824), .B1(KEYINPUT53), .B2(new_n865), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(KEYINPUT54), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n772), .B1(new_n807), .B2(new_n879), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n739), .A2(new_n231), .A3(new_n724), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT107), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT49), .ZN(new_n883));
  INV_X1    g697(.A(new_n790), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n883), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT108), .ZN(new_n887));
  OR3_X1    g701(.A1(new_n885), .A2(new_n658), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n880), .B1(new_n657), .B2(new_n888), .ZN(G75));
  OAI211_X1 g703(.A(G210), .B(G902), .C1(new_n868), .C2(new_n871), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT56), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n464), .A2(new_n471), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(new_n469), .ZN(new_n894));
  XNOR2_X1  g708(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n894), .B(new_n895), .Z(new_n896));
  NAND2_X1  g710(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(new_n896), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n890), .A2(new_n891), .A3(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n215), .A2(G952), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n897), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT119), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n897), .A2(KEYINPUT119), .A3(new_n899), .A4(new_n901), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(G51));
  XNOR2_X1  g720(.A(new_n872), .B(KEYINPUT54), .ZN(new_n907));
  XNOR2_X1  g721(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n440), .B(new_n908), .ZN(new_n909));
  OAI22_X1  g723(.A1(new_n907), .A2(new_n909), .B1(new_n420), .B2(new_n429), .ZN(new_n910));
  OR3_X1    g724(.A1(new_n872), .A2(new_n188), .A3(new_n749), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n900), .B1(new_n910), .B2(new_n911), .ZN(G54));
  INV_X1    g726(.A(KEYINPUT121), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n872), .A2(new_n188), .ZN(new_n914));
  AND2_X1   g728(.A1(KEYINPUT58), .A2(G475), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n913), .B1(new_n916), .B2(new_n533), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n900), .B1(new_n916), .B2(new_n533), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n914), .A2(KEYINPUT121), .A3(new_n524), .A4(new_n915), .ZN(new_n919));
  AND3_X1   g733(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(G60));
  INV_X1    g734(.A(new_n611), .ZN(new_n921));
  NAND2_X1  g735(.A1(G478), .A2(G902), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n922), .B(KEYINPUT59), .Z(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n901), .B1(new_n907), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n921), .B1(new_n879), .B2(new_n924), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n926), .A2(new_n927), .ZN(G63));
  NAND2_X1  g742(.A1(G217), .A2(G902), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT122), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT60), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n931), .B1(new_n868), .B2(new_n871), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n900), .B1(new_n932), .B2(new_n226), .ZN(new_n933));
  OAI211_X1 g747(.A(new_n633), .B(new_n931), .C1(new_n868), .C2(new_n871), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT123), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT61), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n935), .A2(new_n936), .A3(new_n939), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n933), .A2(new_n937), .A3(new_n938), .A4(new_n934), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n940), .A2(new_n941), .ZN(G66));
  AOI21_X1  g756(.A(new_n215), .B1(new_n590), .B2(G224), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n943), .B1(new_n875), .B2(new_n215), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n893), .B1(G898), .B2(new_n215), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n944), .B(new_n945), .Z(G69));
  NAND2_X1  g760(.A1(G900), .A2(G953), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n797), .A2(new_n700), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n840), .B1(new_n755), .B2(new_n948), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n733), .A2(new_n820), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n769), .A2(new_n759), .A3(new_n949), .A4(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n947), .B1(new_n951), .B2(G953), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n311), .B(new_n521), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(KEYINPUT62), .B1(new_n665), .B2(new_n820), .ZN(new_n955));
  OR3_X1    g769(.A1(new_n665), .A2(KEYINPUT62), .A3(new_n820), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n738), .A2(new_n586), .ZN(new_n957));
  AOI211_X1 g771(.A(new_n663), .B(new_n757), .C1(new_n617), .C2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n360), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n759), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n769), .A2(new_n955), .A3(new_n956), .A4(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n953), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n961), .A2(new_n215), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n954), .A2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(G227), .ZN(new_n965));
  OAI21_X1  g779(.A(G953), .B1(new_n965), .B2(new_n642), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT124), .Z(new_n967));
  XNOR2_X1  g781(.A(new_n964), .B(new_n967), .ZN(G72));
  NAND2_X1  g782(.A1(new_n352), .A2(new_n335), .ZN(new_n969));
  XOR2_X1   g783(.A(KEYINPUT125), .B(KEYINPUT63), .Z(new_n970));
  NAND2_X1  g784(.A1(G472), .A2(G902), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n970), .B(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n652), .A2(new_n969), .A3(new_n972), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT126), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n877), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT127), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n972), .B1(new_n961), .B2(new_n875), .ZN(new_n977));
  INV_X1    g791(.A(new_n652), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n972), .B1(new_n951), .B2(new_n875), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n980), .A2(new_n335), .A3(new_n352), .ZN(new_n981));
  AND4_X1   g795(.A1(new_n901), .A2(new_n976), .A3(new_n979), .A4(new_n981), .ZN(G57));
endmodule


