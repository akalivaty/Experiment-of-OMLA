//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0 1 1 0 1 0 1 1 0 0 1 0 0 1 1 0 1 1 0 1 0 1 1 0 1 1 1 1 0 0 0 1 0 1 0 0 1 0 1 1 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n851, new_n852, new_n853, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961;
  INV_X1    g000(.A(KEYINPUT15), .ZN(new_n202));
  XNOR2_X1  g001(.A(G43gat), .B(G50gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT82), .ZN(new_n204));
  AOI21_X1  g003(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(new_n204), .B2(new_n203), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT14), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n207), .B1(G29gat), .B2(G36gat), .ZN(new_n208));
  OR3_X1    g007(.A1(new_n207), .A2(G29gat), .A3(G36gat), .ZN(new_n209));
  XOR2_X1   g008(.A(KEYINPUT83), .B(G36gat), .Z(new_n210));
  INV_X1    g009(.A(G29gat), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n208), .B(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  OR2_X1    g011(.A1(new_n206), .A2(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n203), .A2(KEYINPUT15), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n206), .B1(new_n214), .B2(new_n212), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G15gat), .B(G22gat), .ZN(new_n217));
  OR2_X1    g016(.A1(new_n217), .A2(KEYINPUT85), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(KEYINPUT85), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT16), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n220), .B1(new_n221), .B2(G1gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT86), .ZN(new_n223));
  INV_X1    g022(.A(G1gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n218), .A2(new_n224), .A3(new_n219), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n222), .A2(new_n223), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(G8gat), .ZN(new_n227));
  INV_X1    g026(.A(G8gat), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n222), .A2(new_n223), .A3(new_n225), .A4(new_n228), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n216), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n227), .A2(new_n229), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT17), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n233), .B1(new_n216), .B2(KEYINPUT84), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT84), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n213), .A2(new_n235), .A3(KEYINPUT17), .A4(new_n215), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n230), .B1(new_n232), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(G229gat), .A2(G233gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT87), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n241), .A2(KEYINPUT18), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n232), .A2(new_n216), .ZN(new_n244));
  INV_X1    g043(.A(new_n230), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XOR2_X1   g045(.A(new_n239), .B(KEYINPUT13), .Z(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n238), .B(new_n239), .C1(new_n241), .C2(KEYINPUT18), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n243), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(G113gat), .B(G141gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n251), .B(G197gat), .ZN(new_n252));
  XOR2_X1   g051(.A(KEYINPUT11), .B(G169gat), .Z(new_n253));
  XNOR2_X1  g052(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n255));
  XOR2_X1   g054(.A(new_n254), .B(new_n255), .Z(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n250), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n243), .A2(new_n256), .A3(new_n249), .A4(new_n248), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(G134gat), .B(G162gat), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n263));
  XOR2_X1   g062(.A(new_n262), .B(new_n263), .Z(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G99gat), .B(G106gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(G85gat), .A2(G92gat), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT90), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT7), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(G85gat), .ZN(new_n271));
  INV_X1    g070(.A(G92gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(G99gat), .A2(G106gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT8), .ZN(new_n275));
  AND3_X1   g074(.A1(new_n270), .A2(new_n273), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n267), .A2(new_n268), .ZN(new_n277));
  NAND3_X1  g076(.A1(KEYINPUT90), .A2(G85gat), .A3(G92gat), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n277), .A2(KEYINPUT7), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n266), .B1(new_n276), .B2(new_n279), .ZN(new_n280));
  AOI22_X1  g079(.A1(KEYINPUT8), .A2(new_n274), .B1(new_n271), .B2(new_n272), .ZN(new_n281));
  AND4_X1   g080(.A1(new_n266), .A2(new_n279), .A3(new_n270), .A4(new_n281), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n213), .A2(new_n215), .A3(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT91), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n284), .A2(KEYINPUT91), .A3(new_n285), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n283), .B1(new_n234), .B2(new_n236), .ZN(new_n292));
  XNOR2_X1  g091(.A(G190gat), .B(G218gat), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  NOR3_X1   g093(.A1(new_n291), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n292), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n293), .B1(new_n296), .B2(new_n290), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n265), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT93), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OAI211_X1 g099(.A(KEYINPUT93), .B(new_n265), .C1(new_n295), .C2(new_n297), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n294), .B1(new_n291), .B2(new_n292), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n296), .A2(new_n290), .A3(new_n293), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n303), .A2(new_n264), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT92), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND4_X1  g106(.A1(new_n303), .A2(KEYINPUT92), .A3(new_n264), .A4(new_n304), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AND2_X1   g108(.A1(new_n302), .A2(new_n309), .ZN(new_n310));
  AND2_X1   g109(.A1(G71gat), .A2(G78gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(G71gat), .A2(G78gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(G57gat), .B(G64gat), .ZN(new_n314));
  AOI21_X1  g113(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n313), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(G57gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G64gat), .ZN(new_n318));
  INV_X1    g117(.A(G64gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G57gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(G71gat), .B(G78gat), .ZN(new_n322));
  INV_X1    g121(.A(new_n315), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  AND3_X1   g123(.A1(new_n316), .A2(new_n324), .A3(KEYINPUT89), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT89), .B1(new_n316), .B2(new_n324), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n231), .B1(KEYINPUT21), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n316), .A2(new_n324), .ZN(new_n329));
  XOR2_X1   g128(.A(KEYINPUT88), .B(KEYINPUT21), .Z(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(G231gat), .A2(G233gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n333), .B(G127gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n328), .B(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n336), .B(G155gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(G183gat), .B(G211gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n337), .B(new_n338), .ZN(new_n339));
  OR2_X1    g138(.A1(new_n335), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n335), .A2(new_n339), .ZN(new_n341));
  AND2_X1   g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  AND2_X1   g142(.A1(new_n316), .A2(new_n324), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n344), .B1(new_n280), .B2(new_n282), .ZN(new_n345));
  INV_X1    g144(.A(new_n266), .ZN(new_n346));
  INV_X1    g145(.A(new_n279), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n281), .A2(new_n270), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n346), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n276), .A2(new_n266), .A3(new_n279), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n349), .A2(new_n329), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(KEYINPUT10), .B1(new_n345), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT94), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT10), .ZN(new_n355));
  NOR3_X1   g154(.A1(new_n325), .A2(new_n326), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n354), .B1(new_n356), .B2(new_n283), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT89), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n329), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n316), .A2(new_n324), .A3(KEYINPUT89), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n359), .A2(KEYINPUT10), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n349), .A2(new_n350), .ZN(new_n362));
  NOR3_X1   g161(.A1(new_n361), .A2(KEYINPUT94), .A3(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n353), .B1(new_n357), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(G230gat), .A2(G233gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n365), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n345), .A2(new_n367), .A3(new_n351), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G120gat), .B(G148gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(G176gat), .B(G204gat), .ZN(new_n371));
  XOR2_X1   g170(.A(new_n370), .B(new_n371), .Z(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n366), .A2(new_n368), .A3(new_n372), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n310), .A2(new_n343), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT5), .ZN(new_n379));
  XNOR2_X1  g178(.A(G113gat), .B(G120gat), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT67), .ZN(new_n381));
  AOI21_X1  g180(.A(KEYINPUT1), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n382), .B1(new_n381), .B2(new_n380), .ZN(new_n383));
  XNOR2_X1  g182(.A(G127gat), .B(G134gat), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  XOR2_X1   g185(.A(KEYINPUT68), .B(KEYINPUT1), .Z(new_n387));
  AND2_X1   g186(.A1(new_n387), .A2(new_n384), .ZN(new_n388));
  INV_X1    g187(.A(new_n380), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n386), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(G141gat), .ZN(new_n392));
  INV_X1    g191(.A(G148gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(G141gat), .A2(G148gat), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OR2_X1    g195(.A1(new_n396), .A2(KEYINPUT77), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT2), .ZN(new_n398));
  INV_X1    g197(.A(G155gat), .ZN(new_n399));
  INV_X1    g198(.A(G162gat), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(G155gat), .A2(G162gat), .ZN(new_n402));
  AOI22_X1  g201(.A1(new_n396), .A2(KEYINPUT77), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n397), .A2(new_n403), .ZN(new_n404));
  XOR2_X1   g203(.A(G155gat), .B(G162gat), .Z(new_n405));
  NAND3_X1  g204(.A1(new_n394), .A2(new_n398), .A3(new_n395), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT76), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n405), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n407), .B1(new_n405), .B2(new_n406), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n404), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n391), .A2(new_n411), .ZN(new_n412));
  AOI22_X1  g211(.A1(new_n383), .A2(new_n385), .B1(new_n389), .B2(new_n388), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n405), .A2(new_n406), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(KEYINPUT76), .ZN(new_n415));
  AOI22_X1  g214(.A1(new_n415), .A2(new_n408), .B1(new_n397), .B2(new_n403), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n412), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(G225gat), .A2(G233gat), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n379), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT4), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n417), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT3), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n391), .B1(new_n416), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n416), .A2(new_n424), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n423), .B(new_n419), .C1(new_n425), .C2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n411), .A2(KEYINPUT78), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT78), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n416), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NOR3_X1   g231(.A1(new_n432), .A2(new_n422), .A3(new_n391), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n421), .B1(new_n428), .B2(new_n433), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n429), .A2(new_n431), .A3(new_n422), .A4(new_n413), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n417), .A2(KEYINPUT4), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n413), .B1(new_n411), .B2(KEYINPUT3), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n426), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n437), .A2(new_n379), .A3(new_n419), .A4(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n434), .A2(new_n440), .ZN(new_n441));
  XNOR2_X1  g240(.A(G1gat), .B(G29gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n442), .B(KEYINPUT0), .ZN(new_n443));
  XNOR2_X1  g242(.A(G57gat), .B(G85gat), .ZN(new_n444));
  XOR2_X1   g243(.A(new_n443), .B(new_n444), .Z(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n441), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT6), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n434), .A2(new_n440), .A3(new_n445), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n441), .A2(KEYINPUT6), .A3(new_n446), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  XOR2_X1   g251(.A(G8gat), .B(G36gat), .Z(new_n453));
  XNOR2_X1  g252(.A(new_n453), .B(KEYINPUT75), .ZN(new_n454));
  XNOR2_X1  g253(.A(G64gat), .B(G92gat), .ZN(new_n455));
  XOR2_X1   g254(.A(new_n454), .B(new_n455), .Z(new_n456));
  XNOR2_X1  g255(.A(G211gat), .B(G218gat), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT73), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n457), .B(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(KEYINPUT72), .B(G197gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n460), .B(G204gat), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT22), .ZN(new_n462));
  INV_X1    g261(.A(G211gat), .ZN(new_n463));
  INV_X1    g262(.A(G218gat), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n459), .A2(new_n461), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n459), .B1(new_n465), .B2(new_n461), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g268(.A(KEYINPUT27), .B(G183gat), .ZN(new_n470));
  INV_X1    g269(.A(G190gat), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OR2_X1    g271(.A1(new_n472), .A2(KEYINPUT28), .ZN(new_n473));
  NAND2_X1  g272(.A1(G169gat), .A2(G176gat), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT26), .ZN(new_n475));
  NOR2_X1   g274(.A1(G169gat), .A2(G176gat), .ZN(new_n476));
  NOR4_X1   g275(.A1(KEYINPUT66), .A2(KEYINPUT26), .A3(G169gat), .A4(G176gat), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT66), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n478), .B1(new_n476), .B2(new_n475), .ZN(new_n479));
  OAI221_X1 g278(.A(new_n474), .B1(new_n475), .B2(new_n476), .C1(new_n477), .C2(new_n479), .ZN(new_n480));
  AOI22_X1  g279(.A1(new_n472), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n473), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT65), .ZN(new_n484));
  OR2_X1    g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n486));
  INV_X1    g285(.A(G183gat), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n486), .B1(new_n487), .B2(new_n471), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n483), .A2(new_n484), .ZN(new_n489));
  AND3_X1   g288(.A1(new_n485), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n476), .A2(KEYINPUT23), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT23), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n492), .B1(G169gat), .B2(G176gat), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n491), .A2(new_n474), .A3(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT25), .B1(new_n490), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT64), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n488), .A2(new_n483), .ZN(new_n498));
  NOR2_X1   g297(.A1(KEYINPUT64), .A2(KEYINPUT25), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n497), .B(new_n498), .C1(new_n494), .C2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n482), .A2(new_n495), .A3(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT74), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n482), .A2(KEYINPUT74), .A3(new_n495), .A4(new_n500), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(G226gat), .ZN(new_n506));
  INV_X1    g305(.A(G233gat), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n508), .A2(KEYINPUT29), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n508), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n501), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n469), .B1(new_n510), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n503), .A2(new_n508), .A3(new_n504), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n501), .A2(new_n509), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(new_n469), .A3(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n456), .B1(new_n514), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n456), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n512), .B1(new_n505), .B2(new_n509), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n517), .B(new_n520), .C1(new_n521), .C2(new_n469), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n519), .A2(KEYINPUT30), .A3(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n514), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT30), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n524), .A2(new_n525), .A3(new_n520), .A4(new_n517), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n452), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(G228gat), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n529), .A2(new_n507), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(KEYINPUT29), .B1(new_n416), .B2(new_n424), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n461), .A2(new_n465), .ZN(new_n533));
  INV_X1    g332(.A(new_n459), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(new_n466), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n531), .B1(new_n532), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n535), .A2(KEYINPUT80), .A3(new_n466), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT80), .ZN(new_n539));
  AOI21_X1  g338(.A(KEYINPUT29), .B1(new_n468), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(new_n424), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n537), .B1(new_n542), .B2(new_n432), .ZN(new_n543));
  AOI21_X1  g342(.A(KEYINPUT29), .B1(new_n535), .B2(new_n466), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n411), .B1(new_n544), .B2(KEYINPUT3), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n469), .B1(new_n427), .B2(KEYINPUT29), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n531), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(KEYINPUT79), .B(KEYINPUT31), .ZN(new_n548));
  NOR3_X1   g347(.A1(new_n543), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n548), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT29), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n551), .B1(new_n467), .B2(new_n468), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n416), .B1(new_n552), .B2(new_n424), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n532), .A2(new_n536), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n530), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(KEYINPUT3), .B1(new_n538), .B2(new_n540), .ZN(new_n556));
  INV_X1    g355(.A(new_n432), .ZN(new_n557));
  OAI211_X1 g356(.A(new_n531), .B(new_n546), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n550), .B1(new_n555), .B2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G78gat), .B(G106gat), .ZN(new_n560));
  INV_X1    g359(.A(G50gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n560), .B(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(G22gat), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NOR3_X1   g363(.A1(new_n549), .A2(new_n559), .A3(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n548), .B1(new_n543), .B2(new_n547), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n555), .A2(new_n558), .A3(new_n550), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n563), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n528), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(G227gat), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n572), .A2(new_n507), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n501), .A2(new_n413), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n391), .A2(new_n482), .A3(new_n495), .A4(new_n500), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT34), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI211_X1 g377(.A(KEYINPUT34), .B(new_n573), .C1(new_n574), .C2(new_n575), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n574), .A2(new_n575), .A3(new_n573), .ZN(new_n581));
  XOR2_X1   g380(.A(KEYINPUT69), .B(KEYINPUT33), .Z(new_n582));
  INV_X1    g381(.A(KEYINPUT32), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  XOR2_X1   g384(.A(G71gat), .B(G99gat), .Z(new_n586));
  XNOR2_X1  g385(.A(G15gat), .B(G43gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT70), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n583), .B1(new_n588), .B2(new_n582), .ZN(new_n591));
  AND3_X1   g390(.A1(new_n581), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n590), .B1(new_n581), .B2(new_n591), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n589), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT71), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n580), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  OAI211_X1 g395(.A(new_n589), .B(KEYINPUT71), .C1(new_n592), .C2(new_n593), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n580), .B(new_n589), .C1(new_n593), .C2(new_n592), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n598), .A2(KEYINPUT36), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n594), .B1(new_n578), .B2(new_n579), .ZN(new_n601));
  AOI21_X1  g400(.A(KEYINPUT36), .B1(new_n601), .B2(new_n599), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT38), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT37), .ZN(new_n606));
  OAI211_X1 g405(.A(new_n517), .B(new_n606), .C1(new_n521), .C2(new_n469), .ZN(new_n607));
  AND2_X1   g406(.A1(new_n607), .A2(new_n456), .ZN(new_n608));
  OAI21_X1  g407(.A(KEYINPUT37), .B1(new_n514), .B2(new_n518), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n605), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n515), .A2(new_n536), .A3(new_n516), .ZN(new_n611));
  OAI211_X1 g410(.A(new_n611), .B(KEYINPUT37), .C1(new_n521), .C2(new_n536), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n607), .A2(new_n612), .A3(new_n605), .A4(new_n456), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(new_n522), .ZN(new_n614));
  NOR3_X1   g413(.A1(new_n452), .A2(new_n610), .A3(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n412), .A2(new_n419), .A3(new_n417), .ZN(new_n616));
  AOI22_X1  g415(.A1(new_n435), .A2(new_n436), .B1(new_n426), .B2(new_n438), .ZN(new_n617));
  OAI211_X1 g416(.A(KEYINPUT39), .B(new_n616), .C1(new_n617), .C2(new_n419), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n437), .A2(new_n439), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT39), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n619), .A2(new_n620), .A3(new_n420), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n618), .A2(new_n621), .A3(new_n445), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT40), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n618), .A2(new_n621), .A3(KEYINPUT40), .A4(new_n445), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n624), .A2(new_n447), .A3(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n569), .B1(new_n626), .B2(new_n527), .ZN(new_n627));
  OAI211_X1 g426(.A(new_n571), .B(new_n604), .C1(new_n615), .C2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n566), .A2(new_n563), .A3(new_n567), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n564), .B1(new_n549), .B2(new_n559), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n598), .A2(new_n629), .A3(new_n630), .A4(new_n599), .ZN(new_n631));
  OAI21_X1  g430(.A(KEYINPUT35), .B1(new_n631), .B2(new_n528), .ZN(new_n632));
  AOI22_X1  g431(.A1(new_n450), .A2(new_n451), .B1(new_n523), .B2(new_n526), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT35), .ZN(new_n634));
  AND2_X1   g433(.A1(new_n601), .A2(new_n599), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n633), .A2(new_n634), .A3(new_n569), .A4(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  AOI211_X1 g436(.A(new_n261), .B(new_n378), .C1(new_n628), .C2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n452), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(G1gat), .ZN(G1324gat));
  INV_X1    g440(.A(KEYINPUT42), .ZN(new_n642));
  INV_X1    g441(.A(new_n527), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n638), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(G8gat), .ZN(new_n645));
  XOR2_X1   g444(.A(KEYINPUT16), .B(G8gat), .Z(new_n646));
  NAND3_X1  g445(.A1(new_n638), .A2(new_n643), .A3(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n642), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n648), .B1(new_n642), .B2(new_n647), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n649), .B(KEYINPUT95), .Z(G1325gat));
  INV_X1    g449(.A(new_n604), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n638), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n601), .A2(new_n599), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n653), .A2(G15gat), .ZN(new_n654));
  AOI22_X1  g453(.A1(new_n652), .A2(G15gat), .B1(new_n638), .B2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT96), .ZN(G1326gat));
  NAND2_X1  g455(.A1(new_n638), .A2(new_n570), .ZN(new_n657));
  XNOR2_X1  g456(.A(KEYINPUT43), .B(G22gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(G1327gat));
  AOI21_X1  g458(.A(new_n310), .B1(new_n628), .B2(new_n637), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n343), .A2(new_n261), .A3(new_n376), .ZN(new_n661));
  AND2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n662), .A2(new_n211), .A3(new_n639), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(KEYINPUT97), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT45), .ZN(new_n665));
  AND3_X1   g464(.A1(new_n632), .A2(KEYINPUT99), .A3(new_n636), .ZN(new_n666));
  AOI21_X1  g465(.A(KEYINPUT99), .B1(new_n632), .B2(new_n636), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n628), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT44), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n302), .A2(new_n309), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n668), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n628), .A2(new_n637), .ZN(new_n672));
  OAI211_X1 g471(.A(KEYINPUT98), .B(KEYINPUT44), .C1(new_n672), .C2(new_n310), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT98), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n674), .B1(new_n660), .B2(new_n669), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n671), .A2(new_n673), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(new_n661), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n678), .A2(KEYINPUT100), .A3(new_n639), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT100), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n680), .B1(new_n677), .B2(new_n452), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n679), .A2(G29gat), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n665), .A2(new_n682), .ZN(G1328gat));
  INV_X1    g482(.A(new_n210), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n684), .B1(new_n677), .B2(new_n527), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n684), .B1(KEYINPUT101), .B2(KEYINPUT46), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n662), .A2(new_n643), .A3(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(KEYINPUT101), .A2(KEYINPUT46), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n685), .A2(new_n689), .ZN(G1329gat));
  NAND3_X1  g489(.A1(new_n678), .A2(G43gat), .A3(new_n651), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n662), .A2(new_n635), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n691), .B1(G43gat), .B2(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g493(.A(G50gat), .B1(new_n677), .B2(new_n569), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n662), .A2(new_n561), .A3(new_n570), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT103), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n696), .A2(new_n697), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n695), .A2(KEYINPUT48), .A3(new_n698), .A4(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(KEYINPUT48), .B1(new_n695), .B2(new_n696), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT102), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AOI211_X1 g502(.A(KEYINPUT102), .B(KEYINPUT48), .C1(new_n695), .C2(new_n696), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n700), .B1(new_n703), .B2(new_n704), .ZN(G1331gat));
  NOR4_X1   g504(.A1(new_n670), .A2(new_n342), .A3(new_n260), .A4(new_n377), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n668), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n707), .A2(new_n452), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(new_n317), .ZN(G1332gat));
  XNOR2_X1  g508(.A(new_n707), .B(KEYINPUT104), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n643), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n711), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n712));
  XOR2_X1   g511(.A(KEYINPUT49), .B(G64gat), .Z(new_n713));
  OAI21_X1  g512(.A(new_n712), .B1(new_n711), .B2(new_n713), .ZN(G1333gat));
  NAND3_X1  g513(.A1(new_n710), .A2(G71gat), .A3(new_n651), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n707), .A2(new_n653), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n715), .B1(G71gat), .B2(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(KEYINPUT105), .B(KEYINPUT50), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1334gat));
  NAND2_X1  g518(.A1(new_n710), .A2(new_n570), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g520(.A1(new_n261), .A2(new_n342), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n722), .A2(new_n377), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n676), .A2(new_n639), .A3(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT106), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n271), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n726), .B1(new_n725), .B2(new_n724), .ZN(new_n727));
  INV_X1    g526(.A(new_n722), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n668), .A2(KEYINPUT51), .A3(new_n670), .A4(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(KEYINPUT107), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT99), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n596), .A2(new_n597), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n630), .A2(new_n629), .A3(new_n599), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n634), .B1(new_n734), .B2(new_n633), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n569), .A2(new_n635), .A3(new_n634), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n736), .A2(new_n528), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n731), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n632), .A2(KEYINPUT99), .A3(new_n636), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n310), .B1(new_n740), .B2(new_n628), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT107), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n741), .A2(new_n742), .A3(KEYINPUT51), .A4(new_n728), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n730), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n615), .A2(new_n627), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n599), .A2(KEYINPUT36), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n746), .B1(new_n597), .B2(new_n596), .ZN(new_n747));
  OAI22_X1  g546(.A1(new_n747), .A2(new_n602), .B1(new_n633), .B2(new_n569), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n749), .B1(new_n738), .B2(new_n739), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n750), .A2(new_n310), .A3(new_n722), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n744), .B1(KEYINPUT51), .B2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n639), .A2(new_n271), .A3(new_n376), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n727), .B1(new_n753), .B2(new_n754), .ZN(G1336gat));
  INV_X1    g554(.A(KEYINPUT109), .ZN(new_n756));
  XNOR2_X1  g555(.A(KEYINPUT108), .B(KEYINPUT51), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n756), .B1(new_n751), .B2(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n668), .A2(new_n670), .A3(new_n728), .ZN(new_n759));
  INV_X1    g558(.A(new_n757), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n759), .A2(KEYINPUT109), .A3(new_n760), .ZN(new_n761));
  AOI22_X1  g560(.A1(new_n758), .A2(new_n761), .B1(new_n730), .B2(new_n743), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n527), .A2(G92gat), .A3(new_n377), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(KEYINPUT110), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(KEYINPUT109), .B1(new_n759), .B2(new_n760), .ZN(new_n766));
  AND3_X1   g565(.A1(new_n759), .A2(KEYINPUT109), .A3(new_n760), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n744), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT110), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n768), .A2(new_n769), .A3(new_n763), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n676), .A2(new_n723), .ZN(new_n771));
  OAI21_X1  g570(.A(G92gat), .B1(new_n771), .B2(new_n527), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n765), .A2(new_n770), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(KEYINPUT52), .ZN(new_n774));
  XNOR2_X1  g573(.A(KEYINPUT111), .B(KEYINPUT52), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n772), .B(new_n775), .C1(new_n753), .C2(new_n764), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n774), .A2(new_n776), .ZN(G1337gat));
  OAI21_X1  g576(.A(G99gat), .B1(new_n771), .B2(new_n604), .ZN(new_n778));
  OR3_X1    g577(.A1(new_n653), .A2(new_n377), .A3(G99gat), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n778), .B1(new_n753), .B2(new_n779), .ZN(G1338gat));
  NAND3_X1  g579(.A1(new_n676), .A2(new_n570), .A3(new_n723), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT114), .ZN(new_n782));
  OR2_X1    g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n782), .ZN(new_n784));
  XNOR2_X1  g583(.A(KEYINPUT112), .B(G106gat), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n569), .A2(G106gat), .A3(new_n377), .ZN(new_n787));
  AOI21_X1  g586(.A(KEYINPUT53), .B1(new_n752), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n781), .A2(new_n785), .ZN(new_n790));
  INV_X1    g589(.A(new_n787), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n790), .B1(new_n762), .B2(new_n791), .ZN(new_n792));
  AND3_X1   g591(.A1(new_n792), .A2(KEYINPUT113), .A3(KEYINPUT53), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT113), .B1(new_n792), .B2(KEYINPUT53), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n789), .B1(new_n793), .B2(new_n794), .ZN(G1339gat));
  INV_X1    g594(.A(KEYINPUT55), .ZN(new_n796));
  OAI21_X1  g595(.A(KEYINPUT94), .B1(new_n361), .B2(new_n362), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n327), .A2(new_n354), .A3(new_n283), .A4(KEYINPUT10), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n352), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n799), .A2(new_n367), .ZN(new_n800));
  XNOR2_X1  g599(.A(KEYINPUT116), .B(KEYINPUT54), .ZN(new_n801));
  AOI211_X1 g600(.A(new_n796), .B(new_n372), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n803), .B1(new_n364), .B2(new_n365), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n799), .A2(new_n367), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT115), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(KEYINPUT54), .B1(new_n799), .B2(new_n367), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n345), .A2(new_n351), .ZN(new_n808));
  AOI221_X4 g607(.A(new_n365), .B1(new_n808), .B2(new_n355), .C1(new_n797), .C2(new_n798), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT115), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n807), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n802), .B1(new_n806), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n375), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n810), .B1(new_n807), .B2(new_n809), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n366), .A2(KEYINPUT115), .A3(KEYINPUT54), .A4(new_n805), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n373), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(KEYINPUT55), .B1(new_n816), .B2(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(KEYINPUT117), .B1(new_n813), .B2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n375), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n822), .B1(new_n816), .B2(new_n802), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT117), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n818), .B1(new_n814), .B2(new_n815), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n823), .B(new_n824), .C1(KEYINPUT55), .C2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n821), .A2(new_n260), .A3(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(KEYINPUT118), .B1(new_n238), .B2(new_n239), .ZN(new_n828));
  INV_X1    g627(.A(new_n247), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n244), .A2(new_n245), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n238), .A2(KEYINPUT118), .A3(new_n239), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n254), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n833), .A2(new_n259), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n376), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n670), .B1(new_n827), .B2(new_n835), .ZN(new_n836));
  AND4_X1   g635(.A1(new_n670), .A2(new_n834), .A3(new_n821), .A4(new_n826), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n342), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OR2_X1    g637(.A1(new_n378), .A2(new_n260), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n452), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n840), .A2(new_n527), .A3(new_n734), .ZN(new_n841));
  AOI21_X1  g640(.A(G113gat), .B1(new_n841), .B2(new_n260), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n838), .A2(new_n839), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(new_n569), .ZN(new_n844));
  NOR4_X1   g643(.A1(new_n844), .A2(new_n452), .A3(new_n643), .A4(new_n653), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n260), .A2(G113gat), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n842), .B1(new_n845), .B2(new_n846), .ZN(G1340gat));
  AOI21_X1  g646(.A(G120gat), .B1(new_n841), .B2(new_n376), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n376), .A2(G120gat), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n848), .B1(new_n845), .B2(new_n849), .ZN(G1341gat));
  INV_X1    g649(.A(G127gat), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n841), .A2(new_n851), .A3(new_n343), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n845), .A2(new_n343), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n852), .B1(new_n853), .B2(new_n851), .ZN(G1342gat));
  INV_X1    g653(.A(G134gat), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n841), .A2(new_n855), .A3(new_n670), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n856), .A2(KEYINPUT56), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(KEYINPUT56), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n845), .A2(new_n670), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n857), .B(new_n858), .C1(new_n855), .C2(new_n859), .ZN(G1343gat));
  NAND3_X1  g659(.A1(new_n604), .A2(new_n639), .A3(new_n527), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n823), .B1(KEYINPUT55), .B2(new_n825), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n835), .B1(new_n862), .B2(new_n261), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n310), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n670), .A2(new_n834), .A3(new_n821), .A4(new_n826), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n343), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n378), .A2(new_n260), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n570), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n861), .B1(new_n868), .B2(KEYINPUT57), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n569), .B1(new_n838), .B2(new_n839), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT57), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(G141gat), .B1(new_n873), .B2(new_n261), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n651), .A2(new_n569), .ZN(new_n875));
  AND3_X1   g674(.A1(new_n840), .A2(new_n527), .A3(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n876), .A2(new_n392), .A3(new_n260), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g677(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n878), .B(new_n879), .ZN(G1344gat));
  NAND3_X1  g679(.A1(new_n876), .A2(new_n393), .A3(new_n376), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n873), .A2(new_n377), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n882), .A2(KEYINPUT59), .A3(new_n393), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT59), .ZN(new_n884));
  OR3_X1    g683(.A1(new_n310), .A2(KEYINPUT120), .A3(new_n862), .ZN(new_n885));
  OAI21_X1  g684(.A(KEYINPUT120), .B1(new_n310), .B2(new_n862), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n885), .A2(new_n834), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n343), .B1(new_n887), .B2(new_n864), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n871), .B(new_n570), .C1(new_n888), .C2(new_n867), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n870), .A2(new_n871), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n861), .A2(new_n377), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n884), .B1(new_n892), .B2(G148gat), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n881), .B1(new_n883), .B2(new_n893), .ZN(G1345gat));
  OAI21_X1  g693(.A(G155gat), .B1(new_n873), .B2(new_n342), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n876), .A2(new_n399), .A3(new_n343), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(G1346gat));
  OAI21_X1  g696(.A(G162gat), .B1(new_n873), .B2(new_n310), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n876), .A2(new_n400), .A3(new_n670), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(G1347gat));
  AOI21_X1  g699(.A(new_n639), .B1(new_n838), .B2(new_n839), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n631), .A2(new_n527), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT121), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  OR3_X1    g703(.A1(new_n904), .A2(G169gat), .A3(new_n261), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n643), .A2(new_n452), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n906), .A2(new_n653), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n827), .A2(new_n835), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n310), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n343), .B1(new_n909), .B2(new_n865), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n569), .B(new_n907), .C1(new_n910), .C2(new_n867), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT122), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n843), .A2(KEYINPUT122), .A3(new_n569), .A4(new_n907), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(new_n260), .ZN(new_n916));
  AND3_X1   g715(.A1(new_n916), .A2(KEYINPUT123), .A3(G169gat), .ZN(new_n917));
  AOI21_X1  g716(.A(KEYINPUT123), .B1(new_n916), .B2(G169gat), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n905), .B1(new_n917), .B2(new_n918), .ZN(G1348gat));
  INV_X1    g718(.A(G176gat), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n920), .B1(new_n915), .B2(new_n376), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n904), .A2(G176gat), .A3(new_n377), .ZN(new_n922));
  OR3_X1    g721(.A1(new_n921), .A2(KEYINPUT124), .A3(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(KEYINPUT124), .B1(new_n921), .B2(new_n922), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(G1349gat));
  AND4_X1   g724(.A1(new_n470), .A2(new_n901), .A3(new_n343), .A4(new_n903), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n913), .A2(new_n343), .A3(new_n914), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n926), .B1(new_n927), .B2(G183gat), .ZN(new_n928));
  AOI211_X1 g727(.A(KEYINPUT125), .B(KEYINPUT60), .C1(new_n928), .C2(KEYINPUT126), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(KEYINPUT126), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT125), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT60), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n933), .B1(new_n928), .B2(KEYINPUT125), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n929), .B1(new_n932), .B2(new_n934), .ZN(G1350gat));
  INV_X1    g734(.A(KEYINPUT61), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n915), .A2(new_n670), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n936), .B1(new_n937), .B2(G190gat), .ZN(new_n938));
  AOI211_X1 g737(.A(KEYINPUT61), .B(new_n471), .C1(new_n915), .C2(new_n670), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n670), .A2(new_n471), .ZN(new_n940));
  OAI22_X1  g739(.A1(new_n938), .A2(new_n939), .B1(new_n904), .B2(new_n940), .ZN(G1351gat));
  NOR2_X1   g740(.A1(new_n651), .A2(new_n906), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n889), .A2(new_n890), .A3(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(G197gat), .ZN(new_n944));
  NOR3_X1   g743(.A1(new_n943), .A2(new_n944), .A3(new_n261), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n901), .A2(new_n643), .A3(new_n875), .ZN(new_n946));
  XOR2_X1   g745(.A(new_n946), .B(KEYINPUT127), .Z(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(new_n260), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n945), .B1(new_n948), .B2(new_n944), .ZN(G1352gat));
  NOR3_X1   g748(.A1(new_n946), .A2(G204gat), .A3(new_n377), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT62), .ZN(new_n951));
  OAI21_X1  g750(.A(G204gat), .B1(new_n943), .B2(new_n377), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(G1353gat));
  NAND3_X1  g752(.A1(new_n947), .A2(new_n463), .A3(new_n343), .ZN(new_n954));
  OR2_X1    g753(.A1(new_n943), .A2(new_n342), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n955), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n956));
  INV_X1    g755(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g756(.A(KEYINPUT63), .B1(new_n955), .B2(G211gat), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n954), .B1(new_n957), .B2(new_n958), .ZN(G1354gat));
  NAND3_X1  g758(.A1(new_n947), .A2(new_n464), .A3(new_n670), .ZN(new_n960));
  OAI21_X1  g759(.A(G218gat), .B1(new_n943), .B2(new_n310), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(G1355gat));
endmodule


