//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 1 1 0 0 1 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 0 1 1 0 1 1 0 1 0 1 1 0 0 0 1 1 1 0 1 0 0 1 0 0 1 1 0 0 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:12 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1369, new_n1370, new_n1371,
    new_n1372, new_n1373, new_n1374, new_n1375, new_n1376, new_n1377,
    new_n1378, new_n1379, new_n1380, new_n1381, new_n1382, new_n1383,
    new_n1384;
  OR2_X1    g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  NOR3_X1   g0001(.A1(new_n201), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0002(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0003(.A(G1), .ZN(new_n204));
  INV_X1    g0004(.A(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(KEYINPUT64), .ZN(new_n212));
  INV_X1    g0012(.A(KEYINPUT64), .ZN(new_n213));
  NAND3_X1  g0013(.A1(new_n213), .A2(G1), .A3(G13), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n205), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n201), .A2(G50), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g0020(.A(KEYINPUT65), .B(G77), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G58), .A2(G232), .ZN(new_n227));
  NAND4_X1  g0027(.A1(new_n224), .A2(new_n225), .A3(new_n226), .A4(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n207), .B1(new_n223), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n210), .B(new_n220), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XOR2_X1   g0031(.A(G250), .B(G257), .Z(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT66), .B(KEYINPUT67), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  INV_X1    g0037(.A(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n236), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  OAI21_X1  g0049(.A(G20), .B1(new_n201), .B2(G50), .ZN(new_n250));
  INV_X1    g0050(.A(G150), .ZN(new_n251));
  NOR2_X1   g0051(.A1(G20), .A2(G33), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n250), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  NOR2_X1   g0054(.A1(KEYINPUT8), .A2(G58), .ZN(new_n255));
  XOR2_X1   g0055(.A(KEYINPUT69), .B(G58), .Z(new_n256));
  AOI21_X1  g0056(.A(new_n255), .B1(new_n256), .B2(KEYINPUT8), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(G20), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT70), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n259), .B(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n254), .B1(new_n257), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n216), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n204), .A2(G13), .A3(G20), .ZN(new_n267));
  NAND4_X1  g0067(.A1(new_n212), .A2(new_n214), .A3(new_n267), .A4(new_n263), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n204), .A2(G20), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G50), .ZN(new_n270));
  OAI22_X1  g0070(.A1(new_n268), .A2(new_n270), .B1(G50), .B2(new_n267), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n266), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(KEYINPUT9), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT72), .ZN(new_n274));
  XNOR2_X1  g0074(.A(new_n273), .B(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n272), .A2(KEYINPUT9), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT73), .ZN(new_n277));
  XNOR2_X1  g0077(.A(new_n276), .B(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G190), .ZN(new_n279));
  INV_X1    g0079(.A(G200), .ZN(new_n280));
  INV_X1    g0080(.A(G274), .ZN(new_n281));
  INV_X1    g0081(.A(new_n211), .ZN(new_n282));
  NAND2_X1  g0082(.A1(G33), .A2(G41), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G41), .ZN(new_n285));
  INV_X1    g0085(.A(G45), .ZN(new_n286));
  AOI21_X1  g0086(.A(G1), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n287), .B1(new_n282), .B2(new_n283), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n289), .B1(G226), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n215), .A2(new_n283), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n221), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT3), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G33), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n293), .B1(new_n294), .B2(new_n299), .ZN(new_n300));
  NOR2_X1   g0100(.A1(G222), .A2(G1698), .ZN(new_n301));
  XOR2_X1   g0101(.A(KEYINPUT68), .B(G223), .Z(new_n302));
  AOI21_X1  g0102(.A(new_n301), .B1(new_n302), .B2(G1698), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n303), .A2(new_n298), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n291), .B1(new_n300), .B2(new_n304), .ZN(new_n305));
  MUX2_X1   g0105(.A(new_n279), .B(new_n280), .S(new_n305), .Z(new_n306));
  NAND3_X1  g0106(.A1(new_n275), .A2(new_n278), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(KEYINPUT10), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT10), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n275), .A2(new_n278), .A3(new_n309), .A4(new_n306), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  OR2_X1    g0111(.A1(new_n305), .A2(G179), .ZN(new_n312));
  INV_X1    g0112(.A(new_n272), .ZN(new_n313));
  INV_X1    g0113(.A(G169), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n305), .A2(new_n314), .ZN(new_n315));
  AND3_X1   g0115(.A1(new_n312), .A2(new_n313), .A3(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n311), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n261), .A2(G77), .ZN(new_n319));
  INV_X1    g0119(.A(G68), .ZN(new_n320));
  AOI22_X1  g0120(.A1(new_n252), .A2(G50), .B1(G20), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n265), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  OR2_X1    g0122(.A1(new_n322), .A2(KEYINPUT11), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(KEYINPUT11), .ZN(new_n324));
  INV_X1    g0124(.A(new_n269), .ZN(new_n325));
  NOR3_X1   g0125(.A1(new_n268), .A2(new_n320), .A3(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(KEYINPUT12), .B1(new_n267), .B2(G68), .ZN(new_n327));
  OR3_X1    g0127(.A1(new_n267), .A2(KEYINPUT12), .A3(G68), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n323), .A2(new_n324), .A3(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT13), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n289), .B1(G238), .B2(new_n290), .ZN(new_n333));
  NAND2_X1  g0133(.A1(G33), .A2(G97), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n238), .A2(G1698), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n335), .B1(G226), .B2(G1698), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n334), .B1(new_n336), .B2(new_n298), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n293), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n332), .B1(new_n333), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n333), .A2(new_n332), .A3(new_n338), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G200), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n340), .A2(G190), .A3(new_n341), .ZN(new_n344));
  AND3_X1   g0144(.A1(new_n331), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n341), .ZN(new_n347));
  OAI21_X1  g0147(.A(G169), .B1(new_n347), .B2(new_n339), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT14), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT14), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n342), .A2(new_n350), .A3(G169), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n340), .A2(G179), .A3(new_n341), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n349), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n330), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n346), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n299), .A2(G238), .A3(G1698), .ZN(new_n356));
  INV_X1    g0156(.A(G1698), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n299), .A2(G232), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(G107), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n356), .B(new_n358), .C1(new_n359), .C2(new_n299), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n293), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n289), .B1(G244), .B2(new_n290), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n314), .ZN(new_n364));
  INV_X1    g0164(.A(G77), .ZN(new_n365));
  NOR3_X1   g0165(.A1(new_n268), .A2(new_n365), .A3(new_n325), .ZN(new_n366));
  XOR2_X1   g0166(.A(new_n366), .B(KEYINPUT71), .Z(new_n367));
  XNOR2_X1  g0167(.A(KEYINPUT15), .B(G87), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n294), .A2(G20), .B1(new_n369), .B2(new_n259), .ZN(new_n370));
  XOR2_X1   g0170(.A(KEYINPUT8), .B(G58), .Z(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n370), .B1(new_n253), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n267), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n373), .A2(new_n264), .B1(new_n221), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n367), .A2(new_n375), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n364), .B(new_n376), .C1(G179), .C2(new_n363), .ZN(new_n377));
  INV_X1    g0177(.A(new_n363), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n378), .A2(new_n280), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n367), .B(new_n375), .C1(new_n363), .C2(new_n279), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n377), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  OR3_X1    g0181(.A1(new_n318), .A2(new_n355), .A3(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n257), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n383), .A2(new_n325), .ZN(new_n384));
  INV_X1    g0184(.A(new_n268), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n384), .A2(new_n385), .B1(new_n374), .B2(new_n383), .ZN(new_n386));
  XNOR2_X1  g0186(.A(KEYINPUT69), .B(G58), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n201), .B1(new_n387), .B2(new_n320), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n388), .A2(G20), .B1(G159), .B2(new_n252), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n258), .A2(KEYINPUT74), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT74), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(G33), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n390), .A2(new_n392), .A3(KEYINPUT3), .ZN(new_n393));
  AOI21_X1  g0193(.A(G20), .B1(new_n393), .B2(new_n297), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT7), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(G68), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n394), .A2(new_n395), .ZN(new_n398));
  OAI211_X1 g0198(.A(KEYINPUT16), .B(new_n389), .C1(new_n397), .C2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n264), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n395), .B1(new_n299), .B2(G20), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n390), .A2(new_n392), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT75), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n402), .A2(new_n403), .A3(new_n296), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n395), .A2(G20), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n295), .A2(KEYINPUT75), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n407), .B1(new_n402), .B2(new_n296), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n401), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(G68), .ZN(new_n410));
  AOI21_X1  g0210(.A(KEYINPUT16), .B1(new_n410), .B2(new_n389), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n386), .B1(new_n400), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT76), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT16), .ZN(new_n414));
  XNOR2_X1  g0214(.A(KEYINPUT74), .B(G33), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n415), .A2(KEYINPUT3), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n404), .B(new_n405), .C1(new_n416), .C2(new_n407), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n320), .B1(new_n417), .B2(new_n401), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n388), .A2(G20), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n252), .A2(G159), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n414), .B1(new_n418), .B2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n422), .A2(new_n264), .A3(new_n399), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT76), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n423), .A2(new_n424), .A3(new_n386), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n290), .A2(G232), .B1(new_n284), .B2(new_n287), .ZN(new_n426));
  INV_X1    g0226(.A(new_n297), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n427), .B1(new_n415), .B2(KEYINPUT3), .ZN(new_n428));
  MUX2_X1   g0228(.A(G223), .B(G226), .S(G1698), .Z(new_n429));
  AOI22_X1  g0229(.A1(new_n428), .A2(new_n429), .B1(G33), .B2(G87), .ZN(new_n430));
  OAI211_X1 g0230(.A(G179), .B(new_n426), .C1(new_n430), .C2(new_n292), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n429), .A2(new_n393), .A3(new_n297), .ZN(new_n432));
  NAND2_X1  g0232(.A1(G33), .A2(G87), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n292), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n287), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n282), .A2(new_n283), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n288), .B1(new_n437), .B2(new_n238), .ZN(new_n438));
  OAI21_X1  g0238(.A(G169), .B1(new_n434), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n431), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n413), .A2(new_n425), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT18), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT18), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n413), .A2(new_n443), .A3(new_n425), .A4(new_n440), .ZN(new_n444));
  OAI211_X1 g0244(.A(G190), .B(new_n426), .C1(new_n430), .C2(new_n292), .ZN(new_n445));
  OAI21_X1  g0245(.A(G200), .B1(new_n434), .B2(new_n438), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n386), .B(new_n447), .C1(new_n400), .C2(new_n411), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT17), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n423), .A2(KEYINPUT17), .A3(new_n386), .A4(new_n447), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n442), .A2(new_n444), .A3(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT5), .ZN(new_n455));
  OAI21_X1  g0255(.A(KEYINPUT79), .B1(new_n455), .B2(G41), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT79), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n457), .A2(new_n285), .A3(KEYINPUT5), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n286), .A2(G1), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n455), .A2(G41), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n456), .A2(new_n458), .A3(new_n459), .A4(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n461), .A2(G270), .A3(new_n436), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT83), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n461), .A2(KEYINPUT83), .A3(G270), .A4(new_n436), .ZN(new_n465));
  AND2_X1   g0265(.A1(new_n459), .A2(new_n460), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n466), .A2(new_n284), .A3(new_n458), .A4(new_n456), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(KEYINPUT84), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n462), .A2(new_n463), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT84), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n470), .A2(new_n471), .A3(new_n467), .A4(new_n465), .ZN(new_n472));
  MUX2_X1   g0272(.A(G257), .B(G264), .S(G1698), .Z(new_n473));
  NAND3_X1  g0273(.A1(new_n473), .A2(new_n393), .A3(new_n297), .ZN(new_n474));
  INV_X1    g0274(.A(G303), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n474), .B1(new_n475), .B2(new_n299), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT85), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n475), .B1(new_n295), .B2(new_n297), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n479), .B1(new_n428), .B2(new_n473), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n292), .B1(new_n480), .B2(KEYINPUT85), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n469), .A2(new_n472), .B1(new_n478), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G190), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n258), .A2(G1), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n268), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(G116), .ZN(new_n486));
  INV_X1    g0286(.A(G116), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n374), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(G20), .B1(G33), .B2(G283), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n258), .A2(G97), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n489), .A2(new_n490), .B1(G20), .B2(new_n487), .ZN(new_n491));
  AND3_X1   g0291(.A1(new_n264), .A2(KEYINPUT20), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(KEYINPUT20), .B1(new_n264), .B2(new_n491), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n486), .B(new_n488), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n483), .B(new_n495), .C1(new_n280), .C2(new_n482), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT21), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n494), .A2(G169), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n497), .B1(new_n482), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n469), .A2(new_n472), .ZN(new_n500));
  INV_X1    g0300(.A(G179), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n501), .B1(new_n481), .B2(new_n478), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n500), .A2(new_n494), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n481), .A2(new_n478), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n505), .A2(KEYINPUT21), .A3(G169), .A4(new_n494), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n496), .A2(new_n499), .A3(new_n503), .A4(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n284), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n508), .A2(new_n461), .ZN(new_n509));
  AND2_X1   g0309(.A1(new_n461), .A2(new_n436), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n509), .B1(new_n510), .B2(G257), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n222), .A2(G1698), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n393), .A2(new_n297), .A3(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT4), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n295), .A2(new_n297), .A3(G250), .A4(G1698), .ZN(new_n516));
  AND2_X1   g0316(.A1(KEYINPUT4), .A2(G244), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n295), .A2(new_n297), .A3(new_n517), .A4(new_n357), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G33), .A2(G283), .ZN(new_n519));
  AND3_X1   g0319(.A1(new_n516), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n515), .A2(new_n520), .A3(KEYINPUT78), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n293), .ZN(new_n522));
  AOI21_X1  g0322(.A(KEYINPUT78), .B1(new_n515), .B2(new_n520), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n511), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g0324(.A(KEYINPUT80), .B1(new_n524), .B2(G179), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT78), .ZN(new_n526));
  AOI21_X1  g0326(.A(KEYINPUT4), .B1(new_n428), .B2(new_n512), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n516), .A2(new_n518), .A3(new_n519), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n529), .A2(new_n293), .A3(new_n521), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT80), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n530), .A2(new_n531), .A3(new_n501), .A4(new_n511), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n525), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n359), .B1(new_n417), .B2(new_n401), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT6), .ZN(new_n535));
  INV_X1    g0335(.A(G97), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n536), .A2(new_n359), .ZN(new_n537));
  NOR2_X1   g0337(.A1(G97), .A2(G107), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n535), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n359), .A2(KEYINPUT77), .A3(KEYINPUT6), .A4(G97), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT77), .ZN(new_n541));
  NAND2_X1  g0341(.A1(KEYINPUT6), .A2(G97), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n541), .B1(new_n542), .B2(G107), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n539), .A2(new_n540), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(G20), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n545), .B1(new_n365), .B2(new_n253), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n264), .B1(new_n534), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n267), .A2(G97), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n548), .B1(new_n485), .B2(G97), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n524), .A2(new_n314), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n533), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n461), .A2(G264), .A3(new_n436), .ZN(new_n552));
  INV_X1    g0352(.A(G294), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n415), .A2(new_n553), .ZN(new_n554));
  MUX2_X1   g0354(.A(G250), .B(G257), .S(G1698), .Z(new_n555));
  AOI21_X1  g0355(.A(new_n554), .B1(new_n428), .B2(new_n555), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n467), .B(new_n552), .C1(new_n556), .C2(new_n292), .ZN(new_n557));
  NOR3_X1   g0357(.A1(new_n557), .A2(KEYINPUT87), .A3(G190), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT22), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n205), .A2(G87), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n559), .B1(new_n298), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n402), .A2(new_n205), .A3(G116), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT86), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n563), .B1(new_n205), .B2(G107), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT23), .ZN(new_n565));
  OR2_X1    g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n564), .A2(new_n565), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n561), .A2(new_n562), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n393), .A2(new_n297), .ZN(new_n569));
  NAND2_X1  g0369(.A1(KEYINPUT22), .A2(G87), .ZN(new_n570));
  NOR3_X1   g0370(.A1(new_n569), .A2(G20), .A3(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(KEYINPUT24), .B1(new_n568), .B2(new_n571), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n562), .A2(new_n566), .A3(new_n567), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT24), .ZN(new_n574));
  INV_X1    g0374(.A(new_n570), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n428), .A2(new_n205), .A3(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n573), .A2(new_n574), .A3(new_n576), .A4(new_n561), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n265), .B1(new_n572), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n374), .A2(new_n359), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT25), .ZN(new_n580));
  XNOR2_X1  g0380(.A(new_n579), .B(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n485), .A2(G107), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n558), .A2(new_n578), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n557), .A2(new_n280), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n585), .B(KEYINPUT87), .C1(G190), .C2(new_n557), .ZN(new_n586));
  INV_X1    g0386(.A(new_n583), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n572), .A2(new_n577), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n587), .B1(new_n588), .B2(new_n265), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n555), .A2(new_n393), .A3(new_n297), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n402), .A2(G294), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n292), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n552), .ZN(new_n593));
  NOR3_X1   g0393(.A1(new_n592), .A2(new_n593), .A3(new_n509), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n501), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n557), .A2(new_n314), .ZN(new_n596));
  AND2_X1   g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n584), .A2(new_n586), .B1(new_n589), .B2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n511), .ZN(new_n599));
  AND2_X1   g0399(.A1(new_n521), .A2(new_n293), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n599), .B1(new_n600), .B2(new_n529), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(G190), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n524), .A2(G200), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n602), .A2(new_n547), .A3(new_n549), .A4(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(G238), .A2(G1698), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n605), .B1(new_n222), .B2(G1698), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n606), .A2(new_n393), .A3(new_n297), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n402), .A2(G116), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n292), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n459), .A2(new_n281), .ZN(new_n610));
  INV_X1    g0410(.A(G250), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n611), .B1(new_n286), .B2(G1), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n610), .A2(new_n436), .A3(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n609), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(KEYINPUT81), .B1(new_n615), .B2(new_n501), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT81), .ZN(new_n617));
  NOR4_X1   g0417(.A1(new_n609), .A2(new_n617), .A3(G179), .A4(new_n614), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n369), .A2(new_n267), .ZN(new_n620));
  AOI21_X1  g0420(.A(KEYINPUT19), .B1(new_n259), .B2(G97), .ZN(new_n621));
  OR2_X1    g0421(.A1(KEYINPUT82), .A2(G87), .ZN(new_n622));
  NAND2_X1  g0422(.A1(KEYINPUT82), .A2(G87), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n622), .A2(new_n538), .A3(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT19), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n625), .B1(new_n334), .B2(new_n205), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n621), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n393), .A2(new_n205), .A3(G68), .A4(new_n297), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n620), .B1(new_n629), .B2(new_n264), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n485), .A2(new_n369), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n428), .A2(new_n606), .B1(G116), .B2(new_n402), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n613), .B1(new_n632), .B2(new_n292), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n630), .A2(new_n631), .B1(new_n633), .B2(new_n314), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n629), .A2(new_n264), .ZN(new_n635));
  INV_X1    g0435(.A(new_n620), .ZN(new_n636));
  INV_X1    g0436(.A(G87), .ZN(new_n637));
  NOR3_X1   g0437(.A1(new_n268), .A2(new_n637), .A3(new_n484), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n635), .A2(new_n636), .A3(new_n639), .ZN(new_n640));
  NOR3_X1   g0440(.A1(new_n609), .A2(new_n279), .A3(new_n614), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(G200), .B1(new_n609), .B2(new_n614), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n619), .A2(new_n634), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n551), .A2(new_n598), .A3(new_n604), .A4(new_n644), .ZN(new_n645));
  NOR4_X1   g0445(.A1(new_n382), .A2(new_n454), .A3(new_n507), .A4(new_n645), .ZN(G372));
  NOR2_X1   g0446(.A1(new_n382), .A2(new_n454), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n547), .A2(new_n549), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n648), .B1(new_n601), .B2(G169), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n649), .B1(new_n532), .B2(new_n525), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT89), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n650), .A2(new_n651), .A3(KEYINPUT26), .A4(new_n644), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n615), .A2(new_n501), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n634), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n633), .A2(KEYINPUT88), .A3(G200), .ZN(new_n655));
  AOI211_X1 g0455(.A(new_n620), .B(new_n638), .C1(new_n629), .C2(new_n264), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT88), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n643), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n641), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n655), .A2(new_n656), .A3(new_n658), .A4(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n654), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(KEYINPUT26), .B1(new_n650), .B2(new_n662), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n533), .A2(new_n644), .A3(KEYINPUT26), .A4(new_n550), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(KEYINPUT89), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n652), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n661), .B1(new_n586), .B2(new_n584), .ZN(new_n667));
  OAI211_X1 g0467(.A(new_n596), .B(new_n595), .C1(new_n578), .C2(new_n583), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n506), .A2(new_n668), .A3(new_n499), .A4(new_n503), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n667), .A2(new_n669), .A3(new_n551), .A4(new_n604), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n654), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n666), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n647), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n386), .ZN(new_n674));
  INV_X1    g0474(.A(new_n398), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n320), .B1(new_n394), .B2(new_n395), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n421), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n265), .B1(new_n677), .B2(KEYINPUT16), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n674), .B1(new_n678), .B2(new_n422), .ZN(new_n679));
  INV_X1    g0479(.A(new_n440), .ZN(new_n680));
  OAI21_X1  g0480(.A(KEYINPUT18), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n680), .B1(new_n423), .B2(new_n386), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(new_n443), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n354), .B1(new_n345), .B2(new_n377), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n686), .B(KEYINPUT90), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n685), .B1(new_n687), .B2(new_n452), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n316), .B1(new_n688), .B2(new_n311), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n673), .A2(new_n689), .ZN(G369));
  NAND3_X1  g0490(.A1(new_n506), .A2(new_n499), .A3(new_n503), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n204), .A2(new_n205), .A3(G13), .ZN(new_n692));
  OR2_X1    g0492(.A1(new_n692), .A2(KEYINPUT27), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(KEYINPUT27), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n693), .A2(G213), .A3(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(G343), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n495), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n691), .A2(new_n699), .ZN(new_n700));
  OAI211_X1 g0500(.A(KEYINPUT91), .B(new_n700), .C1(new_n507), .C2(new_n699), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n700), .A2(KEYINPUT91), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n701), .A2(new_n702), .A3(G330), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n589), .A2(new_n697), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n578), .A2(new_n583), .ZN(new_n706));
  INV_X1    g0506(.A(new_n558), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n706), .A2(new_n586), .A3(new_n707), .ZN(new_n708));
  AOI22_X1  g0508(.A1(new_n705), .A2(new_n708), .B1(new_n589), .B2(new_n597), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n668), .A2(new_n697), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n704), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n691), .A2(new_n698), .ZN(new_n713));
  NOR3_X1   g0513(.A1(new_n713), .A2(new_n710), .A3(new_n709), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(new_n710), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n712), .A2(new_n715), .ZN(G399));
  NOR2_X1   g0516(.A1(new_n624), .A2(G116), .ZN(new_n717));
  XNOR2_X1  g0517(.A(new_n717), .B(KEYINPUT92), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n208), .A2(new_n285), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(G1), .ZN(new_n720));
  OAI22_X1  g0520(.A1(new_n718), .A2(new_n720), .B1(new_n218), .B2(new_n719), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT28), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n650), .A2(KEYINPUT95), .A3(KEYINPUT26), .A4(new_n662), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n670), .A2(new_n723), .A3(new_n654), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n662), .A2(new_n533), .A3(KEYINPUT26), .A4(new_n550), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT95), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(KEYINPUT26), .B1(new_n650), .B2(new_n644), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n724), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(KEYINPUT29), .B1(new_n730), .B2(new_n697), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n672), .A2(new_n698), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n731), .B1(new_n732), .B2(KEYINPUT29), .ZN(new_n733));
  INV_X1    g0533(.A(G330), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n645), .A2(new_n507), .A3(new_n697), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT31), .ZN(new_n736));
  INV_X1    g0536(.A(new_n468), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n471), .B1(new_n737), .B2(new_n470), .ZN(new_n738));
  INV_X1    g0538(.A(new_n472), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n502), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(KEYINPUT93), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT93), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n500), .A2(new_n742), .A3(new_n502), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n592), .A2(new_n593), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n530), .A2(new_n511), .A3(new_n615), .A4(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n741), .A2(new_n743), .A3(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT30), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n557), .A2(new_n633), .A3(new_n501), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n749), .B1(new_n530), .B2(new_n511), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n748), .B1(new_n750), .B2(new_n505), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n697), .B1(new_n747), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n501), .B1(new_n609), .B2(new_n614), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n594), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n524), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(KEYINPUT30), .B1(new_n755), .B2(new_n482), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n745), .B1(KEYINPUT93), .B2(new_n740), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n756), .B1(new_n743), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n736), .B1(new_n752), .B2(new_n758), .ZN(new_n759));
  AND3_X1   g0559(.A1(new_n500), .A2(new_n742), .A3(new_n502), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n742), .B1(new_n500), .B2(new_n502), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n760), .A2(new_n761), .A3(new_n745), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(new_n756), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n747), .A2(new_n751), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n763), .A2(new_n764), .A3(KEYINPUT31), .A4(new_n697), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n759), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n735), .B1(new_n766), .B2(KEYINPUT94), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT94), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n759), .A2(new_n765), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n734), .B1(new_n767), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n733), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n722), .B1(new_n771), .B2(G1), .ZN(G364));
  NAND2_X1  g0572(.A1(new_n704), .A2(KEYINPUT96), .ZN(new_n773));
  INV_X1    g0573(.A(KEYINPUT96), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n703), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n719), .ZN(new_n776));
  INV_X1    g0576(.A(G13), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(G20), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n204), .B1(new_n778), .B2(G45), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n776), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n701), .A2(new_n702), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n781), .B1(new_n782), .B2(new_n734), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n773), .A2(new_n775), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n216), .B1(G20), .B2(new_n314), .ZN(new_n785));
  OR2_X1    g0585(.A1(new_n785), .A2(KEYINPUT97), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(KEYINPUT97), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(G13), .A2(G33), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(G20), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n208), .A2(G355), .A3(new_n299), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n794), .B1(G116), .B2(new_n208), .ZN(new_n795));
  OR2_X1    g0595(.A1(new_n245), .A2(new_n286), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n208), .A2(new_n569), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n797), .B1(new_n286), .B2(new_n219), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n795), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n781), .B1(new_n793), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n205), .A2(new_n279), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n501), .A2(G200), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(G322), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n205), .A2(G190), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(new_n802), .ZN(new_n806));
  INV_X1    g0606(.A(G311), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n803), .A2(new_n804), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n801), .ZN(new_n809));
  NOR3_X1   g0609(.A1(new_n809), .A2(new_n280), .A3(G179), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n299), .B(new_n808), .C1(G303), .C2(new_n810), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n805), .A2(new_n501), .A3(G200), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(G283), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n205), .A2(new_n501), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n815), .A2(new_n279), .A3(G200), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  XNOR2_X1  g0617(.A(KEYINPUT33), .B(G317), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n805), .A2(new_n501), .A3(new_n280), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n817), .A2(new_n818), .B1(new_n820), .B2(G329), .ZN(new_n821));
  NOR3_X1   g0621(.A1(new_n279), .A2(G179), .A3(G200), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(new_n205), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NOR4_X1   g0624(.A1(new_n205), .A2(new_n501), .A3(new_n279), .A4(new_n280), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n824), .A2(G294), .B1(new_n825), .B2(G326), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n811), .A2(new_n814), .A3(new_n821), .A4(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n810), .ZN(new_n828));
  AND2_X1   g0628(.A1(new_n622), .A2(new_n623), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n299), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n830), .B(KEYINPUT99), .Z(new_n831));
  NAND2_X1  g0631(.A1(new_n820), .A2(G159), .ZN(new_n832));
  XOR2_X1   g0632(.A(new_n803), .B(KEYINPUT98), .Z(new_n833));
  OAI221_X1 g0633(.A(new_n831), .B1(KEYINPUT32), .B2(new_n832), .C1(new_n387), .C2(new_n833), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n824), .A2(G97), .B1(new_n825), .B2(G50), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n832), .A2(KEYINPUT32), .ZN(new_n836));
  INV_X1    g0636(.A(new_n806), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n817), .A2(G68), .B1(new_n837), .B2(new_n294), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n812), .A2(new_n359), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n835), .A2(new_n836), .A3(new_n838), .A4(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n827), .B1(new_n834), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n800), .B1(new_n842), .B2(new_n788), .ZN(new_n843));
  INV_X1    g0643(.A(new_n782), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n791), .B(KEYINPUT100), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n843), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n784), .A2(new_n846), .ZN(G396));
  INV_X1    g0647(.A(new_n781), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n788), .A2(new_n789), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n848), .B1(new_n849), .B2(new_n365), .ZN(new_n850));
  INV_X1    g0650(.A(new_n788), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n813), .A2(G87), .B1(new_n820), .B2(G311), .ZN(new_n852));
  INV_X1    g0652(.A(G283), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n852), .B1(new_n853), .B2(new_n816), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n828), .A2(new_n359), .B1(new_n803), .B2(new_n553), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n298), .B1(new_n806), .B2(new_n487), .ZN(new_n856));
  INV_X1    g0656(.A(new_n825), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n857), .A2(new_n475), .B1(new_n536), .B2(new_n823), .ZN(new_n858));
  NOR4_X1   g0658(.A1(new_n854), .A2(new_n855), .A3(new_n856), .A4(new_n858), .ZN(new_n859));
  AOI22_X1  g0659(.A1(G137), .A2(new_n825), .B1(new_n837), .B2(G159), .ZN(new_n860));
  INV_X1    g0660(.A(G143), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n860), .B1(new_n251), .B2(new_n816), .C1(new_n833), .C2(new_n861), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n862), .B(KEYINPUT34), .ZN(new_n863));
  INV_X1    g0663(.A(G132), .ZN(new_n864));
  OAI22_X1  g0664(.A1(new_n320), .A2(new_n812), .B1(new_n819), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(G50), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n428), .B1(new_n828), .B2(new_n866), .ZN(new_n867));
  AOI211_X1 g0667(.A(new_n865), .B(new_n867), .C1(new_n256), .C2(new_n824), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n859), .B1(new_n863), .B2(new_n868), .ZN(new_n869));
  OR2_X1    g0669(.A1(new_n377), .A2(new_n697), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n376), .A2(new_n697), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(new_n379), .B2(new_n380), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n377), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  OAI221_X1 g0675(.A(new_n850), .B1(new_n851), .B2(new_n869), .C1(new_n875), .C2(new_n790), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  XNOR2_X1  g0677(.A(new_n732), .B(new_n875), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n878), .A2(new_n770), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n879), .A2(new_n781), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n878), .A2(new_n770), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n877), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(G384));
  NOR2_X1   g0683(.A1(new_n778), .A2(new_n204), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT38), .ZN(new_n885));
  OR2_X1    g0685(.A1(new_n677), .A2(KEYINPUT16), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n674), .B1(new_n886), .B2(new_n678), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n887), .A2(new_n695), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n452), .B1(KEYINPUT18), .B2(new_n441), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n889), .B1(new_n890), .B2(new_n444), .ZN(new_n891));
  XOR2_X1   g0691(.A(new_n695), .B(KEYINPUT101), .Z(new_n892));
  NAND3_X1  g0692(.A1(new_n413), .A2(new_n425), .A3(new_n892), .ZN(new_n893));
  AND3_X1   g0693(.A1(new_n423), .A2(new_n386), .A3(new_n447), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n894), .A2(KEYINPUT37), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n441), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n448), .B1(new_n887), .B2(new_n695), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n887), .A2(new_n680), .ZN(new_n898));
  OAI21_X1  g0698(.A(KEYINPUT37), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n885), .B1(new_n891), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n454), .A2(new_n888), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n896), .A2(new_n899), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n902), .A2(KEYINPUT38), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT40), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n495), .B1(new_n482), .B2(new_n280), .ZN(new_n907));
  AND3_X1   g0707(.A1(new_n500), .A2(G190), .A3(new_n504), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n691), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n648), .B1(G200), .B2(new_n524), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n602), .A2(new_n911), .B1(new_n533), .B2(new_n550), .ZN(new_n912));
  AND3_X1   g0712(.A1(new_n644), .A2(new_n708), .A3(new_n668), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n910), .A2(new_n912), .A3(new_n913), .A4(new_n698), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n914), .A2(new_n759), .A3(new_n765), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n330), .A2(new_n697), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n346), .A2(new_n354), .A3(new_n916), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n330), .B(new_n697), .C1(new_n345), .C2(new_n353), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n874), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  AND2_X1   g0719(.A1(new_n915), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n905), .A2(new_n906), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n915), .A2(new_n919), .ZN(new_n922));
  INV_X1    g0722(.A(new_n893), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n684), .B2(new_n452), .ZN(new_n924));
  AND3_X1   g0724(.A1(new_n441), .A2(new_n893), .A3(new_n895), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT37), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n894), .A2(new_n682), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n926), .B1(new_n893), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n924), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n885), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n922), .B1(new_n904), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n921), .B1(new_n931), .B2(new_n906), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT102), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n647), .A2(new_n915), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n734), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n934), .B2(new_n933), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n647), .A2(new_n733), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n689), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT39), .ZN(new_n939));
  AOI221_X4 g0739(.A(new_n885), .B1(new_n896), .B2(new_n899), .C1(new_n454), .C2(new_n888), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n893), .A2(new_n927), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n896), .B1(new_n941), .B2(new_n926), .ZN(new_n942));
  AOI21_X1  g0742(.A(KEYINPUT38), .B1(new_n942), .B2(new_n924), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n939), .B1(new_n940), .B2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n353), .A2(new_n330), .A3(new_n698), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n901), .A2(KEYINPUT39), .A3(new_n904), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n944), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n917), .A2(new_n918), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n698), .B(new_n875), .C1(new_n666), .C2(new_n671), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n950), .B1(new_n951), .B2(new_n870), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n905), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n685), .A2(new_n892), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n948), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n938), .B(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n884), .B1(new_n936), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n956), .B2(new_n936), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n544), .A2(KEYINPUT35), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n544), .A2(KEYINPUT35), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n959), .A2(G116), .A3(new_n217), .A4(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT36), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n219), .B(new_n294), .C1(new_n320), .C2(new_n387), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(G50), .B2(new_n320), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n964), .A2(G1), .A3(new_n777), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n958), .A2(new_n962), .A3(new_n965), .ZN(G367));
  OAI21_X1  g0766(.A(new_n792), .B1(new_n208), .B2(new_n368), .ZN(new_n967));
  AND3_X1   g0767(.A1(new_n236), .A2(new_n208), .A3(new_n569), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n969), .A2(new_n848), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n640), .A2(new_n697), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n662), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n654), .B2(new_n971), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n823), .A2(new_n320), .B1(new_n803), .B2(new_n251), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT108), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n299), .B1(new_n806), .B2(new_n866), .C1(new_n828), .C2(new_n387), .ZN(new_n976));
  INV_X1    g0776(.A(G159), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n857), .A2(new_n861), .B1(new_n977), .B2(new_n816), .ZN(new_n978));
  INV_X1    g0778(.A(G137), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n221), .A2(new_n812), .B1(new_n819), .B2(new_n979), .ZN(new_n980));
  OR4_X1    g0780(.A1(new_n975), .A2(new_n976), .A3(new_n978), .A4(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n810), .A2(G116), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(KEYINPUT46), .Z(new_n983));
  AOI211_X1 g0783(.A(new_n428), .B(new_n983), .C1(G283), .C2(new_n837), .ZN(new_n984));
  INV_X1    g0784(.A(new_n833), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n985), .A2(G303), .B1(G311), .B2(new_n825), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(KEYINPUT107), .ZN(new_n988));
  AOI22_X1  g0788(.A1(G107), .A2(new_n824), .B1(new_n817), .B2(G294), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n813), .A2(G97), .B1(new_n820), .B2(G317), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n984), .A2(new_n988), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n987), .A2(KEYINPUT107), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n981), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT47), .ZN(new_n994));
  AND2_X1   g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n788), .B1(new_n993), .B2(new_n994), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n970), .B1(new_n845), .B2(new_n973), .C1(new_n995), .C2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT105), .ZN(new_n998));
  INV_X1    g0798(.A(new_n712), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n648), .A2(new_n697), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n912), .A2(new_n1000), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n1001), .A2(KEYINPUT103), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n650), .A2(new_n697), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1001), .A2(KEYINPUT103), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n999), .A2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n973), .A2(KEYINPUT43), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n668), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n698), .B1(new_n1008), .B2(new_n650), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1005), .A2(KEYINPUT42), .A3(new_n714), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(KEYINPUT42), .B1(new_n1005), .B2(new_n714), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1007), .B(new_n1009), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT104), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1012), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n1010), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1017), .A2(KEYINPUT104), .A3(new_n1007), .A4(new_n1009), .ZN(new_n1018));
  AND2_X1   g0818(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1017), .A2(new_n1009), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n973), .B(KEYINPUT43), .Z(new_n1021));
  AND2_X1   g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n998), .B(new_n1006), .C1(new_n1019), .C2(new_n1022), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n1015), .A2(new_n1018), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1006), .ZN(new_n1025));
  OAI21_X1  g0825(.A(KEYINPUT105), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1023), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT44), .ZN(new_n1029));
  OR3_X1    g0829(.A1(new_n1005), .A2(new_n1029), .A3(new_n715), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1029), .B1(new_n1005), .B2(new_n715), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1005), .A2(new_n715), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT45), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1005), .A2(KEYINPUT45), .A3(new_n715), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1032), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(new_n999), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1032), .A2(new_n1037), .A3(new_n712), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n773), .A2(KEYINPUT106), .A3(new_n775), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n711), .B(new_n713), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1043), .B(new_n703), .C1(new_n774), .C2(KEYINPUT106), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(new_n771), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n771), .B1(new_n1041), .B2(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n719), .B(KEYINPUT41), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n780), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n997), .B1(new_n1028), .B2(new_n1052), .ZN(G387));
  INV_X1    g0853(.A(new_n771), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1054), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1055), .A2(new_n776), .A3(new_n1048), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n718), .A2(new_n208), .A3(new_n299), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(G107), .B2(new_n208), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n371), .A2(new_n866), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT50), .ZN(new_n1060));
  AOI211_X1 g0860(.A(G45), .B(new_n718), .C1(G68), .C2(G77), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1060), .B1(new_n1061), .B2(KEYINPUT109), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(KEYINPUT109), .B2(new_n1061), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n797), .B1(new_n241), .B2(G45), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1058), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n781), .B1(new_n1065), .B2(new_n793), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT110), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n817), .A2(G311), .B1(new_n837), .B2(G303), .ZN(new_n1068));
  INV_X1    g0868(.A(G317), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1068), .B1(new_n804), .B2(new_n857), .C1(new_n833), .C2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT48), .ZN(new_n1071));
  OR2_X1    g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n828), .A2(new_n553), .B1(new_n853), .B2(new_n823), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT112), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1072), .A2(new_n1073), .A3(new_n1075), .ZN(new_n1076));
  XOR2_X1   g0876(.A(new_n1076), .B(KEYINPUT113), .Z(new_n1077));
  OR2_X1    g0877(.A1(new_n1077), .A2(KEYINPUT49), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1077), .A2(KEYINPUT49), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n569), .B1(new_n487), .B2(new_n812), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(G326), .B2(new_n820), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1078), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n823), .A2(new_n368), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n803), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1083), .B1(G50), .B2(new_n1084), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT111), .Z(new_n1086));
  OAI22_X1  g0886(.A1(new_n536), .A2(new_n812), .B1(new_n819), .B2(new_n251), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(G159), .B2(new_n825), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n810), .A2(new_n294), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1089), .B(new_n428), .C1(new_n320), .C2(new_n806), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n257), .B2(new_n817), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1086), .A2(new_n1088), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1082), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1067), .B1(new_n1093), .B2(new_n788), .ZN(new_n1094));
  OR2_X1    g0894(.A1(new_n1094), .A2(KEYINPUT114), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n711), .A2(new_n845), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n1094), .B2(KEYINPUT114), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1047), .A2(new_n780), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(KEYINPUT115), .B1(new_n1056), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1056), .A2(KEYINPUT115), .A3(new_n1098), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(new_n1101), .ZN(G393));
  INV_X1    g0902(.A(new_n1040), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n712), .B1(new_n1032), .B2(new_n1037), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1002), .A2(new_n791), .A3(new_n1003), .A4(new_n1004), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n248), .A2(new_n797), .B1(new_n536), .B2(new_n208), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n781), .B1(new_n793), .B2(new_n1107), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n298), .B1(new_n806), .B2(new_n553), .C1(new_n828), .C2(new_n853), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n839), .B(new_n1109), .C1(G322), .C2(new_n820), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n823), .A2(new_n487), .B1(new_n816), .B2(new_n475), .ZN(new_n1111));
  XOR2_X1   g0911(.A(new_n1111), .B(KEYINPUT116), .Z(new_n1112));
  OAI22_X1  g0912(.A1(new_n857), .A2(new_n1069), .B1(new_n803), .B2(new_n807), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT52), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1110), .A2(new_n1112), .A3(new_n1114), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n857), .A2(new_n251), .B1(new_n803), .B2(new_n977), .ZN(new_n1116));
  XOR2_X1   g0916(.A(new_n1116), .B(KEYINPUT51), .Z(new_n1117));
  OAI22_X1  g0917(.A1(new_n823), .A2(new_n365), .B1(new_n812), .B2(new_n637), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n816), .A2(new_n866), .B1(new_n819), .B2(new_n861), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n810), .A2(G68), .B1(new_n371), .B2(new_n837), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1120), .A2(new_n428), .A3(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1115), .B1(new_n1117), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1108), .B1(new_n1123), .B2(new_n788), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n1105), .A2(new_n780), .B1(new_n1106), .B2(new_n1124), .ZN(new_n1125));
  AND2_X1   g0925(.A1(new_n1041), .A2(new_n1048), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n776), .B1(new_n1041), .B2(new_n1048), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1125), .B1(new_n1126), .B2(new_n1127), .ZN(G390));
  NAND3_X1  g0928(.A1(new_n770), .A2(new_n875), .A3(new_n949), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n915), .A2(G330), .ZN(new_n1130));
  AND3_X1   g0930(.A1(new_n917), .A2(KEYINPUT117), .A3(new_n918), .ZN(new_n1131));
  AOI21_X1  g0931(.A(KEYINPUT117), .B1(new_n917), .B2(new_n918), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n1130), .A2(new_n874), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n698), .B(new_n873), .C1(new_n724), .C2(new_n729), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n870), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  AND3_X1   g0936(.A1(new_n1129), .A2(new_n1133), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  AND3_X1   g0938(.A1(new_n915), .A2(new_n919), .A3(G330), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n734), .B(new_n874), .C1(new_n767), .C2(new_n769), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1140), .B1(new_n1141), .B2(new_n949), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n951), .A2(new_n870), .ZN(new_n1143));
  AOI21_X1  g0943(.A(KEYINPUT118), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n698), .B1(new_n762), .B2(new_n756), .ZN(new_n1145));
  AOI21_X1  g0945(.A(KEYINPUT31), .B1(new_n1145), .B2(new_n764), .ZN(new_n1146));
  NOR3_X1   g0946(.A1(new_n752), .A2(new_n758), .A3(new_n736), .ZN(new_n1147));
  OAI21_X1  g0947(.A(KEYINPUT94), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1148), .A2(new_n769), .A3(new_n914), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1149), .A2(G330), .A3(new_n875), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1139), .B1(new_n1150), .B2(new_n950), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT118), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1143), .ZN(new_n1153));
  NOR3_X1   g0953(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1138), .B1(new_n1144), .B2(new_n1154), .ZN(new_n1155));
  AND3_X1   g0955(.A1(new_n901), .A2(KEYINPUT39), .A3(new_n904), .ZN(new_n1156));
  AOI21_X1  g0956(.A(KEYINPUT39), .B1(new_n904), .B2(new_n930), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n1156), .A2(new_n1157), .B1(new_n952), .B2(new_n946), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1135), .A2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n946), .B1(new_n904), .B2(new_n930), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1140), .B1(new_n1158), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1143), .A2(new_n949), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n945), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n944), .A2(new_n947), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n1165), .A2(new_n1166), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1163), .B1(new_n1167), .B2(new_n1129), .ZN(new_n1168));
  AND2_X1   g0968(.A1(new_n915), .A2(G330), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n647), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n937), .A2(new_n1170), .A3(new_n689), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1155), .A2(new_n1168), .A3(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1158), .A2(new_n1162), .A3(new_n1129), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n1167), .B2(new_n1140), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1152), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n949), .B1(new_n770), .B2(new_n875), .ZN(new_n1177));
  OAI211_X1 g0977(.A(KEYINPUT118), .B(new_n1143), .C1(new_n1177), .C2(new_n1139), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1137), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1175), .B1(new_n1179), .B2(new_n1171), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1173), .A2(new_n1180), .A3(new_n776), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1166), .A2(new_n789), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n810), .A2(G150), .ZN(new_n1183));
  XOR2_X1   g0983(.A(new_n1183), .B(KEYINPUT53), .Z(new_n1184));
  INV_X1    g0984(.A(G128), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n857), .A2(new_n1185), .B1(new_n977), .B2(new_n823), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(G137), .B2(new_n817), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(KEYINPUT54), .B(G143), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n806), .A2(new_n1188), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n298), .B(new_n1189), .C1(G132), .C2(new_n1084), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n813), .A2(G50), .B1(new_n820), .B2(G125), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1184), .A2(new_n1187), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n857), .A2(new_n853), .B1(new_n359), .B2(new_n816), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(G294), .B2(new_n820), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n299), .B1(new_n810), .B2(G87), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(G116), .A2(new_n1084), .B1(new_n837), .B2(G97), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n824), .A2(G77), .B1(new_n813), .B2(G68), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .A4(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n851), .B1(new_n1192), .B2(new_n1198), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n848), .B(new_n1199), .C1(new_n383), .C2(new_n849), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n1168), .A2(new_n780), .B1(new_n1182), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1181), .A2(new_n1201), .ZN(G378));
  INV_X1    g1002(.A(KEYINPUT57), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1171), .B1(new_n1155), .B2(new_n1168), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n904), .A2(new_n930), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n906), .B1(new_n1205), .B2(new_n920), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n915), .A2(new_n919), .A3(new_n906), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(new_n904), .B2(new_n901), .ZN(new_n1208));
  OAI21_X1  g1008(.A(G330), .B1(new_n1206), .B2(new_n1208), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n272), .A2(new_n695), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n318), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1210), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n311), .A2(new_n317), .A3(new_n1212), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1211), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1214), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1212), .B1(new_n311), .B2(new_n317), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n316), .B(new_n1210), .C1(new_n308), .C2(new_n310), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1216), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1215), .A2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1209), .A2(new_n1221), .ZN(new_n1222));
  AND3_X1   g1022(.A1(new_n948), .A2(new_n953), .A3(new_n954), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1220), .B(G330), .C1(new_n1206), .C2(new_n1208), .ZN(new_n1224));
  AND3_X1   g1024(.A1(new_n1222), .A2(new_n1223), .A3(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1223), .B1(new_n1222), .B2(new_n1224), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1203), .B1(new_n1204), .B2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1220), .B1(new_n932), .B2(G330), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1224), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n955), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1222), .A2(new_n1223), .A3(new_n1224), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1203), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1172), .B1(new_n1179), .B2(new_n1175), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n719), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1228), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT121), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n779), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1221), .A2(new_n789), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n848), .B1(new_n849), .B2(new_n866), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1240), .B(KEYINPUT120), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n428), .A2(G41), .ZN(new_n1242));
  AOI211_X1 g1042(.A(G50), .B(new_n1242), .C1(new_n258), .C2(new_n285), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1089), .B1(new_n359), .B2(new_n803), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(new_n369), .B2(new_n837), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n857), .A2(new_n487), .B1(new_n853), .B2(new_n819), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(G97), .B2(new_n817), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n824), .A2(G68), .B1(new_n813), .B2(new_n256), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1245), .A2(new_n1247), .A3(new_n1242), .A4(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT58), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1243), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n828), .A2(new_n1188), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n1253), .A2(KEYINPUT119), .B1(G125), .B2(new_n825), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(G150), .A2(new_n824), .B1(new_n817), .B2(G132), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1253), .A2(KEYINPUT119), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n803), .A2(new_n1185), .B1(new_n806), .B2(new_n979), .ZN(new_n1258));
  NOR3_X1   g1058(.A1(new_n1256), .A2(new_n1257), .A3(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1260), .A2(KEYINPUT59), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n258), .B(new_n285), .C1(new_n812), .C2(new_n977), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1262), .B1(G124), .B2(new_n820), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT59), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1263), .B1(new_n1259), .B2(new_n1264), .ZN(new_n1265));
  OAI221_X1 g1065(.A(new_n1251), .B1(new_n1250), .B2(new_n1249), .C1(new_n1261), .C2(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1241), .B1(new_n1266), .B2(new_n788), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1239), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1237), .B1(new_n1238), .B2(new_n1269), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n780), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1271), .A2(KEYINPUT121), .A3(new_n1268), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1270), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1236), .A2(new_n1273), .ZN(G375));
  NAND2_X1  g1074(.A1(new_n1155), .A2(new_n1172), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1179), .A2(new_n1171), .ZN(new_n1276));
  XOR2_X1   g1076(.A(new_n1050), .B(KEYINPUT122), .Z(new_n1277));
  NAND3_X1  g1077(.A1(new_n1275), .A2(new_n1276), .A3(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n848), .B1(new_n849), .B2(new_n320), .ZN(new_n1279));
  OAI22_X1  g1079(.A1(new_n857), .A2(new_n864), .B1(new_n816), .B2(new_n1188), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1280), .B1(G50), .B2(new_n824), .ZN(new_n1281));
  OAI22_X1  g1081(.A1(new_n1185), .A2(new_n819), .B1(new_n812), .B2(new_n387), .ZN(new_n1282));
  OAI221_X1 g1082(.A(new_n428), .B1(new_n251), .B2(new_n806), .C1(new_n828), .C2(new_n977), .ZN(new_n1283));
  AOI211_X1 g1083(.A(new_n1282), .B(new_n1283), .C1(G137), .C2(new_n985), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n299), .B1(new_n1084), .B2(G283), .ZN(new_n1285));
  OAI221_X1 g1085(.A(new_n1285), .B1(new_n359), .B2(new_n806), .C1(new_n828), .C2(new_n536), .ZN(new_n1286));
  AOI211_X1 g1086(.A(new_n1083), .B(new_n1286), .C1(G294), .C2(new_n825), .ZN(new_n1287));
  OAI22_X1  g1087(.A1(new_n816), .A2(new_n487), .B1(new_n819), .B2(new_n475), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1288), .B1(G77), .B2(new_n813), .ZN(new_n1289));
  AOI22_X1  g1089(.A1(new_n1281), .A2(new_n1284), .B1(new_n1287), .B2(new_n1289), .ZN(new_n1290));
  OAI221_X1 g1090(.A(new_n1279), .B1(new_n851), .B2(new_n1290), .C1(new_n1159), .C2(new_n790), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1291), .B1(new_n1179), .B2(new_n779), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1278), .A2(new_n1293), .ZN(G381));
  AND3_X1   g1094(.A1(new_n1181), .A2(KEYINPUT123), .A3(new_n1201), .ZN(new_n1295));
  AOI21_X1  g1095(.A(KEYINPUT123), .B1(new_n1181), .B2(new_n1201), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1297), .A2(new_n1236), .A3(new_n1273), .ZN(new_n1298));
  INV_X1    g1098(.A(G396), .ZN(new_n1299));
  AND3_X1   g1099(.A1(new_n1100), .A2(new_n1299), .A3(new_n1101), .ZN(new_n1300));
  INV_X1    g1100(.A(G390), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1300), .A2(new_n882), .A3(new_n1301), .ZN(new_n1302));
  OR4_X1    g1102(.A1(G387), .A2(new_n1298), .A3(G381), .A4(new_n1302), .ZN(G407));
  OAI211_X1 g1103(.A(G407), .B(G213), .C1(G343), .C2(new_n1298), .ZN(G409));
  INV_X1    g1104(.A(KEYINPUT125), .ZN(new_n1305));
  OAI211_X1 g1105(.A(new_n997), .B(G390), .C1(new_n1028), .C2(new_n1052), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1299), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1306), .B1(new_n1300), .B2(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1054), .B1(new_n1105), .B2(new_n1047), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n779), .B1(new_n1309), .B2(new_n1050), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1310), .A2(new_n1023), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1311));
  AOI21_X1  g1111(.A(G390), .B1(new_n1311), .B2(new_n997), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1305), .B1(new_n1308), .B2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1307), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1100), .A2(new_n1299), .A3(new_n1101), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(G387), .A2(new_n1301), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1316), .A2(new_n1317), .A3(KEYINPUT125), .A4(new_n1306), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1311), .A2(KEYINPUT124), .A3(new_n997), .A4(G390), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT124), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1306), .A2(new_n1320), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1319), .A2(new_n1321), .A3(new_n1317), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1316), .ZN(new_n1323));
  AOI22_X1  g1123(.A1(new_n1313), .A2(new_n1318), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n696), .A2(G213), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1326), .A2(KEYINPUT60), .A3(new_n1171), .A4(new_n1138), .ZN(new_n1327));
  AND2_X1   g1127(.A1(new_n1327), .A2(new_n776), .ZN(new_n1328));
  OAI21_X1  g1128(.A(KEYINPUT60), .B1(new_n1179), .B2(new_n1171), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1329), .A2(new_n1276), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1328), .A2(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(G384), .B1(new_n1331), .B2(new_n1293), .ZN(new_n1332));
  AOI211_X1 g1132(.A(new_n882), .B(new_n1292), .C1(new_n1328), .C2(new_n1330), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1332), .A2(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1234), .A2(new_n1335), .A3(new_n1277), .ZN(new_n1336));
  AOI21_X1  g1136(.A(new_n1269), .B1(new_n1335), .B2(new_n780), .ZN(new_n1337));
  AND2_X1   g1137(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1338));
  NOR3_X1   g1138(.A1(new_n1295), .A2(new_n1296), .A3(new_n1338), .ZN(new_n1339));
  AND3_X1   g1139(.A1(new_n1236), .A2(G378), .A3(new_n1273), .ZN(new_n1340));
  OAI211_X1 g1140(.A(new_n1325), .B(new_n1334), .C1(new_n1339), .C2(new_n1340), .ZN(new_n1341));
  INV_X1    g1141(.A(KEYINPUT62), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1236), .A2(G378), .A3(new_n1273), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT123), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(G378), .A2(new_n1345), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1181), .A2(KEYINPUT123), .A3(new_n1201), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1346), .A2(new_n1347), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1344), .B1(new_n1348), .B2(new_n1338), .ZN(new_n1349));
  NAND4_X1  g1149(.A1(new_n1349), .A2(KEYINPUT62), .A3(new_n1325), .A4(new_n1334), .ZN(new_n1350));
  AND3_X1   g1150(.A1(new_n1343), .A2(KEYINPUT126), .A3(new_n1350), .ZN(new_n1351));
  INV_X1    g1151(.A(KEYINPUT126), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1341), .A2(new_n1352), .A3(new_n1342), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT61), .ZN(new_n1354));
  OAI21_X1  g1154(.A(new_n1325), .B1(new_n1339), .B2(new_n1340), .ZN(new_n1355));
  INV_X1    g1155(.A(G2897), .ZN(new_n1356));
  OAI21_X1  g1156(.A(new_n1334), .B1(new_n1356), .B2(new_n1325), .ZN(new_n1357));
  INV_X1    g1157(.A(new_n1325), .ZN(new_n1358));
  OAI211_X1 g1158(.A(G2897), .B(new_n1358), .C1(new_n1332), .C2(new_n1333), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1355), .A2(new_n1357), .A3(new_n1359), .ZN(new_n1360));
  NAND3_X1  g1160(.A1(new_n1353), .A2(new_n1354), .A3(new_n1360), .ZN(new_n1361));
  OAI21_X1  g1161(.A(new_n1324), .B1(new_n1351), .B2(new_n1361), .ZN(new_n1362));
  INV_X1    g1162(.A(KEYINPUT63), .ZN(new_n1363));
  AOI21_X1  g1163(.A(new_n1324), .B1(new_n1363), .B2(new_n1341), .ZN(new_n1364));
  AND2_X1   g1164(.A1(new_n1360), .A2(new_n1354), .ZN(new_n1365));
  OR2_X1    g1165(.A1(new_n1341), .A2(new_n1363), .ZN(new_n1366));
  NAND3_X1  g1166(.A1(new_n1364), .A2(new_n1365), .A3(new_n1366), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1362), .A2(new_n1367), .ZN(G405));
  NAND2_X1  g1168(.A1(new_n1297), .A2(G375), .ZN(new_n1369));
  INV_X1    g1169(.A(KEYINPUT127), .ZN(new_n1370));
  NAND3_X1  g1170(.A1(new_n1369), .A2(new_n1370), .A3(new_n1344), .ZN(new_n1371));
  INV_X1    g1171(.A(new_n1371), .ZN(new_n1372));
  AOI21_X1  g1172(.A(new_n1370), .B1(new_n1369), .B2(new_n1344), .ZN(new_n1373));
  OAI21_X1  g1173(.A(new_n1334), .B1(new_n1372), .B2(new_n1373), .ZN(new_n1374));
  NAND2_X1  g1174(.A1(new_n1369), .A2(new_n1344), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1375), .A2(KEYINPUT127), .ZN(new_n1376));
  INV_X1    g1176(.A(new_n1334), .ZN(new_n1377));
  NAND3_X1  g1177(.A1(new_n1376), .A2(new_n1377), .A3(new_n1371), .ZN(new_n1378));
  NAND2_X1  g1178(.A1(new_n1374), .A2(new_n1378), .ZN(new_n1379));
  AND2_X1   g1179(.A1(new_n1313), .A2(new_n1318), .ZN(new_n1380));
  AND2_X1   g1180(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1381));
  OR2_X1    g1181(.A1(new_n1380), .A2(new_n1381), .ZN(new_n1382));
  NAND2_X1  g1182(.A1(new_n1379), .A2(new_n1382), .ZN(new_n1383));
  NAND3_X1  g1183(.A1(new_n1374), .A2(new_n1324), .A3(new_n1378), .ZN(new_n1384));
  NAND2_X1  g1184(.A1(new_n1383), .A2(new_n1384), .ZN(G402));
endmodule


