//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 1 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 0 0 1 1 1 0 1 1 0 0 1 0 0 0 1 0 1 1 0 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:39 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n565, new_n566,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1194;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT64), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT65), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT67), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n454));
  XNOR2_X1  g029(.A(new_n453), .B(new_n454), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n452), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n452), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n466), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G137), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n469), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  NOR2_X1   g052(.A1(new_n466), .A2(new_n470), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(G112), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n481), .B1(new_n482), .B2(G2105), .ZN(new_n483));
  OR2_X1    g058(.A1(new_n474), .A2(KEYINPUT68), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n474), .A2(KEYINPUT68), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  AOI211_X1 g062(.A(new_n480), .B(new_n483), .C1(new_n487), .C2(G136), .ZN(G162));
  NAND2_X1  g063(.A1(new_n474), .A2(G138), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n474), .A2(new_n491), .A3(G138), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n494), .B1(new_n495), .B2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT69), .ZN(new_n497));
  OR2_X1    g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n497), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n498), .A2(new_n499), .B1(new_n478), .B2(G126), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n493), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  INV_X1    g077(.A(KEYINPUT6), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n503), .A2(G651), .ZN(new_n504));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT70), .B1(new_n505), .B2(KEYINPUT6), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT70), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(new_n503), .A3(G651), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n504), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n509), .A2(G50), .A3(G543), .ZN(new_n510));
  XNOR2_X1  g085(.A(new_n510), .B(KEYINPUT71), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n512), .B1(new_n513), .B2(KEYINPUT72), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT72), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n515), .A2(KEYINPUT5), .A3(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n517), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n509), .A2(new_n517), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  OAI22_X1  g095(.A1(new_n505), .A2(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n511), .A2(new_n521), .ZN(G166));
  NAND3_X1  g097(.A1(new_n509), .A2(G89), .A3(new_n517), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n517), .A2(G63), .A3(G651), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n523), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(new_n504), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n507), .B1(new_n503), .B2(G651), .ZN(new_n530));
  NOR3_X1   g105(.A1(new_n505), .A2(KEYINPUT70), .A3(KEYINPUT6), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(KEYINPUT73), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT73), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n509), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n533), .A2(G543), .A3(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(G51), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n528), .B1(new_n536), .B2(new_n537), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  NAND2_X1  g114(.A1(G77), .A2(G543), .ZN(new_n540));
  AND2_X1   g115(.A1(new_n514), .A2(new_n516), .ZN(new_n541));
  INV_X1    g116(.A(G64), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n505), .B1(new_n543), .B2(KEYINPUT74), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n544), .B1(KEYINPUT74), .B2(new_n543), .ZN(new_n545));
  NAND4_X1  g120(.A1(new_n533), .A2(G52), .A3(new_n535), .A4(G543), .ZN(new_n546));
  INV_X1    g121(.A(new_n519), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G90), .ZN(new_n548));
  AND3_X1   g123(.A1(new_n546), .A2(KEYINPUT75), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g124(.A(KEYINPUT75), .B1(new_n546), .B2(new_n548), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n545), .B1(new_n549), .B2(new_n550), .ZN(G301));
  INV_X1    g126(.A(G301), .ZN(G171));
  INV_X1    g127(.A(G56), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n553), .B1(new_n514), .B2(new_n516), .ZN(new_n554));
  AND2_X1   g129(.A1(G68), .A2(G543), .ZN(new_n555));
  OAI21_X1  g130(.A(G651), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  XNOR2_X1  g131(.A(KEYINPUT76), .B(G81), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n509), .A2(new_n517), .A3(new_n557), .ZN(new_n558));
  AND2_X1   g133(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(G43), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n536), .B2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  NAND4_X1  g138(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND4_X1  g141(.A1(G319), .A2(G483), .A3(G661), .A4(new_n566), .ZN(G188));
  AOI22_X1  g142(.A1(new_n517), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n568));
  OR2_X1    g143(.A1(new_n568), .A2(new_n505), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n547), .A2(G91), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  AND2_X1   g147(.A1(G53), .A2(G543), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n533), .A2(new_n535), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(KEYINPUT9), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT77), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT9), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n533), .A2(new_n577), .A3(new_n535), .A4(new_n573), .ZN(new_n578));
  AND3_X1   g153(.A1(new_n575), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n576), .B1(new_n575), .B2(new_n578), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n572), .B1(new_n579), .B2(new_n580), .ZN(G299));
  INV_X1    g156(.A(G166), .ZN(G303));
  AOI211_X1 g157(.A(KEYINPUT73), .B(new_n504), .C1(new_n506), .C2(new_n508), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n506), .A2(new_n508), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n534), .B1(new_n584), .B2(new_n529), .ZN(new_n585));
  NOR3_X1   g160(.A1(new_n583), .A2(new_n585), .A3(new_n512), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n586), .A2(KEYINPUT78), .A3(G49), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT78), .ZN(new_n588));
  INV_X1    g163(.A(G49), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n536), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  OR2_X1    g166(.A1(new_n517), .A2(G74), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n547), .A2(G87), .B1(new_n592), .B2(G651), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n591), .A2(new_n593), .ZN(G288));
  INV_X1    g169(.A(G61), .ZN(new_n595));
  OAI21_X1  g170(.A(KEYINPUT79), .B1(new_n541), .B2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(G73), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n597), .B2(new_n512), .ZN(new_n598));
  NOR3_X1   g173(.A1(new_n541), .A2(KEYINPUT79), .A3(new_n595), .ZN(new_n599));
  OAI21_X1  g174(.A(G651), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n509), .A2(G48), .A3(G543), .ZN(new_n601));
  AND2_X1   g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n547), .A2(G86), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(G305));
  NAND2_X1  g179(.A1(new_n586), .A2(G47), .ZN(new_n605));
  NAND2_X1  g180(.A1(G72), .A2(G543), .ZN(new_n606));
  INV_X1    g181(.A(G60), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n541), .B2(new_n607), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n547), .A2(G85), .B1(new_n608), .B2(G651), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n605), .A2(new_n609), .ZN(G290));
  NAND2_X1  g185(.A1(G301), .A2(G868), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n509), .A2(G92), .A3(new_n517), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(KEYINPUT10), .Z(new_n613));
  NAND2_X1  g188(.A1(new_n586), .A2(G54), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n517), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n615));
  OR2_X1    g190(.A1(new_n615), .A2(new_n505), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n613), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(KEYINPUT80), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT80), .ZN(new_n619));
  NAND4_X1  g194(.A1(new_n613), .A2(new_n619), .A3(new_n614), .A4(new_n616), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n611), .B1(new_n622), .B2(G868), .ZN(G284));
  OAI21_X1  g198(.A(new_n611), .B1(new_n622), .B2(G868), .ZN(G321));
  NAND2_X1  g199(.A1(G286), .A2(G868), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT81), .Z(new_n626));
  NOR2_X1   g201(.A1(new_n583), .A2(new_n585), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n577), .B1(new_n627), .B2(new_n573), .ZN(new_n628));
  INV_X1    g203(.A(new_n578), .ZN(new_n629));
  OAI21_X1  g204(.A(KEYINPUT77), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n575), .A2(new_n576), .A3(new_n578), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n571), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n626), .B1(G868), .B2(new_n632), .ZN(G297));
  OAI21_X1  g208(.A(new_n626), .B1(G868), .B2(new_n632), .ZN(G280));
  INV_X1    g209(.A(G559), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n622), .B1(new_n635), .B2(G860), .ZN(G148));
  INV_X1    g211(.A(KEYINPUT82), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(new_n621), .B2(G559), .ZN(new_n638));
  NAND4_X1  g213(.A1(new_n618), .A2(KEYINPUT82), .A3(new_n635), .A4(new_n620), .ZN(new_n639));
  AND3_X1   g214(.A1(new_n638), .A2(G868), .A3(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(G868), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n640), .B1(new_n641), .B2(new_n562), .ZN(G323));
  XNOR2_X1  g217(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g218(.A1(new_n478), .A2(G123), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT84), .ZN(new_n645));
  OR2_X1    g220(.A1(G99), .A2(G2105), .ZN(new_n646));
  OAI211_X1 g221(.A(new_n646), .B(G2104), .C1(G111), .C2(new_n470), .ZN(new_n647));
  INV_X1    g222(.A(G135), .ZN(new_n648));
  OAI211_X1 g223(.A(new_n645), .B(new_n647), .C1(new_n648), .C2(new_n486), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n649), .A2(G2096), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(G2096), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n466), .A2(new_n471), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT83), .B(KEYINPUT12), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n652), .B(new_n653), .Z(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT13), .B(G2100), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n650), .A2(new_n651), .A3(new_n656), .ZN(G156));
  XNOR2_X1  g232(.A(KEYINPUT15), .B(G2435), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT87), .B(G2438), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2427), .B(G2430), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n661), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n662), .A2(KEYINPUT14), .A3(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G1341), .B(G1348), .Z(new_n665));
  XNOR2_X1  g240(.A(G2443), .B(G2446), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n664), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT86), .ZN(new_n670));
  XOR2_X1   g245(.A(G2451), .B(G2454), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  OAI21_X1  g247(.A(G14), .B1(new_n668), .B2(new_n672), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n672), .B2(new_n668), .ZN(G401));
  XOR2_X1   g249(.A(KEYINPUT88), .B(KEYINPUT18), .Z(new_n675));
  XOR2_X1   g250(.A(G2084), .B(G2090), .Z(new_n676));
  XNOR2_X1  g251(.A(G2067), .B(G2678), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AND2_X1   g253(.A1(new_n678), .A2(KEYINPUT17), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n676), .A2(new_n677), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n675), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G2072), .B(G2078), .Z(new_n682));
  AOI21_X1  g257(.A(new_n682), .B1(new_n678), .B2(new_n675), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n681), .B(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G2096), .B(G2100), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(G227));
  XOR2_X1   g261(.A(G1971), .B(G1976), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT19), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1956), .B(G2474), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1961), .B(G1966), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n689), .A2(new_n690), .ZN(new_n692));
  NOR3_X1   g267(.A1(new_n688), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n688), .A2(new_n691), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT20), .Z(new_n695));
  AOI211_X1 g270(.A(new_n693), .B(new_n695), .C1(new_n688), .C2(new_n692), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT89), .ZN(new_n697));
  XOR2_X1   g272(.A(G1981), .B(G1986), .Z(new_n698));
  XNOR2_X1  g273(.A(G1991), .B(G1996), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n697), .B(new_n702), .ZN(G229));
  INV_X1    g278(.A(G16), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G6), .ZN(new_n705));
  INV_X1    g280(.A(G305), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n705), .B1(new_n706), .B2(new_n704), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT32), .B(G1981), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n709), .A2(KEYINPUT91), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n709), .A2(KEYINPUT91), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n704), .A2(G23), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n591), .A2(new_n593), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n713), .B1(new_n714), .B2(new_n704), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT33), .B(G1976), .Z(new_n716));
  OR2_X1    g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n715), .A2(new_n716), .ZN(new_n718));
  NOR2_X1   g293(.A1(G16), .A2(G22), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G166), .B2(G16), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT92), .B(G1971), .Z(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n717), .A2(new_n718), .A3(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(KEYINPUT34), .B1(new_n712), .B2(new_n723), .ZN(new_n724));
  OR4_X1    g299(.A1(KEYINPUT34), .A2(new_n710), .A3(new_n711), .A4(new_n723), .ZN(new_n725));
  INV_X1    g300(.A(G29), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G25), .ZN(new_n727));
  OAI21_X1  g302(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n728));
  INV_X1    g303(.A(G107), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(G2105), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n478), .B2(G119), .ZN(new_n731));
  INV_X1    g306(.A(G131), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n731), .B1(new_n486), .B2(new_n732), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n733), .A2(KEYINPUT90), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(KEYINPUT90), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n727), .B1(new_n736), .B2(new_n726), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT35), .B(G1991), .Z(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n737), .B(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(G290), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G16), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G16), .B2(G24), .ZN(new_n743));
  INV_X1    g318(.A(G1986), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n743), .A2(new_n744), .B1(KEYINPUT93), .B2(KEYINPUT36), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n744), .B2(new_n743), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n740), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n724), .A2(new_n725), .A3(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(KEYINPUT93), .A2(KEYINPUT36), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(G29), .A2(G35), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G162), .B2(G29), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT99), .B(KEYINPUT29), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(G2090), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n704), .A2(G21), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G168), .B2(new_n704), .ZN(new_n758));
  INV_X1    g333(.A(G1966), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(G1341), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n562), .A2(new_n704), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n704), .B2(G19), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n756), .B(new_n760), .C1(new_n761), .C2(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n755), .A2(G2090), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n765), .A2(KEYINPUT100), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(KEYINPUT100), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n764), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT31), .B(G11), .ZN(new_n769));
  XOR2_X1   g344(.A(KEYINPUT98), .B(G28), .Z(new_n770));
  NAND2_X1  g345(.A1(new_n770), .A2(KEYINPUT30), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n771), .A2(new_n726), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n770), .A2(KEYINPUT30), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n769), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT24), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n775), .A2(G34), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n726), .B1(new_n775), .B2(G34), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT97), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n778), .B2(new_n777), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G160), .B2(G29), .ZN(new_n781));
  OAI22_X1  g356(.A1(new_n649), .A2(new_n726), .B1(new_n781), .B2(G2084), .ZN(new_n782));
  AOI211_X1 g357(.A(new_n774), .B(new_n782), .C1(G2084), .C2(new_n781), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n763), .A2(new_n761), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n726), .A2(G32), .ZN(new_n785));
  AND3_X1   g360(.A1(new_n484), .A2(G141), .A3(new_n485), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n478), .A2(G129), .ZN(new_n787));
  NAND3_X1  g362(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT26), .Z(new_n789));
  NAND2_X1  g364(.A1(new_n472), .A2(G105), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n787), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n786), .A2(new_n791), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n785), .B1(new_n792), .B2(new_n726), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT27), .B(G1996), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n783), .A2(new_n784), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n726), .A2(G26), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT28), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n484), .A2(G140), .A3(new_n485), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT94), .ZN(new_n800));
  OAI21_X1  g375(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n801));
  INV_X1    g376(.A(G116), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n801), .B1(new_n802), .B2(G2105), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(new_n478), .B2(G128), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n799), .A2(new_n800), .A3(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n800), .B1(new_n799), .B2(new_n804), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n798), .B1(new_n808), .B2(new_n726), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT95), .B(G2067), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n726), .A2(G27), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G164), .B2(new_n726), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(G2078), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n726), .A2(G33), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT25), .Z(new_n817));
  INV_X1    g392(.A(G139), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(new_n486), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(G115), .A2(G2104), .ZN(new_n820));
  INV_X1    g395(.A(G127), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n820), .B1(new_n466), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n470), .B1(new_n822), .B2(KEYINPUT96), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(KEYINPUT96), .B2(new_n822), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n819), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n815), .B1(new_n826), .B2(new_n726), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(G2072), .ZN(new_n828));
  NOR4_X1   g403(.A1(new_n796), .A2(new_n811), .A3(new_n814), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n704), .A2(G5), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(G171), .B2(new_n704), .ZN(new_n831));
  INV_X1    g406(.A(G1961), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n768), .A2(new_n829), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n704), .A2(G4), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(new_n622), .B2(new_n704), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(G1348), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n704), .A2(G20), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT23), .Z(new_n839));
  AOI21_X1  g414(.A(new_n839), .B1(G299), .B2(G16), .ZN(new_n840));
  INV_X1    g415(.A(G1956), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NOR3_X1   g417(.A1(new_n834), .A2(new_n837), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(new_n748), .B2(new_n749), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n751), .A2(new_n844), .ZN(G311));
  OR2_X1    g420(.A1(new_n748), .A2(new_n749), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n846), .A2(new_n750), .A3(new_n843), .ZN(G150));
  NAND2_X1  g422(.A1(new_n622), .A2(G559), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT38), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n586), .A2(G43), .ZN(new_n850));
  INV_X1    g425(.A(G67), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n851), .B1(new_n514), .B2(new_n516), .ZN(new_n852));
  AND2_X1   g427(.A1(G80), .A2(G543), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI22_X1  g429(.A1(G93), .A2(new_n547), .B1(new_n854), .B2(G651), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n627), .A2(G55), .A3(G543), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n850), .A2(new_n855), .A3(new_n856), .A4(new_n559), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  AOI22_X1  g433(.A1(new_n850), .A2(new_n559), .B1(new_n855), .B2(new_n856), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n849), .B(new_n860), .ZN(new_n861));
  AND2_X1   g436(.A1(new_n861), .A2(KEYINPUT39), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n861), .A2(KEYINPUT39), .ZN(new_n863));
  NOR3_X1   g438(.A1(new_n862), .A2(new_n863), .A3(G860), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n855), .A2(new_n856), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(G860), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT37), .ZN(new_n867));
  OR2_X1    g442(.A1(new_n864), .A2(new_n867), .ZN(G145));
  NAND2_X1  g443(.A1(new_n487), .A2(G142), .ZN(new_n869));
  OAI21_X1  g444(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT101), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(G118), .ZN(new_n873));
  AOI22_X1  g448(.A1(new_n870), .A2(new_n871), .B1(new_n873), .B2(G2105), .ZN(new_n874));
  AOI22_X1  g449(.A1(new_n478), .A2(G130), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n869), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n736), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n876), .B1(new_n734), .B2(new_n735), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n877), .A2(new_n879), .A3(new_n654), .ZN(new_n880));
  INV_X1    g455(.A(new_n654), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n734), .A2(new_n735), .ZN(new_n882));
  INV_X1    g457(.A(new_n876), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n881), .B1(new_n884), .B2(new_n878), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n880), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n792), .ZN(new_n887));
  NOR3_X1   g462(.A1(new_n887), .A2(new_n806), .A3(new_n807), .ZN(new_n888));
  INV_X1    g463(.A(new_n807), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n792), .B1(new_n889), .B2(new_n805), .ZN(new_n890));
  OAI21_X1  g465(.A(G164), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n808), .A2(new_n792), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n887), .B1(new_n806), .B2(new_n807), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n892), .A2(new_n501), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n819), .A2(new_n825), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n891), .A2(new_n894), .A3(new_n826), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n886), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n898), .ZN(new_n900));
  INV_X1    g475(.A(new_n886), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT102), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n902), .B1(new_n900), .B2(new_n901), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n899), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(G162), .B(new_n476), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(new_n649), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(G37), .B1(new_n906), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n899), .A2(KEYINPUT103), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT103), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n886), .A2(new_n897), .A3(new_n912), .A4(new_n898), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n911), .A2(new_n913), .A3(new_n908), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT104), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n900), .A2(new_n901), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(KEYINPUT102), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(new_n903), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n914), .A2(new_n915), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n915), .B1(new_n914), .B2(new_n918), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n910), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(KEYINPUT40), .ZN(G395));
  AOI21_X1  g497(.A(KEYINPUT108), .B1(new_n865), .B2(new_n641), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n714), .A2(new_n741), .ZN(new_n924));
  NAND2_X1  g499(.A1(G288), .A2(G290), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT107), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n924), .A2(KEYINPUT107), .A3(new_n925), .ZN(new_n929));
  XNOR2_X1  g504(.A(G305), .B(G166), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(G305), .B(G303), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n932), .A2(KEYINPUT107), .A3(new_n925), .A4(new_n924), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n931), .A2(new_n933), .A3(KEYINPUT42), .ZN(new_n934));
  AOI21_X1  g509(.A(KEYINPUT42), .B1(new_n931), .B2(new_n933), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n638), .A2(new_n639), .A3(new_n860), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n860), .B1(new_n638), .B2(new_n639), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(G299), .A2(KEYINPUT105), .ZN(new_n940));
  INV_X1    g515(.A(new_n617), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n942), .B(new_n572), .C1(new_n579), .C2(new_n580), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n940), .A2(new_n941), .A3(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(G299), .A2(KEYINPUT105), .A3(new_n617), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OR2_X1    g521(.A1(new_n939), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n943), .A2(new_n941), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n630), .A2(new_n631), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n942), .B1(new_n949), .B2(new_n572), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n945), .ZN(new_n952));
  OAI21_X1  g527(.A(KEYINPUT41), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT41), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n944), .A2(new_n954), .A3(new_n945), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT106), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n944), .A2(new_n954), .A3(new_n945), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n957), .A2(KEYINPUT106), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n939), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n936), .A2(new_n947), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(G868), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n936), .B1(new_n959), .B2(new_n947), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n923), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n947), .A2(new_n959), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n964), .B1(new_n935), .B2(new_n934), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n965), .A2(KEYINPUT108), .A3(G868), .A4(new_n960), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT109), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n963), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n967), .B1(new_n963), .B2(new_n966), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n968), .A2(new_n969), .ZN(G295));
  AND2_X1   g545(.A1(new_n963), .A2(new_n966), .ZN(G331));
  INV_X1    g546(.A(KEYINPUT44), .ZN(new_n972));
  OAI221_X1 g547(.A(new_n545), .B1(G286), .B2(KEYINPUT110), .C1(new_n549), .C2(new_n550), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n865), .A2(new_n561), .ZN(new_n975));
  NAND2_X1  g550(.A1(G286), .A2(KEYINPUT110), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n975), .A2(new_n976), .A3(new_n857), .ZN(new_n977));
  OAI211_X1 g552(.A(KEYINPUT110), .B(G286), .C1(new_n858), .C2(new_n859), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n974), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  AND3_X1   g554(.A1(new_n975), .A2(new_n976), .A3(new_n857), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n976), .B1(new_n975), .B2(new_n857), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n973), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n979), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n983), .B1(new_n956), .B2(new_n958), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n931), .A2(new_n933), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n979), .A2(new_n944), .A3(new_n945), .A4(new_n982), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n987), .B(KEYINPUT111), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n984), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  AND3_X1   g564(.A1(new_n944), .A2(new_n954), .A3(new_n945), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n954), .B1(new_n944), .B2(new_n945), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n983), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n987), .ZN(new_n993));
  AOI21_X1  g568(.A(G37), .B1(new_n993), .B2(new_n985), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n989), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT112), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n989), .A2(new_n994), .A3(KEYINPUT112), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n997), .A2(KEYINPUT43), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n984), .A2(new_n988), .ZN(new_n1000));
  AOI21_X1  g575(.A(G37), .B1(new_n1000), .B2(new_n985), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT43), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1001), .A2(new_n1002), .A3(new_n989), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n972), .B1(new_n999), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1002), .B1(new_n1001), .B2(new_n989), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n989), .A2(new_n994), .A3(new_n1002), .ZN(new_n1006));
  NOR3_X1   g581(.A1(new_n1005), .A2(KEYINPUT44), .A3(new_n1006), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1004), .A2(new_n1007), .ZN(G397));
  INV_X1    g583(.A(G1971), .ZN(new_n1009));
  NAND2_X1  g584(.A1(G160), .A2(G40), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(G1384), .B1(new_n493), .B2(new_n500), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1011), .B1(new_n1012), .B2(KEYINPUT45), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(KEYINPUT45), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1009), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1012), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT50), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT50), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1012), .A2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g595(.A(KEYINPUT114), .B(G2090), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1018), .A2(new_n1011), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1016), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G8), .ZN(new_n1024));
  NOR2_X1   g599(.A1(G166), .A2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1025), .B1(KEYINPUT115), .B2(KEYINPUT55), .ZN(new_n1026));
  XOR2_X1   g601(.A(KEYINPUT115), .B(KEYINPUT55), .Z(new_n1027));
  OAI21_X1  g602(.A(new_n1026), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n1023), .A2(G8), .A3(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1028), .B1(new_n1023), .B2(G8), .ZN(new_n1030));
  XNOR2_X1  g605(.A(KEYINPUT116), .B(G8), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n759), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1032));
  INV_X1    g607(.A(G2084), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1018), .A2(new_n1033), .A3(new_n1011), .A4(new_n1020), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1031), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(G168), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT63), .ZN(new_n1037));
  NOR4_X1   g612(.A1(new_n1029), .A2(new_n1030), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1031), .ZN(new_n1040));
  INV_X1    g615(.A(G1976), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1039), .B(new_n1040), .C1(G288), .C2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n1044));
  OAI21_X1  g619(.A(KEYINPUT117), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT117), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1042), .A2(new_n1046), .A3(KEYINPUT52), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1044), .B1(new_n714), .B2(G1976), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT118), .ZN(new_n1049));
  OR2_X1    g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1042), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n1045), .A2(new_n1047), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  XOR2_X1   g627(.A(KEYINPUT119), .B(G86), .Z(new_n1053));
  NAND2_X1  g628(.A1(new_n547), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n600), .A2(new_n601), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(G1981), .ZN(new_n1056));
  INV_X1    g631(.A(G1981), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n600), .A2(new_n1057), .A3(new_n603), .A4(new_n601), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT49), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1056), .A2(KEYINPUT49), .A3(new_n1058), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1061), .A2(new_n1062), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT120), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT120), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1061), .A2(new_n1067), .A3(new_n1062), .A4(new_n1064), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  AND2_X1   g644(.A1(new_n1052), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1038), .A2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1028), .B1(new_n1023), .B2(new_n1040), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1029), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1036), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1073), .A2(new_n1052), .A3(new_n1069), .A4(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(new_n1037), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1071), .A2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1052), .A2(new_n1069), .A3(new_n1029), .ZN(new_n1078));
  NOR2_X1   g653(.A1(G288), .A2(G1976), .ZN(new_n1079));
  AOI22_X1  g654(.A1(new_n1069), .A2(new_n1079), .B1(new_n1057), .B2(new_n706), .ZN(new_n1080));
  OR2_X1    g655(.A1(new_n1080), .A2(new_n1063), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1077), .A2(KEYINPUT121), .A3(new_n1078), .A4(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT121), .ZN(new_n1083));
  AOI22_X1  g658(.A1(new_n1070), .A2(new_n1038), .B1(new_n1075), .B2(new_n1037), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1078), .B1(new_n1080), .B2(new_n1063), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1083), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT51), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1087), .B1(new_n1035), .B2(G286), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT123), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1089), .A2(new_n1090), .A3(G8), .ZN(new_n1091));
  NAND2_X1  g666(.A1(G286), .A2(new_n1040), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1090), .B1(new_n1089), .B2(G8), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1088), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1035), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1096), .A2(new_n1087), .A3(new_n1092), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT62), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1013), .ZN(new_n1099));
  INV_X1    g674(.A(G2078), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1099), .A2(KEYINPUT53), .A3(new_n1100), .A4(new_n1014), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1011), .B1(new_n1012), .B2(new_n1019), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1020), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NOR3_X1   g679(.A1(new_n1013), .A2(new_n1015), .A3(G2078), .ZN(new_n1105));
  OAI221_X1 g680(.A(new_n1101), .B1(new_n1104), .B2(G1961), .C1(new_n1105), .C2(KEYINPUT53), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(G171), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1098), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1095), .A2(KEYINPUT62), .A3(new_n1097), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1105), .A2(KEYINPUT53), .ZN(new_n1110));
  XNOR2_X1  g685(.A(G301), .B(KEYINPUT54), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1104), .A2(G1961), .ZN(new_n1112));
  NOR3_X1   g687(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1099), .A2(KEYINPUT124), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n1014), .A2(KEYINPUT53), .A3(new_n1100), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT124), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1013), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1114), .A2(new_n1115), .A3(new_n1117), .ZN(new_n1118));
  OR2_X1    g693(.A1(new_n1118), .A2(KEYINPUT125), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(KEYINPUT125), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1113), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1106), .A2(new_n1111), .ZN(new_n1122));
  AND4_X1   g697(.A1(new_n1095), .A2(new_n1121), .A3(new_n1097), .A4(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1104), .A2(G1348), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1039), .A2(G2067), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n941), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT122), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  OAI211_X1 g703(.A(KEYINPUT122), .B(new_n941), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1129));
  NAND2_X1  g704(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT57), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n572), .B(new_n1131), .C1(new_n628), .C2(new_n629), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1018), .A2(new_n1011), .A3(new_n1020), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(new_n841), .ZN(new_n1135));
  XNOR2_X1  g710(.A(KEYINPUT56), .B(G2072), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1099), .A2(new_n1014), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  AOI22_X1  g713(.A1(new_n1128), .A2(new_n1129), .B1(new_n1133), .B2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1138), .A2(new_n1133), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n617), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1141));
  OAI221_X1 g716(.A(new_n941), .B1(G2067), .B2(new_n1039), .C1(new_n1104), .C2(G1348), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1141), .A2(KEYINPUT60), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1133), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT61), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1144), .A2(new_n1145), .A3(new_n1135), .A4(new_n1137), .ZN(new_n1146));
  OAI21_X1  g721(.A(KEYINPUT61), .B1(new_n1138), .B2(new_n1133), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1143), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT59), .ZN(new_n1149));
  INV_X1    g724(.A(G1996), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1099), .A2(new_n1150), .A3(new_n1014), .ZN(new_n1151));
  XOR2_X1   g726(.A(KEYINPUT58), .B(G1341), .Z(new_n1152));
  NAND2_X1  g727(.A1(new_n1039), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1149), .B1(new_n1154), .B2(new_n562), .ZN(new_n1155));
  AOI211_X1 g730(.A(KEYINPUT59), .B(new_n561), .C1(new_n1151), .C2(new_n1153), .ZN(new_n1156));
  OAI22_X1  g731(.A1(new_n1155), .A2(new_n1156), .B1(KEYINPUT60), .B2(new_n1142), .ZN(new_n1157));
  OAI22_X1  g732(.A1(new_n1139), .A2(new_n1140), .B1(new_n1148), .B2(new_n1157), .ZN(new_n1158));
  AOI22_X1  g733(.A1(new_n1108), .A2(new_n1109), .B1(new_n1123), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1070), .A2(new_n1073), .ZN(new_n1160));
  OAI211_X1 g735(.A(new_n1082), .B(new_n1086), .C1(new_n1159), .C2(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n808), .B(G2067), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n792), .B(G1996), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n736), .A2(new_n738), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n882), .A2(new_n739), .ZN(new_n1165));
  AND4_X1   g740(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .A4(new_n1165), .ZN(new_n1166));
  NOR2_X1   g741(.A1(G290), .A2(G1986), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1167), .B(KEYINPUT113), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1168), .B1(G1986), .B2(G290), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1166), .A2(new_n1169), .ZN(new_n1170));
  NOR3_X1   g745(.A1(new_n1012), .A2(new_n1010), .A3(KEYINPUT45), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1161), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1168), .A2(KEYINPUT48), .A3(new_n1171), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1171), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1174), .B1(new_n1166), .B2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(KEYINPUT48), .B1(new_n1168), .B2(new_n1171), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1175), .B1(new_n1162), .B2(new_n792), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT46), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1171), .A2(new_n1150), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1179), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1181), .A2(new_n1180), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1183), .B(KEYINPUT127), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1185));
  XOR2_X1   g760(.A(new_n1185), .B(KEYINPUT47), .Z(new_n1186));
  XNOR2_X1  g761(.A(new_n1164), .B(KEYINPUT126), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1188));
  INV_X1    g763(.A(new_n808), .ZN(new_n1189));
  OAI22_X1  g764(.A1(new_n1187), .A2(new_n1188), .B1(G2067), .B2(new_n1189), .ZN(new_n1190));
  AOI211_X1 g765(.A(new_n1178), .B(new_n1186), .C1(new_n1171), .C2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1173), .A2(new_n1191), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g767(.A1(G229), .A2(new_n461), .A3(G401), .A4(G227), .ZN(new_n1194));
  OAI211_X1 g768(.A(new_n921), .B(new_n1194), .C1(new_n1005), .C2(new_n1006), .ZN(G225));
  INV_X1    g769(.A(G225), .ZN(G308));
endmodule


