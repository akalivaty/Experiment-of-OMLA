

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U561 ( .A1(n534), .A2(G2105), .ZN(n883) );
  XOR2_X1 U562 ( .A(KEYINPUT64), .B(G2104), .Z(n534) );
  XOR2_X1 U563 ( .A(n645), .B(KEYINPUT27), .Z(n527) );
  AND2_X1 U564 ( .A1(n987), .A2(n762), .ZN(n528) );
  NOR2_X1 U565 ( .A1(G299), .A2(n650), .ZN(n647) );
  AND2_X1 U566 ( .A1(n672), .A2(n678), .ZN(n673) );
  INV_X1 U567 ( .A(KEYINPUT14), .ZN(n623) );
  XNOR2_X1 U568 ( .A(n624), .B(n623), .ZN(n625) );
  OR2_X1 U569 ( .A1(n749), .A2(n528), .ZN(n750) );
  XOR2_X1 U570 ( .A(KEYINPUT1), .B(n541), .Z(n789) );
  XNOR2_X1 U571 ( .A(n535), .B(KEYINPUT65), .ZN(n888) );
  OR2_X1 U572 ( .A1(n751), .A2(n750), .ZN(n765) );
  NOR2_X1 U573 ( .A1(G543), .A2(G651), .ZN(n793) );
  XOR2_X1 U574 ( .A(KEYINPUT75), .B(n635), .Z(n977) );
  NOR2_X1 U575 ( .A1(n558), .A2(n557), .ZN(G160) );
  AND2_X1 U576 ( .A1(G2104), .A2(G2105), .ZN(n887) );
  NAND2_X1 U577 ( .A1(G114), .A2(n887), .ZN(n529) );
  XNOR2_X1 U578 ( .A(n529), .B(KEYINPUT85), .ZN(n539) );
  NAND2_X1 U579 ( .A1(n883), .A2(G102), .ZN(n532) );
  NOR2_X1 U580 ( .A1(G2104), .A2(G2105), .ZN(n530) );
  XOR2_X2 U581 ( .A(KEYINPUT17), .B(n530), .Z(n882) );
  NAND2_X1 U582 ( .A1(n882), .A2(G138), .ZN(n531) );
  AND2_X1 U583 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U584 ( .A(KEYINPUT86), .B(n533), .ZN(n537) );
  NAND2_X1 U585 ( .A1(G2105), .A2(n534), .ZN(n535) );
  NAND2_X1 U586 ( .A1(n888), .A2(G126), .ZN(n536) );
  NAND2_X1 U587 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U588 ( .A1(n539), .A2(n538), .ZN(G164) );
  NAND2_X1 U589 ( .A1(G91), .A2(n793), .ZN(n540) );
  XNOR2_X1 U590 ( .A(n540), .B(KEYINPUT70), .ZN(n549) );
  INV_X1 U591 ( .A(G651), .ZN(n542) );
  NOR2_X1 U592 ( .A1(G543), .A2(n542), .ZN(n541) );
  NAND2_X1 U593 ( .A1(G65), .A2(n789), .ZN(n544) );
  XOR2_X1 U594 ( .A(KEYINPUT0), .B(G543), .Z(n597) );
  NOR2_X1 U595 ( .A1(n597), .A2(n542), .ZN(n794) );
  NAND2_X1 U596 ( .A1(G78), .A2(n794), .ZN(n543) );
  NAND2_X1 U597 ( .A1(n544), .A2(n543), .ZN(n547) );
  NOR2_X1 U598 ( .A1(n597), .A2(G651), .ZN(n790) );
  NAND2_X1 U599 ( .A1(G53), .A2(n790), .ZN(n545) );
  XNOR2_X1 U600 ( .A(KEYINPUT71), .B(n545), .ZN(n546) );
  NOR2_X1 U601 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U602 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U603 ( .A(KEYINPUT72), .B(n550), .ZN(G299) );
  NAND2_X1 U604 ( .A1(G101), .A2(n883), .ZN(n551) );
  XOR2_X1 U605 ( .A(KEYINPUT23), .B(n551), .Z(n552) );
  XNOR2_X1 U606 ( .A(n552), .B(KEYINPUT66), .ZN(n554) );
  NAND2_X1 U607 ( .A1(G137), .A2(n882), .ZN(n553) );
  NAND2_X1 U608 ( .A1(n554), .A2(n553), .ZN(n558) );
  NAND2_X1 U609 ( .A1(G113), .A2(n887), .ZN(n556) );
  NAND2_X1 U610 ( .A1(G125), .A2(n888), .ZN(n555) );
  NAND2_X1 U611 ( .A1(n556), .A2(n555), .ZN(n557) );
  NAND2_X1 U612 ( .A1(G61), .A2(n789), .ZN(n560) );
  NAND2_X1 U613 ( .A1(G48), .A2(n790), .ZN(n559) );
  NAND2_X1 U614 ( .A1(n560), .A2(n559), .ZN(n563) );
  NAND2_X1 U615 ( .A1(n794), .A2(G73), .ZN(n561) );
  XOR2_X1 U616 ( .A(KEYINPUT2), .B(n561), .Z(n562) );
  NOR2_X1 U617 ( .A1(n563), .A2(n562), .ZN(n565) );
  NAND2_X1 U618 ( .A1(n793), .A2(G86), .ZN(n564) );
  NAND2_X1 U619 ( .A1(n565), .A2(n564), .ZN(G305) );
  NAND2_X1 U620 ( .A1(G64), .A2(n789), .ZN(n567) );
  NAND2_X1 U621 ( .A1(G52), .A2(n790), .ZN(n566) );
  NAND2_X1 U622 ( .A1(n567), .A2(n566), .ZN(n574) );
  XNOR2_X1 U623 ( .A(KEYINPUT68), .B(KEYINPUT9), .ZN(n572) );
  NAND2_X1 U624 ( .A1(n794), .A2(G77), .ZN(n570) );
  NAND2_X1 U625 ( .A1(n793), .A2(G90), .ZN(n568) );
  XOR2_X1 U626 ( .A(KEYINPUT67), .B(n568), .Z(n569) );
  NAND2_X1 U627 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U628 ( .A(n572), .B(n571), .Z(n573) );
  NOR2_X1 U629 ( .A1(n574), .A2(n573), .ZN(G171) );
  NAND2_X1 U630 ( .A1(G89), .A2(n793), .ZN(n575) );
  XNOR2_X1 U631 ( .A(n575), .B(KEYINPUT78), .ZN(n576) );
  XNOR2_X1 U632 ( .A(n576), .B(KEYINPUT4), .ZN(n578) );
  NAND2_X1 U633 ( .A1(G76), .A2(n794), .ZN(n577) );
  NAND2_X1 U634 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U635 ( .A(n579), .B(KEYINPUT5), .ZN(n584) );
  NAND2_X1 U636 ( .A1(G63), .A2(n789), .ZN(n581) );
  NAND2_X1 U637 ( .A1(G51), .A2(n790), .ZN(n580) );
  NAND2_X1 U638 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U639 ( .A(KEYINPUT6), .B(n582), .Z(n583) );
  NAND2_X1 U640 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U641 ( .A(n585), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U642 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U643 ( .A1(G88), .A2(n793), .ZN(n587) );
  NAND2_X1 U644 ( .A1(G75), .A2(n794), .ZN(n586) );
  NAND2_X1 U645 ( .A1(n587), .A2(n586), .ZN(n591) );
  NAND2_X1 U646 ( .A1(G62), .A2(n789), .ZN(n589) );
  NAND2_X1 U647 ( .A1(G50), .A2(n790), .ZN(n588) );
  NAND2_X1 U648 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U649 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U650 ( .A(n592), .B(KEYINPUT81), .ZN(G303) );
  INV_X1 U651 ( .A(G303), .ZN(G166) );
  NAND2_X1 U652 ( .A1(G49), .A2(n790), .ZN(n594) );
  NAND2_X1 U653 ( .A1(G74), .A2(G651), .ZN(n593) );
  NAND2_X1 U654 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U655 ( .A1(n789), .A2(n595), .ZN(n596) );
  XNOR2_X1 U656 ( .A(n596), .B(KEYINPUT80), .ZN(n599) );
  NAND2_X1 U657 ( .A1(G87), .A2(n597), .ZN(n598) );
  NAND2_X1 U658 ( .A1(n599), .A2(n598), .ZN(G288) );
  NAND2_X1 U659 ( .A1(G60), .A2(n789), .ZN(n601) );
  NAND2_X1 U660 ( .A1(G47), .A2(n790), .ZN(n600) );
  NAND2_X1 U661 ( .A1(n601), .A2(n600), .ZN(n605) );
  NAND2_X1 U662 ( .A1(G85), .A2(n793), .ZN(n603) );
  NAND2_X1 U663 ( .A1(G72), .A2(n794), .ZN(n602) );
  NAND2_X1 U664 ( .A1(n603), .A2(n602), .ZN(n604) );
  OR2_X1 U665 ( .A1(n605), .A2(n604), .ZN(G290) );
  NOR2_X1 U666 ( .A1(G164), .A2(G1384), .ZN(n718) );
  NAND2_X1 U667 ( .A1(G160), .A2(G40), .ZN(n717) );
  INV_X1 U668 ( .A(n717), .ZN(n606) );
  NAND2_X2 U669 ( .A1(n718), .A2(n606), .ZN(n679) );
  NAND2_X1 U670 ( .A1(G8), .A2(n679), .ZN(n711) );
  XNOR2_X1 U671 ( .A(KEYINPUT24), .B(KEYINPUT92), .ZN(n607) );
  XNOR2_X1 U672 ( .A(n607), .B(KEYINPUT91), .ZN(n609) );
  NOR2_X1 U673 ( .A1(G1981), .A2(G305), .ZN(n608) );
  XNOR2_X1 U674 ( .A(n609), .B(n608), .ZN(n610) );
  NOR2_X1 U675 ( .A1(n711), .A2(n610), .ZN(n716) );
  NOR2_X1 U676 ( .A1(G1966), .A2(n711), .ZN(n662) );
  INV_X1 U677 ( .A(n662), .ZN(n672) );
  NAND2_X1 U678 ( .A1(G54), .A2(n790), .ZN(n612) );
  NAND2_X1 U679 ( .A1(G79), .A2(n794), .ZN(n611) );
  NAND2_X1 U680 ( .A1(n612), .A2(n611), .ZN(n617) );
  NAND2_X1 U681 ( .A1(G66), .A2(n789), .ZN(n614) );
  NAND2_X1 U682 ( .A1(G92), .A2(n793), .ZN(n613) );
  NAND2_X1 U683 ( .A1(n614), .A2(n613), .ZN(n615) );
  XOR2_X1 U684 ( .A(KEYINPUT77), .B(n615), .Z(n616) );
  NOR2_X1 U685 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U686 ( .A(KEYINPUT15), .B(n618), .ZN(n973) );
  INV_X1 U687 ( .A(n679), .ZN(n656) );
  NAND2_X1 U688 ( .A1(G2067), .A2(n656), .ZN(n619) );
  XNOR2_X1 U689 ( .A(n619), .B(KEYINPUT98), .ZN(n621) );
  NAND2_X1 U690 ( .A1(G1348), .A2(n679), .ZN(n620) );
  NAND2_X1 U691 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U692 ( .A1(n973), .A2(n622), .ZN(n644) );
  NAND2_X1 U693 ( .A1(n622), .A2(n973), .ZN(n642) );
  NAND2_X1 U694 ( .A1(G56), .A2(n789), .ZN(n624) );
  XNOR2_X1 U695 ( .A(n625), .B(KEYINPUT73), .ZN(n627) );
  NAND2_X1 U696 ( .A1(G43), .A2(n790), .ZN(n626) );
  NAND2_X1 U697 ( .A1(n627), .A2(n626), .ZN(n634) );
  NAND2_X1 U698 ( .A1(n793), .A2(G81), .ZN(n628) );
  XNOR2_X1 U699 ( .A(n628), .B(KEYINPUT12), .ZN(n630) );
  NAND2_X1 U700 ( .A1(G68), .A2(n794), .ZN(n629) );
  NAND2_X1 U701 ( .A1(n630), .A2(n629), .ZN(n631) );
  XOR2_X1 U702 ( .A(KEYINPUT74), .B(n631), .Z(n632) );
  XNOR2_X1 U703 ( .A(KEYINPUT13), .B(n632), .ZN(n633) );
  NOR2_X1 U704 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U705 ( .A(G1996), .B(KEYINPUT96), .Z(n953) );
  NOR2_X1 U706 ( .A1(n679), .A2(n953), .ZN(n636) );
  XOR2_X1 U707 ( .A(KEYINPUT26), .B(n636), .Z(n637) );
  NAND2_X1 U708 ( .A1(n977), .A2(n637), .ZN(n640) );
  NAND2_X1 U709 ( .A1(G1341), .A2(n679), .ZN(n638) );
  XNOR2_X1 U710 ( .A(KEYINPUT97), .B(n638), .ZN(n639) );
  NOR2_X1 U711 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U712 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U713 ( .A1(n644), .A2(n643), .ZN(n649) );
  NAND2_X1 U714 ( .A1(n656), .A2(G2072), .ZN(n645) );
  NAND2_X1 U715 ( .A1(G1956), .A2(n679), .ZN(n646) );
  NAND2_X1 U716 ( .A1(n527), .A2(n646), .ZN(n650) );
  XNOR2_X1 U717 ( .A(n647), .B(KEYINPUT99), .ZN(n648) );
  AND2_X1 U718 ( .A1(n649), .A2(n648), .ZN(n654) );
  XOR2_X1 U719 ( .A(KEYINPUT95), .B(KEYINPUT28), .Z(n652) );
  NAND2_X1 U720 ( .A1(G299), .A2(n650), .ZN(n651) );
  XOR2_X1 U721 ( .A(n652), .B(n651), .Z(n653) );
  NOR2_X1 U722 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U723 ( .A(n655), .B(KEYINPUT29), .ZN(n661) );
  XNOR2_X1 U724 ( .A(G2078), .B(KEYINPUT25), .ZN(n954) );
  NAND2_X1 U725 ( .A1(n656), .A2(n954), .ZN(n657) );
  XNOR2_X1 U726 ( .A(n657), .B(KEYINPUT94), .ZN(n659) );
  INV_X1 U727 ( .A(G1961), .ZN(n1001) );
  NAND2_X1 U728 ( .A1(n1001), .A2(n679), .ZN(n658) );
  NAND2_X1 U729 ( .A1(n659), .A2(n658), .ZN(n666) );
  NAND2_X1 U730 ( .A1(G171), .A2(n666), .ZN(n660) );
  NAND2_X1 U731 ( .A1(n661), .A2(n660), .ZN(n671) );
  NOR2_X1 U732 ( .A1(G2084), .A2(n679), .ZN(n674) );
  NOR2_X1 U733 ( .A1(n662), .A2(n674), .ZN(n663) );
  NAND2_X1 U734 ( .A1(G8), .A2(n663), .ZN(n664) );
  XNOR2_X1 U735 ( .A(KEYINPUT30), .B(n664), .ZN(n665) );
  NOR2_X1 U736 ( .A1(G168), .A2(n665), .ZN(n668) );
  NOR2_X1 U737 ( .A1(G171), .A2(n666), .ZN(n667) );
  NOR2_X1 U738 ( .A1(n668), .A2(n667), .ZN(n669) );
  XOR2_X1 U739 ( .A(KEYINPUT31), .B(n669), .Z(n670) );
  NAND2_X1 U740 ( .A1(n671), .A2(n670), .ZN(n678) );
  XNOR2_X1 U741 ( .A(n673), .B(KEYINPUT100), .ZN(n677) );
  NAND2_X1 U742 ( .A1(G8), .A2(n674), .ZN(n675) );
  XOR2_X1 U743 ( .A(KEYINPUT93), .B(n675), .Z(n676) );
  NAND2_X1 U744 ( .A1(n677), .A2(n676), .ZN(n691) );
  XOR2_X1 U745 ( .A(KEYINPUT103), .B(KEYINPUT32), .Z(n689) );
  NAND2_X1 U746 ( .A1(n678), .A2(G286), .ZN(n686) );
  NOR2_X1 U747 ( .A1(G2090), .A2(n679), .ZN(n680) );
  XNOR2_X1 U748 ( .A(KEYINPUT101), .B(n680), .ZN(n683) );
  NOR2_X1 U749 ( .A1(G1971), .A2(n711), .ZN(n681) );
  NOR2_X1 U750 ( .A1(G166), .A2(n681), .ZN(n682) );
  NAND2_X1 U751 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U752 ( .A(n684), .B(KEYINPUT102), .ZN(n685) );
  NAND2_X1 U753 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U754 ( .A1(n687), .A2(G8), .ZN(n688) );
  XNOR2_X1 U755 ( .A(n689), .B(n688), .ZN(n690) );
  NAND2_X1 U756 ( .A1(n691), .A2(n690), .ZN(n710) );
  NOR2_X1 U757 ( .A1(G1971), .A2(G303), .ZN(n692) );
  XNOR2_X1 U758 ( .A(KEYINPUT104), .B(n692), .ZN(n693) );
  NOR2_X1 U759 ( .A1(KEYINPUT33), .A2(n693), .ZN(n694) );
  NAND2_X1 U760 ( .A1(n710), .A2(n694), .ZN(n697) );
  INV_X1 U761 ( .A(n711), .ZN(n695) );
  NAND2_X1 U762 ( .A1(n695), .A2(KEYINPUT105), .ZN(n696) );
  NAND2_X1 U763 ( .A1(n697), .A2(n696), .ZN(n698) );
  OR2_X1 U764 ( .A1(G1976), .A2(G288), .ZN(n981) );
  NAND2_X1 U765 ( .A1(n698), .A2(n981), .ZN(n707) );
  XNOR2_X1 U766 ( .A(G1981), .B(G305), .ZN(n992) );
  NAND2_X1 U767 ( .A1(G1976), .A2(G288), .ZN(n980) );
  NOR2_X1 U768 ( .A1(KEYINPUT105), .A2(n711), .ZN(n701) );
  NAND2_X1 U769 ( .A1(n980), .A2(n701), .ZN(n699) );
  INV_X1 U770 ( .A(KEYINPUT33), .ZN(n700) );
  NAND2_X1 U771 ( .A1(n699), .A2(n700), .ZN(n704) );
  NOR2_X1 U772 ( .A1(n981), .A2(n700), .ZN(n702) );
  NAND2_X1 U773 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U774 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U775 ( .A1(n992), .A2(n705), .ZN(n706) );
  NAND2_X1 U776 ( .A1(n707), .A2(n706), .ZN(n714) );
  NOR2_X1 U777 ( .A1(G2090), .A2(G303), .ZN(n708) );
  NAND2_X1 U778 ( .A1(G8), .A2(n708), .ZN(n709) );
  NAND2_X1 U779 ( .A1(n710), .A2(n709), .ZN(n712) );
  NAND2_X1 U780 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U781 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U782 ( .A1(n716), .A2(n715), .ZN(n751) );
  NOR2_X1 U783 ( .A1(n718), .A2(n717), .ZN(n762) );
  NAND2_X1 U784 ( .A1(G140), .A2(n882), .ZN(n720) );
  NAND2_X1 U785 ( .A1(G104), .A2(n883), .ZN(n719) );
  NAND2_X1 U786 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U787 ( .A(KEYINPUT34), .B(n721), .ZN(n726) );
  NAND2_X1 U788 ( .A1(G116), .A2(n887), .ZN(n723) );
  NAND2_X1 U789 ( .A1(G128), .A2(n888), .ZN(n722) );
  NAND2_X1 U790 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U791 ( .A(n724), .B(KEYINPUT35), .Z(n725) );
  NOR2_X1 U792 ( .A1(n726), .A2(n725), .ZN(n727) );
  XOR2_X1 U793 ( .A(KEYINPUT36), .B(n727), .Z(n728) );
  XNOR2_X1 U794 ( .A(KEYINPUT87), .B(n728), .ZN(n897) );
  XNOR2_X1 U795 ( .A(G2067), .B(KEYINPUT37), .ZN(n760) );
  NOR2_X1 U796 ( .A1(n897), .A2(n760), .ZN(n931) );
  NAND2_X1 U797 ( .A1(n762), .A2(n931), .ZN(n758) );
  NAND2_X1 U798 ( .A1(G131), .A2(n882), .ZN(n730) );
  NAND2_X1 U799 ( .A1(G95), .A2(n883), .ZN(n729) );
  NAND2_X1 U800 ( .A1(n730), .A2(n729), .ZN(n734) );
  NAND2_X1 U801 ( .A1(G107), .A2(n887), .ZN(n732) );
  NAND2_X1 U802 ( .A1(G119), .A2(n888), .ZN(n731) );
  NAND2_X1 U803 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U804 ( .A1(n734), .A2(n733), .ZN(n867) );
  INV_X1 U805 ( .A(G1991), .ZN(n949) );
  NOR2_X1 U806 ( .A1(n867), .A2(n949), .ZN(n746) );
  NAND2_X1 U807 ( .A1(G105), .A2(n883), .ZN(n735) );
  XOR2_X1 U808 ( .A(KEYINPUT38), .B(n735), .Z(n741) );
  NAND2_X1 U809 ( .A1(n887), .A2(G117), .ZN(n736) );
  XNOR2_X1 U810 ( .A(n736), .B(KEYINPUT88), .ZN(n738) );
  NAND2_X1 U811 ( .A1(G129), .A2(n888), .ZN(n737) );
  NAND2_X1 U812 ( .A1(n738), .A2(n737), .ZN(n739) );
  XOR2_X1 U813 ( .A(KEYINPUT89), .B(n739), .Z(n740) );
  NOR2_X1 U814 ( .A1(n741), .A2(n740), .ZN(n743) );
  NAND2_X1 U815 ( .A1(n882), .A2(G141), .ZN(n742) );
  NAND2_X1 U816 ( .A1(n743), .A2(n742), .ZN(n894) );
  NAND2_X1 U817 ( .A1(G1996), .A2(n894), .ZN(n744) );
  XOR2_X1 U818 ( .A(KEYINPUT90), .B(n744), .Z(n745) );
  NOR2_X1 U819 ( .A1(n746), .A2(n745), .ZN(n939) );
  INV_X1 U820 ( .A(n762), .ZN(n747) );
  NOR2_X1 U821 ( .A1(n939), .A2(n747), .ZN(n755) );
  INV_X1 U822 ( .A(n755), .ZN(n748) );
  NAND2_X1 U823 ( .A1(n758), .A2(n748), .ZN(n749) );
  XNOR2_X1 U824 ( .A(G1986), .B(G290), .ZN(n987) );
  NOR2_X1 U825 ( .A1(n894), .A2(G1996), .ZN(n752) );
  XNOR2_X1 U826 ( .A(n752), .B(KEYINPUT106), .ZN(n922) );
  NOR2_X1 U827 ( .A1(G1986), .A2(G290), .ZN(n753) );
  AND2_X1 U828 ( .A1(n949), .A2(n867), .ZN(n927) );
  NOR2_X1 U829 ( .A1(n753), .A2(n927), .ZN(n754) );
  NOR2_X1 U830 ( .A1(n755), .A2(n754), .ZN(n756) );
  NOR2_X1 U831 ( .A1(n922), .A2(n756), .ZN(n757) );
  XNOR2_X1 U832 ( .A(n757), .B(KEYINPUT39), .ZN(n759) );
  NAND2_X1 U833 ( .A1(n759), .A2(n758), .ZN(n761) );
  NAND2_X1 U834 ( .A1(n897), .A2(n760), .ZN(n932) );
  NAND2_X1 U835 ( .A1(n761), .A2(n932), .ZN(n763) );
  NAND2_X1 U836 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U837 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U838 ( .A(n766), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U839 ( .A(G57), .ZN(G237) );
  INV_X1 U840 ( .A(G132), .ZN(G219) );
  INV_X1 U841 ( .A(G82), .ZN(G220) );
  NAND2_X1 U842 ( .A1(G94), .A2(G452), .ZN(n767) );
  XNOR2_X1 U843 ( .A(n767), .B(KEYINPUT69), .ZN(G173) );
  NAND2_X1 U844 ( .A1(G7), .A2(G661), .ZN(n768) );
  XNOR2_X1 U845 ( .A(n768), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U846 ( .A(G223), .ZN(n830) );
  NAND2_X1 U847 ( .A1(n830), .A2(G567), .ZN(n769) );
  XOR2_X1 U848 ( .A(KEYINPUT11), .B(n769), .Z(G234) );
  NAND2_X1 U849 ( .A1(n977), .A2(G860), .ZN(G153) );
  XOR2_X1 U850 ( .A(G171), .B(KEYINPUT76), .Z(G301) );
  NAND2_X1 U851 ( .A1(G868), .A2(G301), .ZN(n771) );
  INV_X1 U852 ( .A(G868), .ZN(n812) );
  NAND2_X1 U853 ( .A1(n973), .A2(n812), .ZN(n770) );
  NAND2_X1 U854 ( .A1(n771), .A2(n770), .ZN(G284) );
  NOR2_X1 U855 ( .A1(G286), .A2(n812), .ZN(n773) );
  NOR2_X1 U856 ( .A1(G299), .A2(G868), .ZN(n772) );
  NOR2_X1 U857 ( .A1(n773), .A2(n772), .ZN(G297) );
  INV_X1 U858 ( .A(G559), .ZN(n776) );
  NOR2_X1 U859 ( .A1(G860), .A2(n776), .ZN(n774) );
  NOR2_X1 U860 ( .A1(n973), .A2(n774), .ZN(n775) );
  XOR2_X1 U861 ( .A(KEYINPUT16), .B(n775), .Z(G148) );
  INV_X1 U862 ( .A(n973), .ZN(n799) );
  NAND2_X1 U863 ( .A1(n776), .A2(n799), .ZN(n777) );
  NAND2_X1 U864 ( .A1(n777), .A2(G868), .ZN(n779) );
  OR2_X1 U865 ( .A1(n977), .A2(G868), .ZN(n778) );
  NAND2_X1 U866 ( .A1(n779), .A2(n778), .ZN(G282) );
  NAND2_X1 U867 ( .A1(G135), .A2(n882), .ZN(n781) );
  NAND2_X1 U868 ( .A1(G111), .A2(n887), .ZN(n780) );
  NAND2_X1 U869 ( .A1(n781), .A2(n780), .ZN(n786) );
  NAND2_X1 U870 ( .A1(G123), .A2(n888), .ZN(n782) );
  XNOR2_X1 U871 ( .A(n782), .B(KEYINPUT18), .ZN(n784) );
  NAND2_X1 U872 ( .A1(n883), .A2(G99), .ZN(n783) );
  NAND2_X1 U873 ( .A1(n784), .A2(n783), .ZN(n785) );
  NOR2_X1 U874 ( .A1(n786), .A2(n785), .ZN(n926) );
  XNOR2_X1 U875 ( .A(G2096), .B(n926), .ZN(n788) );
  INV_X1 U876 ( .A(G2100), .ZN(n787) );
  NAND2_X1 U877 ( .A1(n788), .A2(n787), .ZN(G156) );
  NAND2_X1 U878 ( .A1(G67), .A2(n789), .ZN(n792) );
  NAND2_X1 U879 ( .A1(G55), .A2(n790), .ZN(n791) );
  NAND2_X1 U880 ( .A1(n792), .A2(n791), .ZN(n798) );
  NAND2_X1 U881 ( .A1(G93), .A2(n793), .ZN(n796) );
  NAND2_X1 U882 ( .A1(G80), .A2(n794), .ZN(n795) );
  NAND2_X1 U883 ( .A1(n796), .A2(n795), .ZN(n797) );
  OR2_X1 U884 ( .A1(n798), .A2(n797), .ZN(n813) );
  NAND2_X1 U885 ( .A1(n799), .A2(G559), .ZN(n810) );
  XOR2_X1 U886 ( .A(n810), .B(n977), .Z(n800) );
  NOR2_X1 U887 ( .A1(G860), .A2(n800), .ZN(n801) );
  XOR2_X1 U888 ( .A(KEYINPUT79), .B(n801), .Z(n802) );
  XOR2_X1 U889 ( .A(n813), .B(n802), .Z(G145) );
  XNOR2_X1 U890 ( .A(KEYINPUT82), .B(KEYINPUT19), .ZN(n804) );
  XNOR2_X1 U891 ( .A(G290), .B(G166), .ZN(n803) );
  XNOR2_X1 U892 ( .A(n804), .B(n803), .ZN(n807) );
  XOR2_X1 U893 ( .A(n977), .B(G299), .Z(n805) );
  XNOR2_X1 U894 ( .A(G288), .B(n805), .ZN(n806) );
  XNOR2_X1 U895 ( .A(n807), .B(n806), .ZN(n809) );
  XOR2_X1 U896 ( .A(G305), .B(n813), .Z(n808) );
  XNOR2_X1 U897 ( .A(n809), .B(n808), .ZN(n900) );
  XOR2_X1 U898 ( .A(n900), .B(n810), .Z(n811) );
  NAND2_X1 U899 ( .A1(G868), .A2(n811), .ZN(n815) );
  NAND2_X1 U900 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U901 ( .A1(n815), .A2(n814), .ZN(G295) );
  NAND2_X1 U902 ( .A1(G2078), .A2(G2084), .ZN(n816) );
  XOR2_X1 U903 ( .A(KEYINPUT20), .B(n816), .Z(n817) );
  NAND2_X1 U904 ( .A1(G2090), .A2(n817), .ZN(n818) );
  XNOR2_X1 U905 ( .A(KEYINPUT21), .B(n818), .ZN(n819) );
  NAND2_X1 U906 ( .A1(n819), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U907 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U908 ( .A1(G220), .A2(G219), .ZN(n820) );
  XNOR2_X1 U909 ( .A(KEYINPUT22), .B(n820), .ZN(n821) );
  NAND2_X1 U910 ( .A1(n821), .A2(G96), .ZN(n822) );
  NOR2_X1 U911 ( .A1(n822), .A2(G218), .ZN(n823) );
  XNOR2_X1 U912 ( .A(n823), .B(KEYINPUT83), .ZN(n837) );
  NAND2_X1 U913 ( .A1(n837), .A2(G2106), .ZN(n827) );
  NAND2_X1 U914 ( .A1(G69), .A2(G120), .ZN(n824) );
  NOR2_X1 U915 ( .A1(G237), .A2(n824), .ZN(n825) );
  NAND2_X1 U916 ( .A1(G108), .A2(n825), .ZN(n838) );
  NAND2_X1 U917 ( .A1(n838), .A2(G567), .ZN(n826) );
  NAND2_X1 U918 ( .A1(n827), .A2(n826), .ZN(n839) );
  NAND2_X1 U919 ( .A1(G661), .A2(G483), .ZN(n828) );
  XNOR2_X1 U920 ( .A(KEYINPUT84), .B(n828), .ZN(n829) );
  NOR2_X1 U921 ( .A1(n839), .A2(n829), .ZN(n836) );
  NAND2_X1 U922 ( .A1(n836), .A2(G36), .ZN(G176) );
  NAND2_X1 U923 ( .A1(n830), .A2(G2106), .ZN(n831) );
  XOR2_X1 U924 ( .A(KEYINPUT109), .B(n831), .Z(G217) );
  NAND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n832) );
  XOR2_X1 U926 ( .A(KEYINPUT110), .B(n832), .Z(n833) );
  NAND2_X1 U927 ( .A1(n833), .A2(G661), .ZN(n834) );
  XOR2_X1 U928 ( .A(KEYINPUT111), .B(n834), .Z(G259) );
  NAND2_X1 U929 ( .A1(G3), .A2(G1), .ZN(n835) );
  NAND2_X1 U930 ( .A1(n836), .A2(n835), .ZN(G188) );
  INV_X1 U932 ( .A(G120), .ZN(G236) );
  INV_X1 U933 ( .A(G96), .ZN(G221) );
  INV_X1 U934 ( .A(G69), .ZN(G235) );
  NOR2_X1 U935 ( .A1(n838), .A2(n837), .ZN(G325) );
  INV_X1 U936 ( .A(G325), .ZN(G261) );
  INV_X1 U937 ( .A(n839), .ZN(G319) );
  XOR2_X1 U938 ( .A(G2096), .B(KEYINPUT43), .Z(n841) );
  XNOR2_X1 U939 ( .A(G2067), .B(KEYINPUT42), .ZN(n840) );
  XNOR2_X1 U940 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U941 ( .A(n842), .B(G2678), .Z(n844) );
  XNOR2_X1 U942 ( .A(G2072), .B(G2090), .ZN(n843) );
  XNOR2_X1 U943 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U944 ( .A(KEYINPUT112), .B(G2100), .Z(n846) );
  XNOR2_X1 U945 ( .A(G2078), .B(G2084), .ZN(n845) );
  XNOR2_X1 U946 ( .A(n846), .B(n845), .ZN(n847) );
  XNOR2_X1 U947 ( .A(n848), .B(n847), .ZN(G227) );
  XOR2_X1 U948 ( .A(G1976), .B(G1971), .Z(n850) );
  XNOR2_X1 U949 ( .A(G1986), .B(G1966), .ZN(n849) );
  XNOR2_X1 U950 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U951 ( .A(G1981), .B(G1956), .Z(n852) );
  XNOR2_X1 U952 ( .A(G1996), .B(G1991), .ZN(n851) );
  XNOR2_X1 U953 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U954 ( .A(n854), .B(n853), .Z(n856) );
  XNOR2_X1 U955 ( .A(G2474), .B(KEYINPUT41), .ZN(n855) );
  XNOR2_X1 U956 ( .A(n856), .B(n855), .ZN(n857) );
  XNOR2_X1 U957 ( .A(KEYINPUT113), .B(n857), .ZN(n858) );
  XNOR2_X1 U958 ( .A(n858), .B(n1001), .ZN(G229) );
  NAND2_X1 U959 ( .A1(G100), .A2(n883), .ZN(n860) );
  NAND2_X1 U960 ( .A1(G112), .A2(n887), .ZN(n859) );
  NAND2_X1 U961 ( .A1(n860), .A2(n859), .ZN(n861) );
  XNOR2_X1 U962 ( .A(KEYINPUT114), .B(n861), .ZN(n866) );
  NAND2_X1 U963 ( .A1(n888), .A2(G124), .ZN(n862) );
  XNOR2_X1 U964 ( .A(n862), .B(KEYINPUT44), .ZN(n864) );
  NAND2_X1 U965 ( .A1(G136), .A2(n882), .ZN(n863) );
  NAND2_X1 U966 ( .A1(n864), .A2(n863), .ZN(n865) );
  NOR2_X1 U967 ( .A1(n866), .A2(n865), .ZN(G162) );
  XOR2_X1 U968 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n869) );
  XNOR2_X1 U969 ( .A(n867), .B(G162), .ZN(n868) );
  XNOR2_X1 U970 ( .A(n869), .B(n868), .ZN(n881) );
  NAND2_X1 U971 ( .A1(G118), .A2(n887), .ZN(n871) );
  NAND2_X1 U972 ( .A1(G130), .A2(n888), .ZN(n870) );
  NAND2_X1 U973 ( .A1(n871), .A2(n870), .ZN(n876) );
  NAND2_X1 U974 ( .A1(G142), .A2(n882), .ZN(n873) );
  NAND2_X1 U975 ( .A1(G106), .A2(n883), .ZN(n872) );
  NAND2_X1 U976 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U977 ( .A(KEYINPUT45), .B(n874), .Z(n875) );
  NOR2_X1 U978 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U979 ( .A(n877), .B(n926), .Z(n879) );
  XNOR2_X1 U980 ( .A(G164), .B(G160), .ZN(n878) );
  XNOR2_X1 U981 ( .A(n879), .B(n878), .ZN(n880) );
  XNOR2_X1 U982 ( .A(n881), .B(n880), .ZN(n896) );
  NAND2_X1 U983 ( .A1(G139), .A2(n882), .ZN(n885) );
  NAND2_X1 U984 ( .A1(G103), .A2(n883), .ZN(n884) );
  NAND2_X1 U985 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U986 ( .A(KEYINPUT115), .B(n886), .Z(n893) );
  NAND2_X1 U987 ( .A1(G115), .A2(n887), .ZN(n890) );
  NAND2_X1 U988 ( .A1(G127), .A2(n888), .ZN(n889) );
  NAND2_X1 U989 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U990 ( .A(KEYINPUT47), .B(n891), .Z(n892) );
  NOR2_X1 U991 ( .A1(n893), .A2(n892), .ZN(n934) );
  XNOR2_X1 U992 ( .A(n894), .B(n934), .ZN(n895) );
  XNOR2_X1 U993 ( .A(n896), .B(n895), .ZN(n898) );
  XOR2_X1 U994 ( .A(n898), .B(n897), .Z(n899) );
  NOR2_X1 U995 ( .A1(G37), .A2(n899), .ZN(G395) );
  XOR2_X1 U996 ( .A(G286), .B(n900), .Z(n901) );
  XNOR2_X1 U997 ( .A(n973), .B(n901), .ZN(n902) );
  XNOR2_X1 U998 ( .A(n902), .B(G171), .ZN(n903) );
  NOR2_X1 U999 ( .A1(G37), .A2(n903), .ZN(G397) );
  XNOR2_X1 U1000 ( .A(G2451), .B(G2427), .ZN(n913) );
  XOR2_X1 U1001 ( .A(G2430), .B(G2443), .Z(n905) );
  XNOR2_X1 U1002 ( .A(KEYINPUT107), .B(G2438), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(n905), .B(n904), .ZN(n909) );
  XOR2_X1 U1004 ( .A(G2435), .B(G2454), .Z(n907) );
  XNOR2_X1 U1005 ( .A(G1341), .B(G1348), .ZN(n906) );
  XNOR2_X1 U1006 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1007 ( .A(n909), .B(n908), .Z(n911) );
  XNOR2_X1 U1008 ( .A(G2446), .B(KEYINPUT108), .ZN(n910) );
  XNOR2_X1 U1009 ( .A(n911), .B(n910), .ZN(n912) );
  XNOR2_X1 U1010 ( .A(n913), .B(n912), .ZN(n914) );
  NAND2_X1 U1011 ( .A1(n914), .A2(G14), .ZN(n920) );
  NAND2_X1 U1012 ( .A1(G319), .A2(n920), .ZN(n917) );
  NOR2_X1 U1013 ( .A1(G227), .A2(G229), .ZN(n915) );
  XNOR2_X1 U1014 ( .A(KEYINPUT49), .B(n915), .ZN(n916) );
  NOR2_X1 U1015 ( .A1(n917), .A2(n916), .ZN(n919) );
  NOR2_X1 U1016 ( .A1(G395), .A2(G397), .ZN(n918) );
  NAND2_X1 U1017 ( .A1(n919), .A2(n918), .ZN(G225) );
  INV_X1 U1018 ( .A(G225), .ZN(G308) );
  INV_X1 U1019 ( .A(G108), .ZN(G238) );
  INV_X1 U1020 ( .A(n920), .ZN(G401) );
  XNOR2_X1 U1021 ( .A(KEYINPUT52), .B(KEYINPUT119), .ZN(n946) );
  XOR2_X1 U1022 ( .A(G2090), .B(G162), .Z(n921) );
  NOR2_X1 U1023 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1024 ( .A(KEYINPUT51), .B(n923), .ZN(n924) );
  XNOR2_X1 U1025 ( .A(n924), .B(KEYINPUT117), .ZN(n944) );
  XNOR2_X1 U1026 ( .A(G2084), .B(G160), .ZN(n925) );
  XNOR2_X1 U1027 ( .A(n925), .B(KEYINPUT116), .ZN(n929) );
  NOR2_X1 U1028 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1029 ( .A1(n929), .A2(n928), .ZN(n930) );
  NOR2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(n933) );
  NAND2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(n942) );
  XOR2_X1 U1032 ( .A(G2072), .B(n934), .Z(n936) );
  XOR2_X1 U1033 ( .A(G164), .B(G2078), .Z(n935) );
  NOR2_X1 U1034 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1035 ( .A(n937), .B(KEYINPUT118), .ZN(n938) );
  XNOR2_X1 U1036 ( .A(n938), .B(KEYINPUT50), .ZN(n940) );
  NAND2_X1 U1037 ( .A1(n940), .A2(n939), .ZN(n941) );
  NOR2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1039 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1040 ( .A(n946), .B(n945), .ZN(n947) );
  INV_X1 U1041 ( .A(KEYINPUT55), .ZN(n969) );
  NAND2_X1 U1042 ( .A1(n947), .A2(n969), .ZN(n948) );
  NAND2_X1 U1043 ( .A1(n948), .A2(G29), .ZN(n1030) );
  XNOR2_X1 U1044 ( .A(G25), .B(n949), .ZN(n950) );
  NAND2_X1 U1045 ( .A1(n950), .A2(G28), .ZN(n960) );
  XNOR2_X1 U1046 ( .A(G2067), .B(G26), .ZN(n952) );
  XNOR2_X1 U1047 ( .A(G33), .B(G2072), .ZN(n951) );
  NOR2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n958) );
  XOR2_X1 U1049 ( .A(n953), .B(G32), .Z(n956) );
  XOR2_X1 U1050 ( .A(n954), .B(G27), .Z(n955) );
  NOR2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n959) );
  NOR2_X1 U1053 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1054 ( .A(KEYINPUT53), .B(n961), .Z(n962) );
  XOR2_X1 U1055 ( .A(KEYINPUT120), .B(n962), .Z(n964) );
  XNOR2_X1 U1056 ( .A(G2090), .B(G35), .ZN(n963) );
  NOR2_X1 U1057 ( .A1(n964), .A2(n963), .ZN(n967) );
  XOR2_X1 U1058 ( .A(G2084), .B(G34), .Z(n965) );
  XNOR2_X1 U1059 ( .A(KEYINPUT54), .B(n965), .ZN(n966) );
  NAND2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1061 ( .A(n969), .B(n968), .ZN(n971) );
  INV_X1 U1062 ( .A(G29), .ZN(n970) );
  NAND2_X1 U1063 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1064 ( .A1(G11), .A2(n972), .ZN(n1028) );
  XNOR2_X1 U1065 ( .A(KEYINPUT56), .B(G16), .ZN(n1000) );
  XNOR2_X1 U1066 ( .A(G1348), .B(KEYINPUT122), .ZN(n974) );
  XNOR2_X1 U1067 ( .A(n974), .B(n973), .ZN(n976) );
  XOR2_X1 U1068 ( .A(G171), .B(G1961), .Z(n975) );
  NOR2_X1 U1069 ( .A1(n976), .A2(n975), .ZN(n998) );
  XNOR2_X1 U1070 ( .A(n977), .B(G1341), .ZN(n990) );
  XOR2_X1 U1071 ( .A(G299), .B(G1956), .Z(n979) );
  XNOR2_X1 U1072 ( .A(G166), .B(G1971), .ZN(n978) );
  NAND2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n984) );
  NAND2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1075 ( .A(KEYINPUT123), .B(n982), .Z(n983) );
  NOR2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1077 ( .A(KEYINPUT124), .B(n985), .Z(n986) );
  NOR2_X1 U1078 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1079 ( .A(KEYINPUT125), .B(n988), .Z(n989) );
  NAND2_X1 U1080 ( .A1(n990), .A2(n989), .ZN(n996) );
  XOR2_X1 U1081 ( .A(G168), .B(G1966), .Z(n991) );
  NOR2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1083 ( .A(KEYINPUT57), .B(n993), .Z(n994) );
  XNOR2_X1 U1084 ( .A(n994), .B(KEYINPUT121), .ZN(n995) );
  NOR2_X1 U1085 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1086 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1087 ( .A1(n1000), .A2(n999), .ZN(n1026) );
  XNOR2_X1 U1088 ( .A(G5), .B(n1001), .ZN(n1021) );
  XOR2_X1 U1089 ( .A(G1966), .B(G21), .Z(n1011) );
  XNOR2_X1 U1090 ( .A(G1348), .B(KEYINPUT59), .ZN(n1002) );
  XNOR2_X1 U1091 ( .A(n1002), .B(G4), .ZN(n1006) );
  XNOR2_X1 U1092 ( .A(G1341), .B(G19), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(G1981), .B(G6), .ZN(n1003) );
  NOR2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1008) );
  XNOR2_X1 U1096 ( .A(G20), .B(G1956), .ZN(n1007) );
  NOR2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1098 ( .A(n1009), .B(KEYINPUT60), .ZN(n1010) );
  NAND2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1100 ( .A(KEYINPUT126), .B(n1012), .ZN(n1019) );
  XNOR2_X1 U1101 ( .A(G1986), .B(G24), .ZN(n1014) );
  XNOR2_X1 U1102 ( .A(G1971), .B(G22), .ZN(n1013) );
  NOR2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1016) );
  XOR2_X1 U1104 ( .A(G1976), .B(G23), .Z(n1015) );
  NAND2_X1 U1105 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1106 ( .A(KEYINPUT58), .B(n1017), .ZN(n1018) );
  NOR2_X1 U1107 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1109 ( .A(KEYINPUT61), .B(n1022), .ZN(n1023) );
  NOR2_X1 U1110 ( .A1(G16), .A2(n1023), .ZN(n1024) );
  XNOR2_X1 U1111 ( .A(n1024), .B(KEYINPUT127), .ZN(n1025) );
  NAND2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1113 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1114 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1115 ( .A(KEYINPUT62), .B(n1031), .Z(G311) );
  INV_X1 U1116 ( .A(G311), .ZN(G150) );
endmodule

