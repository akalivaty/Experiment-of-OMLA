//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 0 1 1 1 1 0 1 1 0 1 0 1 0 1 0 0 0 0 0 0 0 0 0 1 1 1 0 0 0 0 0 0 0 0 1 1 0 1 1 0 1 0 1 0 1 0 0 1 1 0 1 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n817, new_n818, new_n819, new_n821,
    new_n822, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n958, new_n959;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202));
  XOR2_X1   g001(.A(new_n202), .B(KEYINPUT13), .Z(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G15gat), .B(G22gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT16), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n205), .B1(new_n206), .B2(G1gat), .ZN(new_n207));
  INV_X1    g006(.A(G8gat), .ZN(new_n208));
  OAI221_X1 g007(.A(new_n207), .B1(KEYINPUT93), .B2(new_n208), .C1(G1gat), .C2(new_n205), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(KEYINPUT93), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n209), .B(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT92), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT15), .ZN(new_n214));
  OR2_X1    g013(.A1(new_n214), .A2(KEYINPUT90), .ZN(new_n215));
  AOI22_X1  g014(.A1(new_n214), .A2(KEYINPUT90), .B1(G43gat), .B2(G50gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G50gat), .ZN(new_n218));
  XNOR2_X1  g017(.A(KEYINPUT91), .B(G43gat), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  OR2_X1    g019(.A1(G43gat), .A2(G50gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(G43gat), .A2(G50gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT15), .ZN(new_n224));
  OR3_X1    g023(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G29gat), .A2(G36gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n224), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n213), .B1(new_n220), .B2(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n214), .B1(new_n221), .B2(new_n222), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n231), .B1(G29gat), .B2(G36gat), .ZN(new_n232));
  XOR2_X1   g031(.A(KEYINPUT91), .B(G43gat), .Z(new_n233));
  OAI211_X1 g032(.A(new_n215), .B(new_n216), .C1(new_n233), .C2(G50gat), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n232), .A2(new_n234), .A3(KEYINPUT92), .A4(new_n227), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n230), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n225), .A2(KEYINPUT89), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(new_n226), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n225), .A2(KEYINPUT89), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n228), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(new_n231), .ZN(new_n241));
  AND2_X1   g040(.A1(new_n236), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n212), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n236), .A2(new_n241), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n211), .A2(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n204), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT17), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n236), .A2(new_n247), .A3(new_n241), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n247), .B1(new_n236), .B2(new_n241), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n212), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n250), .A2(new_n202), .A3(new_n245), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT18), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n246), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G113gat), .B(G141gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT87), .B(G197gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(KEYINPUT11), .B(G169gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  XOR2_X1   g057(.A(KEYINPUT88), .B(KEYINPUT12), .Z(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n250), .A2(KEYINPUT18), .A3(new_n202), .A4(new_n245), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n253), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n260), .B1(new_n253), .B2(new_n261), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT94), .ZN(new_n265));
  NOR3_X1   g064(.A1(new_n263), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n253), .A2(new_n261), .ZN(new_n267));
  INV_X1    g066(.A(new_n260), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(KEYINPUT94), .B1(new_n269), .B2(new_n262), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n266), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT74), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT71), .ZN(new_n274));
  NAND3_X1  g073(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n275));
  AOI21_X1  g074(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n276));
  OAI221_X1 g075(.A(new_n275), .B1(G183gat), .B2(G190gat), .C1(new_n276), .C2(KEYINPUT65), .ZN(new_n277));
  AND2_X1   g076(.A1(new_n276), .A2(KEYINPUT65), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT66), .ZN(new_n279));
  NOR2_X1   g078(.A1(G169gat), .A2(G176gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT23), .ZN(new_n281));
  OAI22_X1  g080(.A1(new_n277), .A2(new_n278), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(G169gat), .A2(G176gat), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n280), .B1(KEYINPUT23), .B2(new_n285), .ZN(new_n286));
  OR2_X1    g085(.A1(new_n286), .A2(new_n279), .ZN(new_n287));
  INV_X1    g086(.A(new_n276), .ZN(new_n288));
  INV_X1    g087(.A(G183gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT67), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT67), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(G183gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n288), .B(new_n275), .C1(new_n293), .C2(G190gat), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT25), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n286), .A2(new_n295), .ZN(new_n296));
  AOI22_X1  g095(.A1(new_n287), .A2(new_n283), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n281), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n284), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT27), .B(G183gat), .ZN(new_n300));
  INV_X1    g099(.A(G190gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n300), .A2(KEYINPUT28), .A3(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT68), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT27), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n304), .B1(new_n290), .B2(new_n292), .ZN(new_n305));
  NOR2_X1   g104(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n306));
  OAI211_X1 g105(.A(new_n303), .B(new_n301), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT28), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n306), .ZN(new_n310));
  XNOR2_X1  g109(.A(KEYINPUT67), .B(G183gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n310), .B1(new_n311), .B2(new_n304), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n303), .B1(new_n312), .B2(new_n301), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n302), .B1(new_n309), .B2(new_n313), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n280), .A2(KEYINPUT26), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(new_n285), .ZN(new_n316));
  AOI22_X1  g115(.A1(new_n280), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT69), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n318), .B(new_n319), .ZN(new_n320));
  AND3_X1   g119(.A1(new_n314), .A2(KEYINPUT70), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT70), .B1(new_n314), .B2(new_n320), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n299), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(G113gat), .B(G120gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n324), .A2(KEYINPUT1), .ZN(new_n325));
  XNOR2_X1  g124(.A(G127gat), .B(G134gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n326), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n328), .B1(KEYINPUT1), .B2(new_n324), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n323), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n330), .ZN(new_n332));
  OAI211_X1 g131(.A(new_n332), .B(new_n299), .C1(new_n321), .C2(new_n322), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(G227gat), .A2(G233gat), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n274), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  AOI211_X1 g136(.A(KEYINPUT71), .B(new_n335), .C1(new_n331), .C2(new_n333), .ZN(new_n338));
  OAI21_X1  g137(.A(KEYINPUT32), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  XOR2_X1   g138(.A(KEYINPUT72), .B(KEYINPUT33), .Z(new_n340));
  OAI21_X1  g139(.A(new_n340), .B1(new_n337), .B2(new_n338), .ZN(new_n341));
  XOR2_X1   g140(.A(G15gat), .B(G43gat), .Z(new_n342));
  XNOR2_X1  g141(.A(G71gat), .B(G99gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n342), .B(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n339), .A2(new_n341), .A3(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n344), .ZN(new_n346));
  OAI221_X1 g145(.A(KEYINPUT32), .B1(new_n340), .B2(new_n346), .C1(new_n337), .C2(new_n338), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n331), .A2(new_n335), .A3(new_n333), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT34), .B1(new_n336), .B2(KEYINPUT73), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n349), .B(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n348), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n345), .A2(new_n351), .A3(new_n347), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n273), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n345), .A2(new_n351), .A3(new_n347), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(new_n273), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(KEYINPUT85), .B1(new_n355), .B2(new_n358), .ZN(new_n359));
  AND3_X1   g158(.A1(new_n345), .A2(new_n351), .A3(new_n347), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n351), .B1(new_n345), .B2(new_n347), .ZN(new_n361));
  OAI21_X1  g160(.A(KEYINPUT74), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT85), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n362), .A2(new_n363), .A3(new_n357), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n359), .A2(new_n364), .ZN(new_n365));
  OR2_X1    g164(.A1(KEYINPUT79), .A2(G148gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(KEYINPUT79), .A2(G148gat), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n366), .A2(G141gat), .A3(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(G148gat), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n369), .A2(G141gat), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  OR3_X1    g170(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(G155gat), .A2(G162gat), .ZN(new_n373));
  AOI22_X1  g172(.A1(new_n368), .A2(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  XOR2_X1   g173(.A(G155gat), .B(G162gat), .Z(new_n375));
  XNOR2_X1  g174(.A(G141gat), .B(G148gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(KEYINPUT77), .B(KEYINPUT2), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n375), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT78), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n375), .B(KEYINPUT78), .C1(new_n376), .C2(new_n377), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n374), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(new_n332), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT4), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n382), .A2(KEYINPUT4), .A3(new_n332), .ZN(new_n386));
  INV_X1    g185(.A(new_n374), .ZN(new_n387));
  INV_X1    g186(.A(new_n381), .ZN(new_n388));
  OR2_X1    g187(.A1(KEYINPUT77), .A2(KEYINPUT2), .ZN(new_n389));
  NAND2_X1  g188(.A1(KEYINPUT77), .A2(KEYINPUT2), .ZN(new_n390));
  INV_X1    g189(.A(G141gat), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n391), .A2(G148gat), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n389), .B(new_n390), .C1(new_n370), .C2(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT78), .B1(new_n393), .B2(new_n375), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n387), .B1(new_n388), .B2(new_n394), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n395), .A2(KEYINPUT3), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT3), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n330), .B1(new_n382), .B2(new_n397), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n385), .B(new_n386), .C1(new_n396), .C2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(G225gat), .A2(G233gat), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT5), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n395), .A2(new_n330), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n400), .B1(new_n403), .B2(new_n383), .ZN(new_n404));
  OAI22_X1  g203(.A1(new_n399), .A2(new_n401), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  AND2_X1   g204(.A1(new_n385), .A2(new_n386), .ZN(new_n406));
  OR2_X1    g205(.A1(new_n398), .A2(new_n396), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n406), .A2(KEYINPUT5), .A3(new_n407), .A4(new_n400), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  XOR2_X1   g208(.A(G1gat), .B(G29gat), .Z(new_n410));
  XNOR2_X1  g209(.A(G57gat), .B(G85gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n410), .B(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n413));
  XOR2_X1   g212(.A(new_n412), .B(new_n413), .Z(new_n414));
  NAND2_X1  g213(.A1(new_n409), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT6), .ZN(new_n416));
  INV_X1    g215(.A(new_n414), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n405), .A2(new_n408), .A3(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n415), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n405), .A2(new_n408), .A3(KEYINPUT6), .A4(new_n417), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  AND2_X1   g221(.A1(G226gat), .A2(G233gat), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n423), .B(new_n299), .C1(new_n321), .C2(new_n322), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n314), .A2(new_n320), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(new_n299), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n423), .A2(KEYINPUT29), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n424), .A2(new_n428), .ZN(new_n429));
  AND2_X1   g228(.A1(G211gat), .A2(G218gat), .ZN(new_n430));
  AND2_X1   g229(.A1(G197gat), .A2(G204gat), .ZN(new_n431));
  NOR2_X1   g230(.A1(G197gat), .A2(G204gat), .ZN(new_n432));
  OAI22_X1  g231(.A1(KEYINPUT22), .A2(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  XOR2_X1   g232(.A(G211gat), .B(G218gat), .Z(new_n434));
  XOR2_X1   g233(.A(new_n433), .B(new_n434), .Z(new_n435));
  INV_X1    g234(.A(KEYINPUT75), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n433), .A2(KEYINPUT75), .A3(new_n434), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n429), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n425), .A2(new_n423), .A3(new_n299), .ZN(new_n442));
  INV_X1    g241(.A(new_n299), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT70), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n425), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n314), .A2(KEYINPUT70), .A3(new_n320), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n443), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n427), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n442), .B(new_n439), .C1(new_n447), .C2(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n441), .A2(KEYINPUT76), .A3(new_n449), .ZN(new_n450));
  AOI211_X1 g249(.A(KEYINPUT76), .B(new_n439), .C1(new_n424), .C2(new_n428), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g252(.A(G8gat), .B(G36gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(G64gat), .B(G92gat), .ZN(new_n455));
  XOR2_X1   g254(.A(new_n454), .B(new_n455), .Z(new_n456));
  NAND2_X1  g255(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT76), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n458), .B1(new_n429), .B2(new_n440), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n451), .B1(new_n459), .B2(new_n449), .ZN(new_n460));
  INV_X1    g259(.A(new_n456), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n457), .A2(new_n462), .A3(KEYINPUT30), .ZN(new_n463));
  OR3_X1    g262(.A1(new_n460), .A2(KEYINPUT30), .A3(new_n461), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n422), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n396), .A2(KEYINPUT29), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n467), .A2(new_n440), .ZN(new_n468));
  OR2_X1    g267(.A1(new_n468), .A2(KEYINPUT81), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(KEYINPUT81), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n397), .B1(new_n435), .B2(KEYINPUT29), .ZN(new_n471));
  AOI22_X1  g270(.A1(new_n471), .A2(new_n395), .B1(G228gat), .B2(G233gat), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n469), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  OR2_X1    g272(.A1(new_n439), .A2(KEYINPUT29), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n382), .B1(new_n474), .B2(new_n397), .ZN(new_n475));
  OAI211_X1 g274(.A(G228gat), .B(G233gat), .C1(new_n475), .C2(new_n468), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(KEYINPUT31), .B(G50gat), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  XNOR2_X1  g278(.A(G78gat), .B(G106gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n480), .B(G22gat), .ZN(new_n481));
  INV_X1    g280(.A(new_n478), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n473), .A2(new_n476), .A3(new_n482), .ZN(new_n483));
  AND3_X1   g282(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n481), .B1(new_n479), .B2(new_n483), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NOR3_X1   g286(.A1(new_n466), .A2(new_n487), .A3(KEYINPUT35), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n365), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n353), .A2(new_n465), .A3(new_n486), .A4(new_n354), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT35), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT86), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n490), .A2(KEYINPUT86), .A3(KEYINPUT35), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n489), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT37), .ZN(new_n497));
  INV_X1    g296(.A(new_n442), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n498), .B1(new_n323), .B2(new_n427), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n497), .B1(new_n499), .B2(new_n440), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n429), .A2(new_n439), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT38), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  XNOR2_X1  g301(.A(KEYINPUT82), .B(KEYINPUT37), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n502), .B(new_n461), .C1(new_n460), .C2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT83), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n453), .A2(new_n503), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n508), .A2(KEYINPUT83), .A3(new_n461), .A4(new_n502), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n461), .B1(new_n450), .B2(new_n452), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n421), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n507), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT84), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n507), .A2(new_n509), .A3(new_n511), .A4(KEYINPUT84), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n508), .A2(new_n461), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n453), .A2(new_n497), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT38), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n514), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  AND2_X1   g318(.A1(new_n463), .A2(new_n464), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n399), .A2(new_n401), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n403), .A2(new_n383), .A3(new_n400), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n521), .A2(KEYINPUT39), .A3(new_n522), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n523), .B(new_n414), .C1(KEYINPUT39), .C2(new_n521), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT40), .ZN(new_n525));
  OR2_X1    g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(new_n525), .ZN(new_n527));
  AND3_X1   g326(.A1(new_n526), .A2(new_n418), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n487), .B1(new_n520), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n519), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n466), .A2(new_n487), .ZN(new_n531));
  AOI21_X1  g330(.A(KEYINPUT36), .B1(new_n362), .B2(new_n357), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT36), .ZN(new_n533));
  NOR3_X1   g332(.A1(new_n360), .A2(new_n361), .A3(new_n533), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n530), .B(new_n531), .C1(new_n532), .C2(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n272), .B1(new_n496), .B2(new_n535), .ZN(new_n536));
  XOR2_X1   g335(.A(G57gat), .B(G64gat), .Z(new_n537));
  INV_X1    g336(.A(KEYINPUT9), .ZN(new_n538));
  INV_X1    g337(.A(G71gat), .ZN(new_n539));
  INV_X1    g338(.A(G78gat), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(G71gat), .B(G78gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n544), .A2(KEYINPUT21), .ZN(new_n545));
  AND2_X1   g344(.A1(G231gat), .A2(G233gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  XOR2_X1   g346(.A(G127gat), .B(G155gat), .Z(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT20), .ZN(new_n549));
  XOR2_X1   g348(.A(new_n547), .B(new_n549), .Z(new_n550));
  XNOR2_X1  g349(.A(G183gat), .B(G211gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n211), .B1(KEYINPUT21), .B2(new_n544), .ZN(new_n553));
  XNOR2_X1  g352(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(new_n552), .B(new_n555), .Z(new_n556));
  XOR2_X1   g355(.A(G99gat), .B(G106gat), .Z(new_n557));
  NAND2_X1  g356(.A1(G99gat), .A2(G106gat), .ZN(new_n558));
  INV_X1    g357(.A(G85gat), .ZN(new_n559));
  INV_X1    g358(.A(G92gat), .ZN(new_n560));
  AOI22_X1  g359(.A1(KEYINPUT8), .A2(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(KEYINPUT98), .ZN(new_n562));
  NAND2_X1  g361(.A1(KEYINPUT97), .A2(KEYINPUT7), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n563), .A2(G85gat), .A3(G92gat), .ZN(new_n564));
  NOR2_X1   g363(.A1(KEYINPUT97), .A2(KEYINPUT7), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n557), .B1(new_n562), .B2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT99), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT98), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n561), .B(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n565), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n564), .B(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n557), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n570), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n567), .A2(new_n568), .A3(new_n574), .ZN(new_n575));
  OAI211_X1 g374(.A(KEYINPUT99), .B(new_n557), .C1(new_n562), .C2(new_n566), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(new_n244), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT41), .ZN(new_n579));
  NAND2_X1  g378(.A1(G232gat), .A2(G233gat), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n248), .A2(new_n249), .ZN(new_n581));
  OAI221_X1 g380(.A(new_n578), .B1(new_n579), .B2(new_n580), .C1(new_n581), .C2(new_n577), .ZN(new_n582));
  XNOR2_X1  g381(.A(G190gat), .B(G218gat), .ZN(new_n583));
  OR2_X1    g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(KEYINPUT100), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n580), .A2(new_n579), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT96), .ZN(new_n587));
  XNOR2_X1  g386(.A(G134gat), .B(G162gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n582), .A2(new_n583), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n584), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n585), .A2(new_n584), .A3(new_n591), .A4(new_n589), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n556), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G120gat), .B(G148gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(G176gat), .B(G204gat), .ZN(new_n599));
  XOR2_X1   g398(.A(new_n598), .B(new_n599), .Z(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(new_n542), .B(new_n543), .Z(new_n602));
  NAND3_X1  g401(.A1(new_n575), .A2(new_n576), .A3(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT10), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n567), .A2(new_n544), .A3(new_n574), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT101), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n603), .A2(KEYINPUT101), .A3(new_n604), .A4(new_n605), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n602), .A2(new_n604), .ZN(new_n610));
  AOI22_X1  g409(.A1(new_n608), .A2(new_n609), .B1(new_n577), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(G230gat), .A2(G233gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT103), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n613), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n615), .B1(new_n603), .B2(new_n605), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n601), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT104), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n608), .A2(new_n609), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n577), .A2(new_n610), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(KEYINPUT102), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT102), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n611), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n622), .A2(new_n624), .A3(new_n615), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n616), .A2(new_n601), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n618), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n615), .B1(new_n611), .B2(new_n623), .ZN(new_n628));
  AND3_X1   g427(.A1(new_n619), .A2(new_n623), .A3(new_n620), .ZN(new_n629));
  OAI211_X1 g428(.A(new_n618), .B(new_n626), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n617), .B1(new_n627), .B2(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n597), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n536), .A2(KEYINPUT105), .A3(new_n633), .ZN(new_n634));
  AOI22_X1  g433(.A1(new_n365), .A2(new_n488), .B1(new_n493), .B2(new_n494), .ZN(new_n635));
  INV_X1    g434(.A(new_n535), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n271), .B(new_n633), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT105), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n634), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(new_n422), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(G1gat), .ZN(G1324gat));
  INV_X1    g441(.A(KEYINPUT106), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n640), .A2(new_n520), .ZN(new_n644));
  XOR2_X1   g443(.A(KEYINPUT16), .B(G8gat), .Z(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n643), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(KEYINPUT42), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT42), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n643), .B(new_n649), .C1(new_n644), .C2(new_n646), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n644), .A2(G8gat), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n648), .A2(new_n650), .A3(new_n651), .ZN(G1325gat));
  INV_X1    g451(.A(new_n640), .ZN(new_n653));
  INV_X1    g452(.A(new_n365), .ZN(new_n654));
  OR3_X1    g453(.A1(new_n653), .A2(G15gat), .A3(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(KEYINPUT107), .B1(new_n532), .B2(new_n534), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n533), .B1(new_n355), .B2(new_n358), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT107), .ZN(new_n658));
  INV_X1    g457(.A(new_n534), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(G15gat), .B1(new_n653), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n655), .A2(new_n662), .ZN(G1326gat));
  AOI21_X1  g462(.A(KEYINPUT105), .B1(new_n536), .B2(new_n633), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n637), .A2(new_n638), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n487), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(KEYINPUT108), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT108), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n640), .A2(new_n668), .A3(new_n487), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT43), .B(G22gat), .ZN(new_n670));
  AND3_X1   g469(.A1(new_n667), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n670), .B1(new_n667), .B2(new_n669), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n671), .A2(new_n672), .ZN(G1327gat));
  INV_X1    g472(.A(new_n556), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n593), .A2(new_n594), .ZN(new_n675));
  NOR3_X1   g474(.A1(new_n674), .A2(new_n632), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n536), .A2(new_n676), .ZN(new_n677));
  NOR3_X1   g476(.A1(new_n677), .A2(G29gat), .A3(new_n421), .ZN(new_n678));
  XOR2_X1   g477(.A(new_n678), .B(KEYINPUT45), .Z(new_n679));
  NAND2_X1  g478(.A1(new_n530), .A2(new_n531), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n680), .B1(new_n656), .B2(new_n660), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n595), .B1(new_n681), .B2(new_n635), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OAI211_X1 g483(.A(KEYINPUT44), .B(new_n595), .C1(new_n635), .C2(new_n636), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n632), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n269), .A2(new_n262), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n687), .A2(new_n556), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT109), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(G29gat), .B1(new_n691), .B2(new_n421), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n679), .A2(new_n692), .ZN(G1328gat));
  INV_X1    g492(.A(new_n520), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n677), .A2(G36gat), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT46), .ZN(new_n696));
  OAI21_X1  g495(.A(G36gat), .B1(new_n691), .B2(new_n694), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(G1329gat));
  INV_X1    g497(.A(new_n661), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n684), .A2(new_n699), .A3(new_n685), .A4(new_n690), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(new_n233), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n654), .A2(new_n233), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n536), .A2(new_n676), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(KEYINPUT47), .B1(new_n704), .B2(KEYINPUT110), .ZN(new_n705));
  INV_X1    g504(.A(new_n703), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n706), .B1(new_n700), .B2(new_n233), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT110), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT47), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n705), .A2(new_n710), .ZN(G1330gat));
  NAND4_X1  g510(.A1(new_n684), .A2(new_n487), .A3(new_n685), .A4(new_n690), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(G50gat), .ZN(new_n713));
  AOI21_X1  g512(.A(KEYINPUT48), .B1(new_n713), .B2(KEYINPUT111), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n487), .A2(new_n218), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n713), .B1(new_n677), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  OAI221_X1 g516(.A(new_n713), .B1(KEYINPUT111), .B2(KEYINPUT48), .C1(new_n677), .C2(new_n715), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(G1331gat));
  OAI21_X1  g518(.A(new_n496), .B1(new_n699), .B2(new_n680), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n597), .A2(new_n688), .A3(new_n687), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(new_n422), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g524(.A1(new_n723), .A2(new_n520), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n726), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n727));
  XOR2_X1   g526(.A(KEYINPUT49), .B(G64gat), .Z(new_n728));
  OAI21_X1  g527(.A(new_n727), .B1(new_n726), .B2(new_n728), .ZN(G1333gat));
  OAI21_X1  g528(.A(G71gat), .B1(new_n722), .B2(new_n661), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n365), .A2(new_n539), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n730), .B1(new_n722), .B2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT50), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n732), .B(new_n733), .ZN(G1334gat));
  NAND2_X1  g533(.A1(new_n723), .A2(new_n487), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g535(.A1(new_n674), .A2(new_n687), .A3(new_n688), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n686), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(G85gat), .B1(new_n738), .B2(new_n421), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n674), .A2(new_n688), .ZN(new_n740));
  OAI211_X1 g539(.A(new_n595), .B(new_n740), .C1(new_n681), .C2(new_n635), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT51), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n741), .A2(new_n742), .ZN(new_n744));
  OR2_X1    g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(new_n632), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n422), .A2(new_n559), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n739), .B1(new_n746), .B2(new_n747), .ZN(G1336gat));
  NOR3_X1   g547(.A1(new_n694), .A2(new_n687), .A3(G92gat), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT52), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n684), .A2(new_n520), .A3(new_n685), .A4(new_n737), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(G92gat), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n750), .A2(new_n751), .A3(new_n753), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n749), .B(KEYINPUT112), .ZN(new_n755));
  AOI22_X1  g554(.A1(new_n745), .A2(new_n755), .B1(new_n752), .B2(G92gat), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n754), .B1(new_n756), .B2(new_n751), .ZN(G1337gat));
  OAI21_X1  g556(.A(G99gat), .B1(new_n738), .B2(new_n661), .ZN(new_n758));
  OR2_X1    g557(.A1(new_n654), .A2(G99gat), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n758), .B1(new_n746), .B2(new_n759), .ZN(G1338gat));
  NOR2_X1   g559(.A1(new_n486), .A2(G106gat), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n632), .B(new_n761), .C1(new_n743), .C2(new_n744), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n684), .A2(new_n487), .A3(new_n685), .A4(new_n737), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(G106gat), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n762), .A2(KEYINPUT113), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n765), .A2(new_n766), .A3(KEYINPUT53), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT53), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n762), .B(new_n764), .C1(KEYINPUT113), .C2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n769), .ZN(G1339gat));
  NOR3_X1   g569(.A1(new_n597), .A2(new_n688), .A3(new_n632), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n243), .A2(new_n245), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n250), .A2(new_n245), .ZN(new_n773));
  INV_X1    g572(.A(new_n202), .ZN(new_n774));
  AOI22_X1  g573(.A1(new_n772), .A2(new_n204), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n263), .B1(new_n258), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n632), .A2(new_n777), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n626), .B1(new_n628), .B2(new_n629), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(KEYINPUT104), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(new_n630), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT54), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n782), .B1(new_n611), .B2(new_n613), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n783), .B1(new_n628), .B2(new_n629), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n600), .B1(new_n614), .B2(new_n782), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n784), .A2(KEYINPUT55), .A3(new_n785), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n781), .A2(new_n788), .A3(new_n688), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n778), .A2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT114), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n595), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n778), .A2(new_n790), .A3(KEYINPUT114), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n781), .A2(new_n788), .A3(new_n789), .ZN(new_n796));
  INV_X1    g595(.A(new_n777), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n796), .A2(new_n675), .A3(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n771), .B1(new_n800), .B2(new_n556), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n801), .A2(new_n487), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n520), .A2(new_n421), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n802), .A2(new_n365), .A3(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(G113gat), .B1(new_n804), .B2(new_n272), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n801), .A2(new_n421), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n360), .A2(new_n361), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n486), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n810), .A2(new_n520), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(new_n688), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n813), .A2(G113gat), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n814), .B(KEYINPUT115), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n805), .B1(new_n812), .B2(new_n815), .ZN(G1340gat));
  INV_X1    g615(.A(G120gat), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n804), .A2(new_n817), .A3(new_n687), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n811), .A2(new_n632), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n818), .B1(new_n819), .B2(new_n817), .ZN(G1341gat));
  OAI21_X1  g619(.A(G127gat), .B1(new_n804), .B2(new_n556), .ZN(new_n821));
  OR2_X1    g620(.A1(new_n556), .A2(G127gat), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n821), .B1(new_n812), .B2(new_n822), .ZN(G1342gat));
  NOR2_X1   g622(.A1(new_n675), .A2(new_n520), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n824), .B(KEYINPUT116), .ZN(new_n825));
  OR3_X1    g624(.A1(new_n810), .A2(G134gat), .A3(new_n825), .ZN(new_n826));
  OR2_X1    g625(.A1(new_n826), .A2(KEYINPUT56), .ZN(new_n827));
  OAI21_X1  g626(.A(G134gat), .B1(new_n804), .B2(new_n675), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(KEYINPUT56), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(G1343gat));
  INV_X1    g629(.A(KEYINPUT119), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n831), .B1(new_n801), .B2(new_n421), .ZN(new_n832));
  INV_X1    g631(.A(new_n771), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n798), .B1(new_n793), .B2(new_n794), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n833), .B1(new_n834), .B2(new_n674), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n835), .A2(KEYINPUT119), .A3(new_n422), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n699), .A2(new_n486), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n832), .A2(new_n694), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n271), .A2(new_n391), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n803), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n841), .B1(new_n656), .B2(new_n660), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n835), .A2(new_n487), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n486), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n271), .A2(new_n781), .A3(new_n788), .A4(new_n789), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n595), .B1(new_n847), .B2(new_n778), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n556), .B1(new_n848), .B2(new_n798), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT117), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n771), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI211_X1 g650(.A(KEYINPUT117), .B(new_n556), .C1(new_n848), .C2(new_n798), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n846), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OAI22_X1  g652(.A1(new_n843), .A2(KEYINPUT57), .B1(new_n853), .B2(KEYINPUT118), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(KEYINPUT118), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  OAI211_X1 g655(.A(new_n688), .B(new_n842), .C1(new_n854), .C2(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n840), .B1(new_n857), .B2(G141gat), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT58), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n661), .A2(new_n803), .ZN(new_n860));
  AOI21_X1  g659(.A(KEYINPUT57), .B1(new_n835), .B2(new_n487), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n849), .A2(new_n850), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n862), .A2(new_n833), .A3(new_n852), .ZN(new_n863));
  AOI21_X1  g662(.A(KEYINPUT118), .B1(new_n863), .B2(new_n845), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n860), .B1(new_n865), .B2(new_n855), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n391), .B1(new_n866), .B2(new_n271), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n859), .B1(new_n838), .B2(new_n839), .ZN(new_n868));
  OAI22_X1  g667(.A1(new_n858), .A2(new_n859), .B1(new_n867), .B2(new_n868), .ZN(G1344gat));
  NAND2_X1  g668(.A1(new_n366), .A2(new_n367), .ZN(new_n870));
  OR3_X1    g669(.A1(new_n838), .A2(new_n870), .A3(new_n687), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT59), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT120), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n687), .B1(new_n842), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n860), .A2(KEYINPUT120), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n847), .A2(new_n778), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n675), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n674), .B1(new_n878), .B2(new_n799), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n597), .A2(new_n271), .A3(new_n632), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n487), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AOI22_X1  g680(.A1(new_n835), .A2(new_n845), .B1(new_n881), .B2(new_n844), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n876), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n369), .B1(new_n883), .B2(KEYINPUT121), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT121), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n885), .B1(new_n876), .B2(new_n882), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n872), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n870), .A2(new_n872), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n888), .B1(new_n866), .B2(new_n632), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n871), .B1(new_n887), .B2(new_n889), .ZN(G1345gat));
  INV_X1    g689(.A(G155gat), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n891), .B1(new_n866), .B2(new_n674), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n838), .A2(G155gat), .A3(new_n556), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n892), .A2(new_n893), .ZN(G1346gat));
  INV_X1    g693(.A(G162gat), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n895), .B1(new_n866), .B2(new_n595), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n836), .A2(new_n837), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n825), .A2(G162gat), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n897), .A2(new_n832), .A3(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(KEYINPUT122), .B1(new_n896), .B2(new_n900), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n595), .B(new_n842), .C1(new_n854), .C2(new_n856), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(G162gat), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n903), .A2(new_n904), .A3(new_n899), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n901), .A2(new_n905), .ZN(G1347gat));
  NOR2_X1   g705(.A1(new_n694), .A2(new_n422), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n365), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT123), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n802), .A2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(G169gat), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n910), .A2(new_n911), .A3(new_n272), .ZN(new_n912));
  INV_X1    g711(.A(new_n907), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n801), .A2(new_n808), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(G169gat), .B1(new_n914), .B2(new_n688), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n912), .A2(new_n915), .ZN(G1348gat));
  NAND4_X1  g715(.A1(new_n802), .A2(G176gat), .A3(new_n632), .A4(new_n909), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n917), .A2(KEYINPUT124), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n917), .A2(KEYINPUT124), .ZN(new_n919));
  AOI21_X1  g718(.A(G176gat), .B1(new_n914), .B2(new_n632), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(G1349gat));
  OAI21_X1  g720(.A(new_n293), .B1(new_n910), .B2(new_n556), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n914), .A2(new_n300), .A3(new_n674), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n924), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g724(.A(G190gat), .B1(new_n910), .B2(new_n675), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(KEYINPUT61), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n914), .A2(new_n301), .A3(new_n595), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(G1351gat));
  AOI21_X1  g728(.A(new_n913), .B1(new_n656), .B2(new_n660), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n843), .A2(new_n930), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n931), .A2(G197gat), .A3(new_n813), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT125), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n881), .A2(new_n844), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n934), .B1(new_n801), .B2(new_n846), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(new_n930), .ZN(new_n936));
  OAI21_X1  g735(.A(G197gat), .B1(new_n936), .B2(new_n272), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n933), .A2(new_n937), .ZN(G1352gat));
  NOR3_X1   g737(.A1(new_n931), .A2(G204gat), .A3(new_n687), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT62), .ZN(new_n940));
  OR2_X1    g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g740(.A(G204gat), .B1(new_n936), .B2(new_n687), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n939), .A2(new_n940), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(G1353gat));
  NOR2_X1   g743(.A1(new_n556), .A2(G211gat), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n835), .A2(new_n487), .A3(new_n930), .A4(new_n945), .ZN(new_n946));
  XOR2_X1   g745(.A(new_n946), .B(KEYINPUT126), .Z(new_n947));
  NAND3_X1  g746(.A1(new_n935), .A2(new_n674), .A3(new_n930), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT63), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n948), .A2(new_n949), .A3(G211gat), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n949), .B1(new_n948), .B2(G211gat), .ZN(new_n952));
  OAI21_X1  g751(.A(KEYINPUT127), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(new_n952), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT127), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n954), .A2(new_n955), .A3(new_n950), .A4(new_n947), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n953), .A2(new_n956), .ZN(G1354gat));
  OAI21_X1  g756(.A(G218gat), .B1(new_n936), .B2(new_n675), .ZN(new_n958));
  OR2_X1    g757(.A1(new_n675), .A2(G218gat), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n958), .B1(new_n931), .B2(new_n959), .ZN(G1355gat));
endmodule


