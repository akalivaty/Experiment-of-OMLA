//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 1 1 0 0 1 0 0 1 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 0 0 1 1 1 0 1 1 1 0 1 0 0 0 0 1 1 0 1 0 0 0 1 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:03 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1208, new_n1209, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  AND2_X1   g0009(.A1(G50), .A2(G226), .ZN(new_n210));
  INV_X1    g0010(.A(G58), .ZN(new_n211));
  INV_X1    g0011(.A(G232), .ZN(new_n212));
  INV_X1    g0012(.A(G77), .ZN(new_n213));
  INV_X1    g0013(.A(G244), .ZN(new_n214));
  OAI22_X1  g0014(.A1(new_n211), .A2(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n210), .B(new_n215), .C1(G116), .C2(G270), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G87), .A2(G250), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G97), .A2(G257), .ZN(new_n218));
  XNOR2_X1  g0018(.A(KEYINPUT64), .B(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  OR2_X1    g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND4_X1  g0021(.A1(new_n216), .A2(new_n217), .A3(new_n218), .A4(new_n221), .ZN(new_n222));
  AND2_X1   g0022(.A1(G107), .A2(G264), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n206), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT1), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g0028(.A1(G58), .A2(G68), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G50), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n209), .B(new_n225), .C1(new_n228), .C2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT65), .B(G264), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n237), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(G50), .ZN(new_n250));
  AOI21_X1  g0050(.A(new_n227), .B1(new_n229), .B2(new_n250), .ZN(new_n251));
  NOR2_X1   g0051(.A1(G20), .A2(G33), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n251), .B1(G150), .B2(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT8), .B(G58), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(KEYINPUT68), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT68), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n256), .A2(new_n211), .A3(KEYINPUT8), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(G20), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n253), .B1(new_n258), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(new_n226), .ZN(new_n264));
  INV_X1    g0064(.A(G1), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(G13), .A3(G20), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n262), .A2(new_n264), .B1(new_n250), .B2(new_n267), .ZN(new_n268));
  AND2_X1   g0068(.A1(new_n263), .A2(new_n226), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n265), .A2(G20), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G50), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n268), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g0074(.A(new_n274), .B(KEYINPUT9), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n226), .B1(G33), .B2(G41), .ZN(new_n276));
  INV_X1    g0076(.A(G41), .ZN(new_n277));
  INV_X1    g0077(.A(G45), .ZN(new_n278));
  AOI21_X1  g0078(.A(G1), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(KEYINPUT66), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n265), .B1(G41), .B2(G45), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT66), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n276), .B1(new_n280), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G226), .ZN(new_n285));
  OR2_X1    g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(KEYINPUT3), .A2(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G1698), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G222), .ZN(new_n290));
  NAND2_X1  g0090(.A1(G223), .A2(G1698), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n288), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n292), .B(new_n276), .C1(G77), .C2(new_n288), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n279), .A2(G274), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n285), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  XOR2_X1   g0095(.A(new_n295), .B(KEYINPUT67), .Z(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G190), .ZN(new_n297));
  INV_X1    g0097(.A(G200), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n275), .B(new_n297), .C1(new_n298), .C2(new_n296), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n299), .B(KEYINPUT10), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n296), .A2(G169), .ZN(new_n301));
  INV_X1    g0101(.A(G179), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n301), .B1(new_n302), .B2(new_n296), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n274), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n300), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT74), .ZN(new_n306));
  AND3_X1   g0106(.A1(KEYINPUT73), .A2(G58), .A3(G68), .ZN(new_n307));
  AOI21_X1  g0107(.A(KEYINPUT73), .B1(G58), .B2(G68), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n227), .B1(new_n309), .B2(new_n230), .ZN(new_n310));
  INV_X1    g0110(.A(new_n252), .ZN(new_n311));
  INV_X1    g0111(.A(G159), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n306), .B1(new_n310), .B2(new_n313), .ZN(new_n314));
  AND2_X1   g0114(.A1(KEYINPUT3), .A2(G33), .ZN(new_n315));
  NOR2_X1   g0115(.A1(KEYINPUT3), .A2(G33), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(KEYINPUT7), .B1(new_n317), .B2(new_n227), .ZN(new_n318));
  AND4_X1   g0118(.A1(KEYINPUT7), .A2(new_n286), .A3(new_n227), .A4(new_n287), .ZN(new_n319));
  OAI21_X1  g0119(.A(G68), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n313), .ZN(new_n321));
  NOR3_X1   g0121(.A1(new_n307), .A2(new_n308), .A3(new_n229), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n321), .B(KEYINPUT74), .C1(new_n227), .C2(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n314), .A2(new_n320), .A3(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT16), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n314), .A2(KEYINPUT16), .A3(new_n320), .A4(new_n323), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n326), .A2(new_n264), .A3(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n258), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n272), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n258), .A2(new_n267), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n328), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n288), .B1(G226), .B2(new_n289), .ZN(new_n333));
  NOR2_X1   g0133(.A1(G223), .A2(G1698), .ZN(new_n334));
  INV_X1    g0134(.A(G87), .ZN(new_n335));
  OAI22_X1  g0135(.A1(new_n333), .A2(new_n334), .B1(new_n259), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n276), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n284), .A2(G232), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n337), .A2(new_n294), .A3(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G169), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OR2_X1    g0141(.A1(new_n339), .A2(G179), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n332), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(KEYINPUT75), .A2(KEYINPUT18), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(KEYINPUT75), .A2(KEYINPUT18), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n343), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  AND3_X1   g0148(.A1(new_n328), .A2(new_n330), .A3(new_n331), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n339), .A2(G200), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n337), .A2(G190), .A3(new_n294), .A4(new_n338), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n349), .A2(KEYINPUT17), .A3(new_n350), .A4(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT17), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n328), .A2(new_n330), .A3(new_n331), .A4(new_n351), .ZN(new_n354));
  INV_X1    g0154(.A(new_n350), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n332), .A2(new_n344), .A3(new_n341), .A4(new_n342), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n352), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  XOR2_X1   g0158(.A(KEYINPUT15), .B(G87), .Z(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n260), .ZN(new_n360));
  XNOR2_X1  g0160(.A(new_n360), .B(KEYINPUT69), .ZN(new_n361));
  OAI221_X1 g0161(.A(new_n361), .B1(new_n227), .B2(new_n213), .C1(new_n254), .C2(new_n311), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n362), .A2(new_n264), .B1(new_n213), .B2(new_n267), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n272), .A2(G77), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n289), .A2(G232), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n288), .B(new_n366), .C1(new_n219), .C2(new_n289), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n367), .B(new_n276), .C1(G107), .C2(new_n288), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n284), .A2(G244), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n368), .A2(new_n294), .A3(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(G190), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n365), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n370), .A2(G200), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  NOR4_X1   g0176(.A1(new_n305), .A2(new_n348), .A3(new_n358), .A4(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n261), .A2(new_n213), .ZN(new_n378));
  OAI22_X1  g0178(.A1(new_n311), .A2(new_n250), .B1(new_n227), .B2(G68), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n264), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  XNOR2_X1  g0180(.A(new_n380), .B(KEYINPUT11), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n267), .A2(new_n220), .ZN(new_n382));
  AND2_X1   g0182(.A1(new_n382), .A2(KEYINPUT12), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n382), .A2(KEYINPUT12), .ZN(new_n384));
  OAI221_X1 g0184(.A(new_n381), .B1(new_n220), .B2(new_n271), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  OAI211_X1 g0185(.A(G1), .B(G13), .C1(new_n259), .C2(new_n277), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n279), .A2(KEYINPUT66), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n281), .A2(new_n282), .ZN(new_n388));
  OAI211_X1 g0188(.A(G238), .B(new_n386), .C1(new_n387), .C2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n294), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n212), .A2(G1698), .ZN(new_n391));
  OAI221_X1 g0191(.A(new_n391), .B1(G226), .B2(G1698), .C1(new_n315), .C2(new_n316), .ZN(new_n392));
  NAND2_X1  g0192(.A1(G33), .A2(G97), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n386), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(KEYINPUT13), .B1(new_n390), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n394), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT13), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n396), .A2(new_n397), .A3(new_n294), .A4(new_n389), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n385), .B1(G200), .B2(new_n399), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n399), .A2(new_n371), .ZN(new_n401));
  OR2_X1    g0201(.A1(new_n401), .A2(KEYINPUT70), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(KEYINPUT70), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n400), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n395), .A2(new_n398), .A3(G179), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT71), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n395), .A2(new_n398), .A3(KEYINPUT71), .A4(G179), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT14), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n410), .B1(new_n399), .B2(G169), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  AOI211_X1 g0212(.A(KEYINPUT14), .B(new_n340), .C1(new_n395), .C2(new_n398), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  AND4_X1   g0214(.A1(KEYINPUT72), .A2(new_n409), .A3(new_n412), .A4(new_n414), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n411), .A2(new_n413), .ZN(new_n416));
  AOI21_X1  g0216(.A(KEYINPUT72), .B1(new_n416), .B2(new_n409), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n385), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n370), .A2(new_n340), .ZN(new_n419));
  OR2_X1    g0219(.A1(new_n370), .A2(G179), .ZN(new_n420));
  AND3_X1   g0220(.A1(new_n365), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  AND4_X1   g0222(.A1(new_n377), .A2(new_n404), .A3(new_n418), .A4(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT22), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT83), .ZN(new_n425));
  AOI21_X1  g0225(.A(G20), .B1(new_n286), .B2(new_n287), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n425), .B1(new_n426), .B2(G87), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n227), .B(G87), .C1(new_n315), .C2(new_n316), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n428), .A2(KEYINPUT83), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n424), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(KEYINPUT23), .B1(new_n227), .B2(G107), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT23), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n432), .A2(new_n203), .A3(G20), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n227), .A2(G33), .A3(G116), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n431), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT84), .ZN(new_n436));
  XNOR2_X1  g0236(.A(new_n435), .B(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n426), .A2(new_n425), .A3(G87), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n428), .A2(KEYINPUT83), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n438), .A2(KEYINPUT22), .A3(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n430), .A2(new_n437), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT24), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT24), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n430), .A2(new_n437), .A3(new_n443), .A4(new_n440), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n269), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  XNOR2_X1  g0245(.A(new_n445), .B(KEYINPUT85), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n265), .A2(G33), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n269), .A2(new_n266), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT25), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n450), .B1(new_n266), .B2(G107), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n267), .A2(KEYINPUT25), .A3(new_n203), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n449), .A2(G107), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n288), .B1(G257), .B2(new_n289), .ZN(new_n454));
  NOR2_X1   g0254(.A1(G250), .A2(G1698), .ZN(new_n455));
  INV_X1    g0255(.A(G294), .ZN(new_n456));
  OAI22_X1  g0256(.A1(new_n454), .A2(new_n455), .B1(new_n259), .B2(new_n456), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n278), .A2(G1), .ZN(new_n458));
  XNOR2_X1  g0258(.A(KEYINPUT5), .B(G41), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n276), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  AOI22_X1  g0260(.A1(new_n457), .A2(new_n276), .B1(G264), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n459), .A2(G274), .A3(new_n458), .ZN(new_n462));
  XNOR2_X1  g0262(.A(new_n462), .B(KEYINPUT78), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(new_n298), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n465), .A2(G190), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n446), .A2(new_n453), .A3(new_n467), .A4(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(G33), .A2(G283), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n470), .B(new_n227), .C1(G33), .C2(new_n202), .ZN(new_n471));
  INV_X1    g0271(.A(G116), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(G20), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n471), .A2(new_n264), .A3(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT20), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n471), .A2(KEYINPUT20), .A3(new_n264), .A4(new_n473), .ZN(new_n477));
  AOI22_X1  g0277(.A1(G116), .A2(new_n449), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n266), .A2(G116), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT81), .ZN(new_n480));
  XNOR2_X1  g0280(.A(new_n479), .B(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n340), .B1(new_n478), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n289), .A2(G257), .ZN(new_n483));
  NAND2_X1  g0283(.A1(G264), .A2(G1698), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n483), .B(new_n484), .C1(new_n315), .C2(new_n316), .ZN(new_n485));
  INV_X1    g0285(.A(G303), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n286), .A2(new_n486), .A3(new_n287), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT80), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n386), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n485), .A2(KEYINPUT80), .A3(new_n487), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n460), .A2(G270), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n492), .A2(new_n463), .A3(new_n493), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n482), .A2(KEYINPUT21), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(KEYINPUT21), .B1(new_n482), .B2(new_n494), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n490), .A2(new_n491), .B1(new_n460), .B2(G270), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n269), .A2(G116), .A3(new_n266), .A4(new_n447), .ZN(new_n498));
  INV_X1    g0298(.A(new_n476), .ZN(new_n499));
  INV_X1    g0299(.A(new_n477), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n481), .B(new_n498), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  AND4_X1   g0301(.A1(G179), .A2(new_n497), .A3(new_n501), .A4(new_n463), .ZN(new_n502));
  NOR3_X1   g0302(.A1(new_n495), .A2(new_n496), .A3(new_n502), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n492), .A2(new_n463), .A3(G190), .A4(new_n493), .ZN(new_n504));
  INV_X1    g0304(.A(new_n501), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n298), .B1(new_n497), .B2(new_n463), .ZN(new_n507));
  OAI21_X1  g0307(.A(KEYINPUT82), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n494), .A2(G200), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT82), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n509), .A2(new_n510), .A3(new_n505), .A4(new_n504), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT4), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n513), .A2(G1698), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n514), .B(G244), .C1(new_n316), .C2(new_n315), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n214), .B1(new_n286), .B2(new_n287), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n515), .B(new_n470), .C1(new_n516), .C2(KEYINPUT4), .ZN(new_n517));
  OAI21_X1  g0317(.A(G250), .B1(new_n315), .B2(new_n316), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n289), .B1(new_n518), .B2(KEYINPUT4), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n276), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n460), .A2(G257), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n520), .A2(new_n463), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n340), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n520), .A2(new_n463), .A3(new_n302), .A4(new_n521), .ZN(new_n524));
  AND2_X1   g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT6), .ZN(new_n526));
  AND2_X1   g0326(.A1(G97), .A2(G107), .ZN(new_n527));
  NOR2_X1   g0327(.A1(G97), .A2(G107), .ZN(new_n528));
  OAI211_X1 g0328(.A(KEYINPUT76), .B(new_n526), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n526), .A2(KEYINPUT76), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G97), .A2(G107), .ZN(new_n531));
  NAND2_X1  g0331(.A1(KEYINPUT6), .A2(G107), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n204), .A2(new_n530), .A3(new_n531), .A4(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(G20), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n311), .A2(new_n213), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n535), .A2(KEYINPUT77), .A3(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(G107), .B1(new_n318), .B2(new_n319), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT77), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n227), .B1(new_n529), .B2(new_n533), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n540), .B1(new_n541), .B2(new_n536), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n538), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n264), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n266), .A2(G97), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n448), .A2(new_n202), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n544), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n525), .A2(new_n549), .ZN(new_n550));
  AOI211_X1 g0350(.A(new_n545), .B(new_n547), .C1(new_n543), .C2(new_n264), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n522), .A2(G200), .ZN(new_n552));
  INV_X1    g0352(.A(new_n522), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(G190), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n551), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  AND4_X1   g0355(.A1(new_n503), .A2(new_n512), .A3(new_n550), .A4(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n442), .A2(new_n444), .ZN(new_n557));
  AOI21_X1  g0357(.A(KEYINPUT85), .B1(new_n557), .B2(new_n264), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT85), .ZN(new_n559));
  AOI211_X1 g0359(.A(new_n559), .B(new_n269), .C1(new_n442), .C2(new_n444), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n453), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n464), .A2(G179), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n562), .B1(new_n340), .B2(new_n464), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(G238), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n289), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n214), .A2(G1698), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n566), .B(new_n567), .C1(new_n315), .C2(new_n316), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n259), .A2(new_n472), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n386), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  OR3_X1    g0371(.A1(new_n278), .A2(G1), .A3(G274), .ZN(new_n572));
  INV_X1    g0372(.A(G250), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(new_n278), .B2(G1), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n572), .A2(new_n386), .A3(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(G200), .B1(new_n571), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n528), .A2(new_n335), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n393), .A2(new_n227), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n578), .A2(new_n579), .A3(KEYINPUT19), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n227), .B(G68), .C1(new_n315), .C2(new_n316), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT19), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(new_n393), .B2(G20), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n359), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n584), .A2(new_n264), .B1(new_n267), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n449), .A2(G87), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n577), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(KEYINPUT79), .ZN(new_n589));
  INV_X1    g0389(.A(new_n571), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n590), .A2(G190), .A3(new_n575), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT79), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n577), .A2(new_n586), .A3(new_n592), .A4(new_n587), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n589), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n449), .A2(new_n359), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n586), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n571), .A2(new_n576), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n302), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n340), .B1(new_n571), .B2(new_n576), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n596), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  AND2_X1   g0400(.A1(new_n594), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n469), .A2(new_n556), .A3(new_n564), .A4(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n423), .A2(new_n603), .ZN(G372));
  NAND2_X1  g0404(.A1(new_n352), .A2(new_n356), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n418), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n421), .A2(new_n404), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT88), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n343), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n332), .A2(KEYINPUT88), .A3(new_n341), .A4(new_n342), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n611), .A2(KEYINPUT18), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(KEYINPUT18), .B1(new_n611), .B2(new_n612), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n609), .A2(new_n615), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n616), .A2(new_n300), .B1(new_n274), .B2(new_n303), .ZN(new_n617));
  XNOR2_X1  g0417(.A(new_n617), .B(KEYINPUT89), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n564), .A2(new_n503), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n555), .A2(new_n550), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n591), .A2(new_n577), .A3(new_n586), .A4(new_n587), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n600), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n619), .A2(new_n469), .A3(new_n620), .A4(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n523), .A2(new_n524), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n551), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g0425(.A(KEYINPUT86), .B(KEYINPUT26), .Z(new_n626));
  NAND3_X1  g0426(.A1(new_n601), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n525), .A2(new_n549), .A3(new_n622), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT26), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n600), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(KEYINPUT87), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT87), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n631), .A2(new_n634), .A3(new_n600), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n623), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n423), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n618), .A2(new_n637), .ZN(G369));
  INV_X1    g0438(.A(G13), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n639), .A2(G20), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n226), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT27), .ZN(new_n643));
  NOR3_X1   g0443(.A1(new_n642), .A2(KEYINPUT90), .A3(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(G213), .B1(new_n641), .B2(KEYINPUT27), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT90), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n646), .B1(new_n641), .B2(KEYINPUT27), .ZN(new_n647));
  NOR3_X1   g0447(.A1(new_n644), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(G343), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n561), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n469), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n564), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n561), .A2(new_n563), .A3(new_n649), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  OR3_X1    g0455(.A1(new_n495), .A2(new_n496), .A3(new_n502), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n505), .A2(new_n649), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n503), .A2(new_n512), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n658), .B1(new_n659), .B2(new_n657), .ZN(new_n660));
  XNOR2_X1  g0460(.A(KEYINPUT91), .B(G330), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n655), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n503), .A2(new_n650), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n469), .A2(new_n564), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n654), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n663), .A2(new_n666), .ZN(G399));
  INV_X1    g0467(.A(new_n207), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n668), .A2(G41), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(G1), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n528), .A2(new_n335), .A3(new_n472), .ZN(new_n672));
  OAI22_X1  g0472(.A1(new_n671), .A2(new_n672), .B1(new_n231), .B2(new_n670), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n673), .B(KEYINPUT28), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n634), .B1(new_n631), .B2(new_n600), .ZN(new_n675));
  INV_X1    g0475(.A(new_n600), .ZN(new_n676));
  AOI211_X1 g0476(.A(KEYINPUT87), .B(new_n676), .C1(new_n627), .C2(new_n630), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n650), .B1(new_n678), .B2(new_n623), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n679), .A2(KEYINPUT29), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(KEYINPUT92), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT92), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT94), .ZN(new_n683));
  XOR2_X1   g0483(.A(new_n600), .B(KEYINPUT93), .Z(new_n684));
  AOI21_X1  g0484(.A(new_n626), .B1(new_n601), .B2(new_n625), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n628), .A2(new_n629), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n684), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  OAI211_X1 g0487(.A(new_n453), .B(new_n468), .C1(new_n558), .C2(new_n560), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n620), .B1(new_n688), .B2(new_n466), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n622), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n691), .B1(new_n564), .B2(new_n503), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n687), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n683), .B1(new_n693), .B2(new_n650), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n656), .B1(new_n561), .B2(new_n563), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n689), .A2(new_n695), .A3(new_n691), .ZN(new_n696));
  OAI211_X1 g0496(.A(KEYINPUT94), .B(new_n649), .C1(new_n696), .C2(new_n687), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n682), .B1(new_n698), .B2(KEYINPUT29), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n681), .B1(new_n699), .B2(new_n680), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n494), .A2(new_n302), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n701), .A2(new_n461), .A3(new_n597), .A4(new_n553), .ZN(new_n702));
  XOR2_X1   g0502(.A(new_n702), .B(KEYINPUT30), .Z(new_n703));
  NAND4_X1  g0503(.A1(new_n464), .A2(new_n302), .A3(new_n494), .A4(new_n522), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(new_n597), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n650), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  OAI211_X1 g0506(.A(KEYINPUT31), .B(new_n706), .C1(new_n602), .C2(new_n650), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n706), .A2(KEYINPUT31), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(new_n661), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n700), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n674), .B1(new_n712), .B2(G1), .ZN(G364));
  NAND3_X1  g0513(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(new_n371), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(G326), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n317), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n227), .A2(new_n371), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n298), .A2(G179), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(new_n486), .ZN(new_n722));
  OR3_X1    g0522(.A1(new_n227), .A2(KEYINPUT96), .A3(G190), .ZN(new_n723));
  OAI21_X1  g0523(.A(KEYINPUT96), .B1(new_n227), .B2(G190), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n725), .A2(G179), .A3(G200), .ZN(new_n726));
  XNOR2_X1  g0526(.A(new_n726), .B(KEYINPUT98), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n728), .A2(G329), .ZN(new_n729));
  NOR3_X1   g0529(.A1(new_n725), .A2(G179), .A3(new_n298), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(G283), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n714), .A2(G190), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  OR2_X1    g0535(.A1(KEYINPUT33), .A2(G317), .ZN(new_n736));
  NAND2_X1  g0536(.A1(KEYINPUT33), .A2(G317), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OR4_X1    g0538(.A1(new_n722), .A2(new_n729), .A3(new_n733), .A4(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n302), .A2(G200), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n719), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  AOI211_X1 g0542(.A(new_n718), .B(new_n739), .C1(G322), .C2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n227), .A2(G190), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(new_n740), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G311), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n302), .A2(new_n298), .A3(G190), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G20), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  OAI211_X1 g0550(.A(new_n743), .B(new_n747), .C1(new_n456), .C2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n288), .B1(new_n735), .B2(new_n220), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n750), .A2(new_n202), .ZN(new_n753));
  AOI22_X1  g0553(.A1(new_n746), .A2(G77), .B1(G50), .B2(new_n715), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n754), .B1(new_n211), .B2(new_n741), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n753), .B1(new_n756), .B2(KEYINPUT95), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n730), .A2(G107), .ZN(new_n758));
  OAI211_X1 g0558(.A(new_n757), .B(new_n758), .C1(KEYINPUT95), .C2(new_n756), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n721), .A2(new_n335), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n726), .A2(G159), .ZN(new_n761));
  XNOR2_X1  g0561(.A(KEYINPUT97), .B(KEYINPUT32), .ZN(new_n762));
  XOR2_X1   g0562(.A(new_n761), .B(new_n762), .Z(new_n763));
  OR4_X1    g0563(.A1(new_n752), .A2(new_n759), .A3(new_n760), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n751), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n226), .B1(G20), .B2(new_n340), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n668), .A2(new_n288), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n769), .B1(new_n278), .B2(new_n232), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n770), .B1(new_n245), .B2(new_n278), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n288), .A2(G355), .A3(new_n207), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n771), .B(new_n772), .C1(G116), .C2(new_n207), .ZN(new_n773));
  NOR2_X1   g0573(.A1(G13), .A2(G33), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(G20), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n766), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n773), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n776), .B(KEYINPUT99), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  OR2_X1    g0580(.A1(new_n660), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n671), .B1(G45), .B2(new_n640), .ZN(new_n782));
  NAND4_X1  g0582(.A1(new_n767), .A2(new_n778), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  XOR2_X1   g0583(.A(new_n783), .B(KEYINPUT100), .Z(new_n784));
  INV_X1    g0584(.A(new_n662), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n660), .A2(new_n661), .ZN(new_n786));
  NOR3_X1   g0586(.A1(new_n785), .A2(new_n786), .A3(new_n782), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(G396));
  NAND2_X1  g0589(.A1(new_n421), .A2(new_n649), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n649), .B1(new_n363), .B2(new_n364), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n791), .B1(new_n373), .B2(new_n374), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n790), .B1(new_n792), .B2(new_n421), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n679), .B(new_n794), .ZN(new_n795));
  OR2_X1    g0595(.A1(new_n795), .A2(new_n710), .ZN(new_n796));
  INV_X1    g0596(.A(new_n782), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OR2_X1    g0598(.A1(new_n798), .A2(KEYINPUT104), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n795), .A2(new_n710), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n798), .A2(KEYINPUT104), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n766), .A2(new_n774), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n797), .B1(new_n213), .B2(new_n803), .ZN(new_n804));
  XOR2_X1   g0604(.A(new_n804), .B(KEYINPUT101), .Z(new_n805));
  NOR2_X1   g0605(.A1(new_n794), .A2(new_n775), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n746), .A2(G116), .B1(G283), .B2(new_n734), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(new_n731), .B2(new_n335), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n317), .B1(new_n716), .B2(new_n486), .C1(new_n750), .C2(new_n202), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n808), .B(new_n809), .C1(new_n728), .C2(G311), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n810), .B1(new_n203), .B2(new_n721), .C1(new_n456), .C2(new_n741), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n317), .B1(new_n728), .B2(G132), .ZN(new_n812));
  INV_X1    g0612(.A(new_n721), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n730), .A2(G68), .B1(G50), .B2(new_n813), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT103), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n812), .B(new_n815), .C1(new_n211), .C2(new_n750), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n742), .A2(G143), .B1(G150), .B2(new_n734), .ZN(new_n817));
  INV_X1    g0617(.A(G137), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n817), .B1(new_n818), .B2(new_n716), .C1(new_n312), .C2(new_n745), .ZN(new_n819));
  XNOR2_X1  g0619(.A(KEYINPUT102), .B(KEYINPUT34), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n819), .B(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n811), .B1(new_n816), .B2(new_n821), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n805), .B(new_n806), .C1(new_n766), .C2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n802), .A2(new_n824), .ZN(G384));
  INV_X1    g0625(.A(KEYINPUT38), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT105), .ZN(new_n827));
  AND3_X1   g0627(.A1(new_n332), .A2(new_n827), .A3(new_n648), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n827), .B1(new_n332), .B2(new_n648), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n358), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n831), .B1(new_n832), .B2(new_n347), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n343), .B(new_n834), .C1(new_n828), .C2(new_n829), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n332), .A2(new_n648), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n354), .A2(new_n355), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT37), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n343), .A2(new_n840), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n835), .A2(KEYINPUT37), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n826), .B1(new_n833), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n830), .B1(new_n358), .B2(new_n348), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n835), .A2(KEYINPUT37), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n839), .A2(new_n841), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n844), .B(KEYINPUT38), .C1(new_n845), .C2(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n843), .A2(new_n848), .A3(KEYINPUT39), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT39), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n611), .A2(new_n612), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT18), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n611), .A2(KEYINPUT18), .A3(new_n612), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n854), .A2(new_n606), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n834), .A2(new_n836), .ZN(new_n857));
  OAI21_X1  g0657(.A(KEYINPUT37), .B1(new_n852), .B2(new_n857), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n856), .A2(new_n837), .B1(new_n846), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n848), .B1(new_n859), .B2(KEYINPUT38), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n850), .B1(new_n851), .B2(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n418), .A2(new_n650), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n615), .A2(new_n648), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n385), .A2(new_n650), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n418), .A2(new_n404), .A3(new_n865), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n385), .B(new_n650), .C1(new_n415), .C2(new_n417), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n636), .A2(new_n649), .A3(new_n794), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n869), .B1(new_n870), .B2(new_n790), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n843), .A2(new_n848), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n864), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n863), .A2(new_n873), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n423), .B(new_n681), .C1(new_n699), .C2(new_n680), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n618), .ZN(new_n876));
  XOR2_X1   g0676(.A(new_n874), .B(new_n876), .Z(new_n877));
  AOI21_X1  g0677(.A(new_n793), .B1(new_n866), .B2(new_n867), .ZN(new_n878));
  AND3_X1   g0678(.A1(new_n878), .A2(new_n707), .A3(new_n708), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT40), .B1(new_n879), .B2(new_n872), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT106), .ZN(new_n881));
  NOR3_X1   g0681(.A1(new_n833), .A2(new_n842), .A3(new_n826), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n858), .A2(new_n846), .ZN(new_n883));
  NOR3_X1   g0683(.A1(new_n613), .A2(new_n614), .A3(new_n605), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n883), .B1(new_n884), .B2(new_n836), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n882), .B1(new_n826), .B2(new_n885), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n878), .A2(new_n707), .A3(KEYINPUT40), .A4(new_n708), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n881), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AND4_X1   g0688(.A1(KEYINPUT40), .A2(new_n878), .A3(new_n707), .A4(new_n708), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n889), .A2(new_n860), .A3(KEYINPUT106), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n880), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n423), .A2(new_n709), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n891), .B(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n661), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n877), .B(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n895), .B1(new_n265), .B2(new_n640), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n472), .B1(new_n534), .B2(KEYINPUT35), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n897), .B(new_n228), .C1(KEYINPUT35), .C2(new_n534), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n898), .B(KEYINPUT36), .ZN(new_n899));
  NOR4_X1   g0699(.A1(new_n231), .A2(new_n213), .A3(new_n307), .A4(new_n308), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n220), .A2(G50), .ZN(new_n901));
  OAI211_X1 g0701(.A(G1), .B(new_n639), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n896), .A2(new_n899), .A3(new_n902), .ZN(G367));
  AOI21_X1  g0703(.A(KEYINPUT46), .B1(new_n813), .B2(G116), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(G107), .B2(new_n749), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n813), .A2(KEYINPUT46), .A3(G116), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n905), .B(new_n906), .C1(new_n732), .C2(new_n745), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n288), .B1(new_n726), .B2(G317), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n202), .B2(new_n731), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT110), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n907), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI221_X1 g0711(.A(new_n911), .B1(new_n910), .B2(new_n909), .C1(new_n456), .C2(new_n735), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(G311), .B2(new_n715), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n486), .B2(new_n741), .ZN(new_n914));
  XOR2_X1   g0714(.A(new_n914), .B(KEYINPUT111), .Z(new_n915));
  INV_X1    g0715(.A(new_n726), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n916), .A2(new_n818), .ZN(new_n917));
  AOI22_X1  g0717(.A1(G150), .A2(new_n742), .B1(new_n813), .B2(G58), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n312), .B2(new_n735), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n731), .A2(new_n213), .ZN(new_n920));
  AOI211_X1 g0720(.A(new_n919), .B(new_n920), .C1(G143), .C2(new_n715), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n317), .B1(new_n746), .B2(G50), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n749), .A2(G68), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n915), .B1(new_n917), .B2(new_n924), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n925), .B(KEYINPUT47), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n926), .A2(new_n766), .ZN(new_n927));
  OAI221_X1 g0727(.A(new_n777), .B1(new_n207), .B2(new_n585), .C1(new_n241), .C2(new_n769), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n649), .B1(new_n586), .B2(new_n587), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n676), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n930), .B1(new_n691), .B2(new_n929), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n782), .B(new_n928), .C1(new_n931), .C2(new_n780), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n927), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n620), .B1(new_n551), .B2(new_n649), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n625), .A2(new_n650), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n666), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT45), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n666), .A2(new_n936), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT44), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n939), .B(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(new_n663), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n655), .B1(new_n503), .B2(new_n650), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n665), .A2(KEYINPUT109), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n665), .A2(KEYINPUT109), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n947), .A2(new_n785), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n785), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n712), .B1(new_n943), .B2(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n669), .B(KEYINPUT41), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n265), .B1(new_n640), .B2(G45), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n469), .A2(new_n564), .A3(new_n620), .A4(new_n664), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n957), .A2(KEYINPUT42), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n550), .B1(new_n934), .B2(new_n564), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n649), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n957), .A2(KEYINPUT42), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n958), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n931), .A2(KEYINPUT43), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT107), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n931), .A2(KEYINPUT43), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(KEYINPUT108), .Z(new_n967));
  NAND3_X1  g0767(.A1(new_n962), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n965), .B1(new_n962), .B2(new_n967), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n663), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n972), .A2(new_n936), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n971), .B(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n933), .B1(new_n956), .B2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(G387));
  AOI21_X1  g0777(.A(new_n670), .B1(new_n711), .B2(new_n951), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n711), .B2(new_n951), .ZN(new_n979));
  AOI22_X1  g0779(.A1(G97), .A2(new_n730), .B1(new_n726), .B2(G150), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n721), .A2(new_n213), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(new_n329), .B2(new_n734), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n585), .A2(new_n750), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n741), .A2(new_n250), .B1(new_n745), .B2(new_n220), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n317), .B1(new_n715), .B2(G159), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n980), .A2(new_n982), .A3(new_n985), .A4(new_n986), .ZN(new_n987));
  AOI22_X1  g0787(.A1(new_n742), .A2(G317), .B1(G311), .B2(new_n734), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n486), .B2(new_n745), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(G322), .B2(new_n715), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n990), .B(KEYINPUT48), .Z(new_n991));
  OAI221_X1 g0791(.A(new_n991), .B1(new_n732), .B2(new_n750), .C1(new_n456), .C2(new_n721), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n992), .B(KEYINPUT49), .Z(new_n993));
  OAI221_X1 g0793(.A(new_n317), .B1(new_n731), .B2(new_n472), .C1(new_n717), .C2(new_n916), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n987), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n766), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n254), .A2(G50), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n997), .B(KEYINPUT50), .Z(new_n998));
  NOR2_X1   g0798(.A1(new_n220), .A2(new_n213), .ZN(new_n999));
  NOR4_X1   g0799(.A1(new_n998), .A2(G45), .A3(new_n999), .A4(new_n672), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n768), .B1(new_n237), .B2(new_n278), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n288), .A2(new_n672), .A3(new_n207), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1000), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n207), .A2(G107), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n777), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n797), .B1(new_n655), .B2(new_n779), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n996), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n979), .B(new_n1007), .C1(new_n955), .C2(new_n951), .ZN(G393));
  NAND2_X1  g0808(.A1(new_n936), .A2(new_n776), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n742), .A2(G159), .B1(G150), .B2(new_n715), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n1010), .B(KEYINPUT51), .Z(new_n1011));
  OAI221_X1 g0811(.A(new_n1011), .B1(new_n335), .B2(new_n731), .C1(new_n254), .C2(new_n745), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n750), .A2(new_n213), .ZN(new_n1013));
  AND2_X1   g0813(.A1(new_n726), .A2(G143), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n288), .B1(new_n721), .B2(new_n220), .C1(new_n250), .C2(new_n735), .ZN(new_n1015));
  NOR4_X1   g0815(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .A4(new_n1015), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n742), .A2(G311), .B1(G317), .B2(new_n715), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT52), .Z(new_n1018));
  NAND2_X1  g0818(.A1(new_n813), .A2(G283), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n726), .A2(G322), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1018), .A2(new_n758), .A3(new_n1019), .A4(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n750), .A2(new_n472), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n735), .A2(new_n486), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n317), .B1(new_n745), .B2(new_n456), .ZN(new_n1024));
  NOR4_X1   g0824(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n766), .B1(new_n1016), .B2(new_n1025), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n777), .B1(new_n202), .B2(new_n207), .C1(new_n248), .C2(new_n769), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1009), .A2(new_n782), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n942), .B(new_n972), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n712), .A2(new_n1030), .A3(new_n950), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n943), .B1(new_n711), .B2(new_n951), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1031), .A2(new_n1032), .A3(new_n669), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(KEYINPUT113), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT113), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1031), .A2(new_n1032), .A3(new_n1035), .A4(new_n669), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1029), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1030), .B(KEYINPUT112), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n955), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1037), .A2(new_n1040), .ZN(G390));
  OAI21_X1  g0841(.A(new_n849), .B1(new_n886), .B2(KEYINPUT39), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n774), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n258), .A2(new_n803), .ZN(new_n1044));
  XOR2_X1   g0844(.A(KEYINPUT54), .B(G143), .Z(new_n1045));
  AOI22_X1  g0845(.A1(new_n728), .A2(G125), .B1(new_n746), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n813), .A2(G150), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT117), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT53), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1046), .A2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n288), .B1(new_n731), .B2(new_n250), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT116), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n1051), .A2(new_n1052), .B1(G159), .B2(new_n749), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n715), .A2(G128), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1053), .B(new_n1054), .C1(new_n1052), .C2(new_n1051), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n735), .A2(new_n818), .ZN(new_n1056));
  INV_X1    g0856(.A(G132), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n741), .A2(new_n1057), .ZN(new_n1058));
  NOR4_X1   g0858(.A1(new_n1050), .A2(new_n1055), .A3(new_n1056), .A4(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1013), .B1(new_n728), .B2(G294), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n730), .A2(G68), .B1(G97), .B2(new_n746), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n317), .B1(new_n741), .B2(new_n472), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n760), .B(new_n1062), .C1(G107), .C2(new_n734), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1060), .A2(new_n1061), .A3(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(G283), .B2(new_n715), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n766), .B1(new_n1059), .B2(new_n1065), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1043), .A2(new_n782), .A3(new_n1044), .A4(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT114), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n862), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n790), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n679), .B2(new_n794), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1069), .B1(new_n1071), .B2(new_n869), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n694), .A2(new_n697), .A3(new_n790), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n792), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n422), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1073), .A2(new_n1075), .A3(new_n868), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n885), .A2(new_n826), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n862), .B1(new_n1077), .B2(new_n848), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n1042), .A2(new_n1072), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n709), .A2(G330), .A3(new_n878), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1068), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n871), .A2(new_n862), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1082), .B1(new_n861), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1080), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1084), .A2(KEYINPUT114), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1081), .A2(new_n1086), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n707), .A2(new_n708), .A3(new_n661), .A4(new_n794), .ZN(new_n1088));
  OR2_X1    g0888(.A1(new_n1088), .A2(new_n869), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1082), .B(new_n1089), .C1(new_n861), .C2(new_n1083), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(KEYINPUT115), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT115), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1079), .A2(new_n1092), .A3(new_n1089), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1087), .A2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1067), .B1(new_n1095), .B2(new_n955), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1088), .A2(new_n869), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1080), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1071), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n707), .A2(new_n708), .A3(G330), .A4(new_n794), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n1073), .A2(new_n1075), .B1(new_n869), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n1089), .ZN(new_n1103));
  AND2_X1   g0903(.A1(new_n1100), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n423), .A2(G330), .A3(new_n709), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n875), .A2(new_n618), .A3(new_n1105), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1087), .A2(new_n1094), .A3(new_n1107), .ZN(new_n1108));
  AND2_X1   g0908(.A1(new_n1108), .A2(new_n669), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1107), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1095), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1096), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(G378));
  XOR2_X1   g0913(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n305), .B(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n274), .A2(new_n648), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1116), .B(new_n1117), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1118), .A2(new_n775), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n734), .A2(G97), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n923), .A2(new_n277), .A3(new_n317), .A4(new_n1120), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n981), .B(new_n1121), .C1(new_n728), .C2(G283), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n730), .A2(G58), .ZN(new_n1123));
  XOR2_X1   g0923(.A(new_n1123), .B(KEYINPUT118), .Z(new_n1124));
  NAND2_X1  g0924(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(G116), .B2(new_n715), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n1126), .B1(new_n203), .B2(new_n741), .C1(new_n585), .C2(new_n745), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1127), .B(KEYINPUT58), .ZN(new_n1128));
  AOI21_X1  g0928(.A(G50), .B1(new_n287), .B2(new_n277), .ZN(new_n1129));
  AOI21_X1  g0929(.A(G41), .B1(new_n726), .B2(G124), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n813), .A2(new_n1045), .B1(G132), .B2(new_n734), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n742), .A2(G128), .B1(new_n749), .B2(G150), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n715), .A2(G125), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n746), .A2(G137), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1131), .A2(new_n1132), .A3(new_n1133), .A4(new_n1134), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n259), .B(new_n1130), .C1(new_n1135), .C2(KEYINPUT59), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(G159), .B2(new_n730), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1135), .A2(KEYINPUT59), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1129), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1128), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n766), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n803), .A2(new_n250), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  NOR4_X1   g0944(.A1(new_n1119), .A2(new_n797), .A3(new_n1142), .A4(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n879), .A2(new_n872), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT40), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NOR3_X1   g0948(.A1(new_n886), .A2(new_n881), .A3(new_n887), .ZN(new_n1149));
  AOI21_X1  g0949(.A(KEYINPUT106), .B1(new_n889), .B2(new_n860), .ZN(new_n1150));
  OAI211_X1 g0950(.A(G330), .B(new_n1148), .C1(new_n1149), .C2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1151), .A2(new_n1118), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1118), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(new_n891), .B2(G330), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n874), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1151), .A2(new_n1118), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n891), .A2(G330), .A3(new_n1153), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1156), .A2(new_n1157), .A3(new_n863), .A4(new_n873), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n1155), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1145), .B1(new_n1159), .B2(new_n1039), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1106), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1108), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1162), .A2(KEYINPUT57), .A3(new_n1159), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n669), .ZN(new_n1164));
  AOI21_X1  g0964(.A(KEYINPUT57), .B1(new_n1162), .B2(new_n1159), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1160), .B1(new_n1164), .B2(new_n1165), .ZN(G375));
  NOR2_X1   g0966(.A1(new_n920), .A2(new_n288), .ZN(new_n1167));
  XOR2_X1   g0967(.A(new_n1167), .B(KEYINPUT120), .Z(new_n1168));
  AOI22_X1  g0968(.A1(new_n728), .A2(G303), .B1(G107), .B2(new_n746), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n983), .B1(G116), .B2(new_n734), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(G294), .B2(new_n715), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n1172), .B1(new_n202), .B2(new_n721), .C1(new_n732), .C2(new_n741), .ZN(new_n1173));
  XOR2_X1   g0973(.A(new_n1173), .B(KEYINPUT121), .Z(new_n1174));
  NOR2_X1   g0974(.A1(new_n716), .A2(new_n1057), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1124), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(G150), .B2(new_n746), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n721), .A2(new_n312), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n317), .B(new_n1178), .C1(new_n728), .C2(G128), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1177), .B(new_n1179), .C1(new_n250), .C2(new_n750), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT122), .ZN(new_n1181));
  OR2_X1    g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1045), .A2(new_n734), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n742), .A2(G137), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .A4(new_n1185), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1174), .B1(new_n1175), .B2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n797), .B1(new_n1187), .B2(new_n766), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(new_n775), .B2(new_n868), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(new_n220), .B2(new_n803), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1104), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1190), .B1(new_n1191), .B2(new_n1039), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1193));
  XOR2_X1   g0993(.A(new_n953), .B(KEYINPUT119), .Z(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1110), .A2(new_n1193), .A3(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1192), .A2(new_n1196), .ZN(G381));
  NOR2_X1   g0997(.A1(G375), .A2(G378), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1037), .A2(new_n976), .A3(new_n1040), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1198), .A2(new_n1200), .ZN(new_n1201));
  OR3_X1    g1001(.A1(G393), .A2(G384), .A3(G396), .ZN(new_n1202));
  NOR3_X1   g1002(.A1(new_n1201), .A2(G381), .A3(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT123), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NOR4_X1   g1005(.A1(new_n1201), .A2(KEYINPUT123), .A3(G381), .A4(new_n1202), .ZN(new_n1206));
  OR2_X1    g1006(.A1(new_n1205), .A2(new_n1206), .ZN(G407));
  INV_X1    g1007(.A(G343), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1198), .A2(new_n1208), .ZN(new_n1209));
  OAI211_X1 g1009(.A(G213), .B(new_n1209), .C1(new_n1205), .C2(new_n1206), .ZN(G409));
  NAND2_X1  g1010(.A1(G375), .A2(G378), .ZN(new_n1211));
  INV_X1    g1011(.A(G213), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1212), .A2(G343), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1155), .A2(new_n1158), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(new_n1161), .B2(new_n1108), .ZN(new_n1216));
  AOI21_X1  g1016(.A(KEYINPUT124), .B1(new_n1216), .B2(new_n1195), .ZN(new_n1217));
  AND4_X1   g1017(.A1(KEYINPUT124), .A2(new_n1162), .A3(new_n1159), .A4(new_n1195), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1112), .B(new_n1160), .C1(new_n1217), .C2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1193), .A2(KEYINPUT125), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(KEYINPUT60), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT60), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1193), .A2(KEYINPUT125), .A3(new_n1222), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1221), .A2(new_n669), .A3(new_n1110), .A4(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1224), .A2(G384), .A3(new_n1192), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(G384), .B1(new_n1224), .B2(new_n1192), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1211), .A2(new_n1214), .A3(new_n1219), .A4(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1213), .A2(G2897), .ZN(new_n1230));
  XOR2_X1   g1030(.A(new_n1230), .B(KEYINPUT126), .Z(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1224), .A2(new_n1192), .ZN(new_n1233));
  INV_X1    g1033(.A(G384), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1231), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1235), .A2(new_n1225), .A3(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1232), .A2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1213), .B1(G375), .B2(G378), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1238), .B1(new_n1239), .B2(new_n1219), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT63), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1229), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT61), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(G390), .A2(G387), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(G393), .B(G396), .ZN(new_n1245));
  AND3_X1   g1045(.A1(new_n1244), .A2(new_n1199), .A3(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1245), .B1(new_n1244), .B2(new_n1199), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1239), .A2(KEYINPUT63), .A3(new_n1219), .A4(new_n1228), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1242), .A2(new_n1243), .A3(new_n1248), .A4(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1160), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n670), .B1(new_n1216), .B2(KEYINPUT57), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1165), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1251), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1219), .B(new_n1214), .C1(new_n1254), .C2(new_n1112), .ZN(new_n1255));
  AND2_X1   g1055(.A1(new_n1232), .A2(new_n1237), .ZN(new_n1256));
  AOI21_X1  g1056(.A(KEYINPUT61), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  AND2_X1   g1057(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1229), .A2(new_n1258), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1258), .A2(new_n1260), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1239), .A2(new_n1219), .A3(new_n1228), .A4(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1257), .A2(new_n1259), .A3(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1247), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1244), .A2(new_n1245), .A3(new_n1199), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1263), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1250), .A2(new_n1267), .ZN(G405));
  NAND2_X1  g1068(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1112), .B1(new_n1269), .B2(new_n1160), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1248), .B1(new_n1198), .B2(new_n1270), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1198), .A2(new_n1270), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1266), .A2(new_n1272), .ZN(new_n1273));
  AND3_X1   g1073(.A1(new_n1271), .A2(new_n1273), .A3(new_n1228), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1228), .B1(new_n1271), .B2(new_n1273), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1274), .A2(new_n1275), .ZN(G402));
endmodule


