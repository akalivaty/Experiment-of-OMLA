//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 0 1 0 0 1 0 0 0 1 1 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:09 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n223, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n231, new_n232,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1251, new_n1252, new_n1253, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(G20), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n206), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n209), .B1(new_n212), .B2(new_n213), .C1(KEYINPUT1), .C2(new_n220), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n221), .B1(KEYINPUT1), .B2(new_n220), .ZN(G361));
  XNOR2_X1  g0022(.A(G238), .B(G244), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(G232), .ZN(new_n224));
  XOR2_X1   g0024(.A(KEYINPUT2), .B(G226), .Z(new_n225));
  XNOR2_X1  g0025(.A(new_n224), .B(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(G250), .B(G257), .ZN(new_n227));
  XNOR2_X1  g0027(.A(G264), .B(G270), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n226), .B(new_n229), .ZN(G358));
  NAND2_X1  g0030(.A1(new_n202), .A2(G68), .ZN(new_n231));
  INV_X1    g0031(.A(G68), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(G50), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G58), .B(G77), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G87), .B(G97), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G351));
  NAND2_X1  g0040(.A1(G33), .A2(G41), .ZN(new_n241));
  NAND3_X1  g0041(.A1(new_n241), .A2(G1), .A3(G13), .ZN(new_n242));
  INV_X1    g0042(.A(KEYINPUT66), .ZN(new_n243));
  NOR2_X1   g0043(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g0044(.A(KEYINPUT66), .B1(new_n211), .B2(new_n241), .ZN(new_n245));
  NOR2_X1   g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(G1698), .ZN(new_n248));
  OR2_X1    g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  AOI21_X1  g0050(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G223), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n249), .A2(new_n250), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(G222), .A3(new_n248), .ZN(new_n254));
  INV_X1    g0054(.A(G77), .ZN(new_n255));
  OAI211_X1 g0055(.A(new_n252), .B(new_n254), .C1(new_n255), .C2(new_n253), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT65), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n247), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n258), .B1(new_n257), .B2(new_n256), .ZN(new_n259));
  INV_X1    g0059(.A(G274), .ZN(new_n260));
  AND2_X1   g0060(.A1(KEYINPUT64), .A2(G41), .ZN(new_n261));
  NOR2_X1   g0061(.A1(KEYINPUT64), .A2(G41), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G45), .ZN(new_n264));
  AOI211_X1 g0064(.A(G1), .B(new_n260), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n242), .ZN(new_n266));
  INV_X1    g0066(.A(G41), .ZN(new_n267));
  AOI21_X1  g0067(.A(G1), .B1(new_n267), .B2(new_n264), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n265), .B1(G226), .B2(new_n269), .ZN(new_n270));
  AND2_X1   g0070(.A1(new_n259), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G190), .ZN(new_n272));
  INV_X1    g0072(.A(G33), .ZN(new_n273));
  OAI21_X1  g0073(.A(KEYINPUT68), .B1(new_n273), .B2(G20), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT68), .ZN(new_n275));
  INV_X1    g0075(.A(G20), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n275), .A2(new_n276), .A3(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT8), .B(G58), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n203), .A2(G20), .ZN(new_n281));
  NOR2_X1   g0081(.A1(G20), .A2(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G150), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n280), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n210), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT67), .ZN(new_n288));
  XNOR2_X1  g0088(.A(new_n287), .B(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n285), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G13), .ZN(new_n291));
  NOR3_X1   g0091(.A1(new_n291), .A2(new_n276), .A3(G1), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n290), .B1(new_n202), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT73), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT9), .ZN(new_n295));
  INV_X1    g0095(.A(new_n292), .ZN(new_n296));
  INV_X1    g0096(.A(G1), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G20), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n289), .A2(G50), .A3(new_n296), .A4(new_n298), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n293), .A2(new_n294), .A3(new_n295), .A4(new_n299), .ZN(new_n300));
  OAI221_X1 g0100(.A(new_n299), .B1(G50), .B2(new_n296), .C1(new_n289), .C2(new_n285), .ZN(new_n301));
  NAND2_X1  g0101(.A1(KEYINPUT73), .A2(KEYINPUT9), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n294), .A2(new_n295), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n301), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n300), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n259), .A2(new_n270), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G200), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n272), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(KEYINPUT10), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT10), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n272), .A2(new_n305), .A3(new_n310), .A4(new_n307), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G169), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n306), .A2(new_n313), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n314), .B(new_n301), .C1(G179), .C2(new_n306), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n289), .A2(G77), .A3(new_n296), .A4(new_n298), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT71), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n317), .B(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n279), .ZN(new_n320));
  AOI22_X1  g0120(.A1(new_n320), .A2(new_n282), .B1(G20), .B2(G77), .ZN(new_n321));
  XNOR2_X1  g0121(.A(KEYINPUT15), .B(G87), .ZN(new_n322));
  XNOR2_X1  g0122(.A(new_n322), .B(KEYINPUT70), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n321), .B1(new_n323), .B2(new_n278), .ZN(new_n324));
  INV_X1    g0124(.A(new_n289), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n324), .A2(new_n325), .B1(new_n255), .B2(new_n292), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n319), .A2(new_n326), .ZN(new_n327));
  AND2_X1   g0127(.A1(KEYINPUT3), .A2(G33), .ZN(new_n328));
  NOR2_X1   g0128(.A1(KEYINPUT3), .A2(G33), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n251), .A2(G238), .B1(new_n330), .B2(G107), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n253), .A2(G232), .A3(new_n248), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n246), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n265), .B1(G244), .B2(new_n269), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n313), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n327), .A2(KEYINPUT72), .A3(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G179), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n334), .A2(new_n335), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(KEYINPUT72), .B1(new_n327), .B2(new_n337), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n327), .B1(G200), .B2(new_n336), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n334), .A2(new_n335), .A3(G190), .ZN(new_n346));
  XOR2_X1   g0146(.A(new_n346), .B(KEYINPUT69), .Z(new_n347));
  NAND2_X1  g0147(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n325), .A2(new_n292), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n279), .B1(new_n297), .B2(G20), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n350), .A2(new_n351), .B1(new_n292), .B2(new_n279), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT78), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n249), .A2(new_n354), .A3(new_n250), .ZN(new_n355));
  OAI21_X1  g0155(.A(KEYINPUT78), .B1(new_n328), .B2(new_n329), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n355), .A2(new_n356), .A3(new_n276), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT7), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NOR4_X1   g0159(.A1(new_n328), .A2(new_n329), .A3(new_n358), .A4(G20), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT79), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n362), .A2(new_n363), .A3(G68), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n360), .B1(new_n357), .B2(new_n358), .ZN(new_n365));
  OAI21_X1  g0165(.A(KEYINPUT79), .B1(new_n365), .B2(new_n232), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n282), .A2(G159), .ZN(new_n368));
  XNOR2_X1  g0168(.A(new_n368), .B(KEYINPUT80), .ZN(new_n369));
  INV_X1    g0169(.A(G58), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n370), .A2(new_n232), .ZN(new_n371));
  OAI21_X1  g0171(.A(G20), .B1(new_n371), .B2(new_n201), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n369), .A2(KEYINPUT16), .A3(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n289), .B1(new_n367), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n358), .B1(new_n253), .B2(G20), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n361), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(G68), .ZN(new_n378));
  AND2_X1   g0178(.A1(new_n369), .A2(new_n372), .ZN(new_n379));
  AOI21_X1  g0179(.A(KEYINPUT16), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n353), .B1(new_n375), .B2(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n265), .B1(G232), .B2(new_n269), .ZN(new_n383));
  OR2_X1    g0183(.A1(G223), .A2(G1698), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n253), .B(new_n384), .C1(G226), .C2(new_n248), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(G33), .A2(G87), .ZN(new_n387));
  XNOR2_X1  g0187(.A(new_n387), .B(KEYINPUT81), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n246), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n383), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(G169), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(new_n339), .B2(new_n390), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT18), .B1(new_n382), .B2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n363), .B1(new_n362), .B2(G68), .ZN(new_n395));
  NOR3_X1   g0195(.A1(new_n365), .A2(KEYINPUT79), .A3(new_n232), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n374), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n397), .A2(new_n325), .A3(new_n381), .ZN(new_n398));
  INV_X1    g0198(.A(G200), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n390), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n400), .B1(G190), .B2(new_n390), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n398), .A2(new_n401), .A3(new_n352), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT17), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n398), .A2(new_n352), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT18), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n405), .A2(new_n406), .A3(new_n392), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n382), .A2(KEYINPUT17), .A3(new_n401), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n394), .A2(new_n404), .A3(new_n407), .A4(new_n408), .ZN(new_n409));
  OR3_X1    g0209(.A1(new_n316), .A2(new_n349), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n292), .A2(new_n232), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT12), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n411), .A2(KEYINPUT77), .A3(new_n412), .ZN(new_n413));
  XOR2_X1   g0213(.A(KEYINPUT77), .B(KEYINPUT12), .Z(new_n414));
  OAI21_X1  g0214(.A(new_n413), .B1(new_n411), .B2(new_n414), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n282), .A2(G50), .B1(G20), .B2(new_n232), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n416), .B1(new_n278), .B2(new_n255), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n325), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT11), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n415), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n350), .A2(G68), .A3(new_n298), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n420), .B(new_n421), .C1(new_n419), .C2(new_n418), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT13), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n265), .B1(G238), .B2(new_n269), .ZN(new_n424));
  OAI211_X1 g0224(.A(G226), .B(new_n248), .C1(new_n328), .C2(new_n329), .ZN(new_n425));
  NAND2_X1  g0225(.A1(G33), .A2(G97), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI211_X1 g0227(.A(G232), .B(G1698), .C1(new_n328), .C2(new_n329), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT74), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT74), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n253), .A2(new_n430), .A3(G232), .A4(G1698), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n427), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT75), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n246), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  AOI211_X1 g0234(.A(KEYINPUT75), .B(new_n427), .C1(new_n429), .C2(new_n431), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n423), .B(new_n424), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT76), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n424), .B1(new_n434), .B2(new_n435), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT13), .ZN(new_n440));
  AND2_X1   g0240(.A1(new_n425), .A2(new_n426), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n430), .B1(new_n251), .B2(G232), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n428), .A2(KEYINPUT74), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT75), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n432), .A2(new_n433), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n445), .A2(new_n446), .A3(new_n246), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n447), .A2(KEYINPUT76), .A3(new_n423), .A4(new_n424), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n438), .A2(new_n440), .A3(new_n448), .A4(G179), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n313), .B1(new_n440), .B2(new_n436), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT14), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  AOI211_X1 g0252(.A(KEYINPUT14), .B(new_n313), .C1(new_n440), .C2(new_n436), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n422), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n440), .A2(new_n436), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n422), .B1(new_n455), .B2(G200), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n438), .A2(new_n440), .A3(new_n448), .A4(G190), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n410), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT89), .ZN(new_n462));
  INV_X1    g0262(.A(new_n323), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n463), .A2(new_n296), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(G20), .B1(new_n249), .B2(new_n250), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT19), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n276), .B1(new_n426), .B2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(G87), .ZN(new_n469));
  INV_X1    g0269(.A(G97), .ZN(new_n470));
  INV_X1    g0270(.A(G107), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n466), .A2(G68), .B1(new_n468), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n274), .A2(new_n277), .A3(G97), .ZN(new_n474));
  AND3_X1   g0274(.A1(new_n474), .A2(KEYINPUT87), .A3(new_n467), .ZN(new_n475));
  AOI21_X1  g0275(.A(KEYINPUT87), .B1(new_n474), .B2(new_n467), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n473), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT88), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n289), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  OAI211_X1 g0279(.A(KEYINPUT88), .B(new_n473), .C1(new_n475), .C2(new_n476), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n297), .A2(G33), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n289), .A2(new_n296), .A3(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(G87), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n297), .A2(G45), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n486), .A2(G274), .ZN(new_n487));
  AOI21_X1  g0287(.A(G250), .B1(new_n297), .B2(G45), .ZN(new_n488));
  NOR3_X1   g0288(.A1(new_n266), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  OAI211_X1 g0289(.A(G244), .B(G1698), .C1(new_n328), .C2(new_n329), .ZN(new_n490));
  OAI211_X1 g0290(.A(G238), .B(new_n248), .C1(new_n328), .C2(new_n329), .ZN(new_n491));
  NAND2_X1  g0291(.A1(G33), .A2(G116), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n489), .B1(new_n246), .B2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(G190), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n496), .B1(G200), .B2(new_n494), .ZN(new_n497));
  AND4_X1   g0297(.A1(new_n465), .A2(new_n481), .A3(new_n485), .A4(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n494), .A2(new_n339), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n499), .B1(G169), .B2(new_n494), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n464), .B1(new_n479), .B2(new_n480), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n484), .A2(new_n463), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n462), .B1(new_n498), .B2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT84), .ZN(new_n505));
  OAI211_X1 g0305(.A(G244), .B(new_n248), .C1(new_n328), .C2(new_n329), .ZN(new_n506));
  AOI21_X1  g0306(.A(KEYINPUT4), .B1(new_n506), .B2(KEYINPUT83), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n506), .A2(KEYINPUT83), .A3(KEYINPUT4), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n251), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n505), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AND3_X1   g0312(.A1(new_n506), .A2(KEYINPUT83), .A3(KEYINPUT4), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n505), .B(new_n511), .C1(new_n513), .C2(new_n507), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n246), .B1(new_n512), .B2(new_n515), .ZN(new_n516));
  OR2_X1    g0316(.A1(KEYINPUT64), .A2(G41), .ZN(new_n517));
  NAND2_X1  g0317(.A1(KEYINPUT64), .A2(G41), .ZN(new_n518));
  AOI21_X1  g0318(.A(KEYINPUT5), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT5), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n297), .B(G45), .C1(new_n520), .C2(G41), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n266), .A2(new_n260), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n521), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n520), .B1(new_n261), .B2(new_n262), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n266), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n527), .A2(KEYINPUT85), .A3(G257), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(KEYINPUT85), .B1(new_n527), .B2(G257), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n524), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n516), .A2(G179), .A3(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n511), .B1(new_n513), .B2(new_n507), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(KEYINPUT84), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n247), .B1(new_n535), .B2(new_n514), .ZN(new_n536));
  OAI21_X1  g0336(.A(G169), .B1(new_n536), .B2(new_n531), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n533), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n282), .A2(G77), .ZN(new_n539));
  XOR2_X1   g0339(.A(new_n539), .B(KEYINPUT82), .Z(new_n540));
  INV_X1    g0340(.A(KEYINPUT6), .ZN(new_n541));
  NOR3_X1   g0341(.A1(new_n541), .A2(new_n470), .A3(G107), .ZN(new_n542));
  XNOR2_X1  g0342(.A(G97), .B(G107), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n542), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n540), .B1(new_n276), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n471), .B1(new_n361), .B2(new_n376), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n325), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n484), .A2(G97), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n292), .A2(new_n470), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(KEYINPUT86), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT86), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n547), .A2(new_n552), .A3(new_n548), .A4(new_n549), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n538), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n466), .A2(G68), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n468), .A2(new_n472), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n474), .A2(new_n467), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT87), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n474), .A2(KEYINPUT87), .A3(new_n467), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n558), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n325), .B1(new_n563), .B2(KEYINPUT88), .ZN(new_n564));
  INV_X1    g0364(.A(new_n480), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n502), .B(new_n465), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n500), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n501), .A2(new_n485), .A3(new_n497), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n568), .A2(KEYINPUT89), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n516), .A2(G190), .A3(new_n532), .ZN(new_n571));
  OAI21_X1  g0371(.A(G200), .B1(new_n536), .B2(new_n531), .ZN(new_n572));
  INV_X1    g0372(.A(new_n550), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n504), .A2(new_n555), .A3(new_n570), .A4(new_n574), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n276), .B(G87), .C1(new_n328), .C2(new_n329), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(KEYINPUT22), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT22), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n253), .A2(new_n578), .A3(new_n276), .A4(G87), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT24), .ZN(new_n581));
  OR3_X1    g0381(.A1(new_n492), .A2(KEYINPUT91), .A3(G20), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT23), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(new_n276), .B2(G107), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n471), .A2(KEYINPUT23), .A3(G20), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(KEYINPUT91), .B1(new_n492), .B2(G20), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n582), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n580), .A2(new_n581), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n581), .B1(new_n580), .B2(new_n588), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n325), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n292), .A2(new_n471), .ZN(new_n592));
  XNOR2_X1  g0392(.A(new_n592), .B(KEYINPUT25), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n593), .B1(new_n484), .B2(G107), .ZN(new_n594));
  OAI211_X1 g0394(.A(G264), .B(new_n242), .C1(new_n519), .C2(new_n521), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT92), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n527), .A2(KEYINPUT92), .A3(G264), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n253), .A2(G257), .A3(G1698), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n253), .A2(G250), .A3(new_n248), .ZN(new_n600));
  INV_X1    g0400(.A(G294), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n599), .B(new_n600), .C1(new_n273), .C2(new_n601), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n597), .A2(new_n598), .B1(new_n602), .B2(new_n246), .ZN(new_n603));
  AOI21_X1  g0403(.A(G200), .B1(new_n603), .B2(new_n524), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n602), .A2(new_n246), .ZN(new_n605));
  AND4_X1   g0405(.A1(new_n495), .A2(new_n605), .A3(new_n524), .A4(new_n595), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n591), .B(new_n594), .C1(new_n604), .C2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n597), .A2(new_n598), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n608), .A2(G179), .A3(new_n524), .A4(new_n605), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n605), .A2(new_n524), .A3(new_n595), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n609), .B1(new_n610), .B2(new_n313), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n591), .A2(new_n594), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n607), .A2(new_n613), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n289), .A2(G116), .A3(new_n296), .A4(new_n482), .ZN(new_n615));
  INV_X1    g0415(.A(G116), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n292), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(G20), .B1(G33), .B2(G283), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n273), .A2(G97), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g0420(.A(new_n620), .B(KEYINPUT90), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n286), .A2(new_n210), .B1(G20), .B2(new_n616), .ZN(new_n622));
  AOI21_X1  g0422(.A(KEYINPUT20), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n620), .A2(KEYINPUT90), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT90), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n625), .B1(new_n618), .B2(new_n619), .ZN(new_n626));
  OAI211_X1 g0426(.A(KEYINPUT20), .B(new_n622), .C1(new_n624), .C2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n615), .B(new_n617), .C1(new_n623), .C2(new_n628), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n527), .A2(G270), .B1(new_n522), .B2(new_n523), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n251), .A2(G264), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n253), .A2(G257), .A3(new_n248), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n330), .A2(G303), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n246), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n313), .B1(new_n630), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n629), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT21), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n630), .A2(new_n635), .A3(G179), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n629), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n629), .A2(KEYINPUT21), .A3(new_n636), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n630), .A2(new_n635), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(G200), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n622), .B1(new_n624), .B2(new_n626), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT20), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n648), .A2(new_n627), .B1(new_n616), .B2(new_n292), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n630), .A2(new_n635), .A3(G190), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n645), .A2(new_n615), .A3(new_n649), .A4(new_n650), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n639), .A2(new_n642), .A3(new_n643), .A4(new_n651), .ZN(new_n652));
  NOR4_X1   g0452(.A1(new_n461), .A2(new_n575), .A3(new_n614), .A4(new_n652), .ZN(G372));
  INV_X1    g0453(.A(new_n315), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n394), .A2(new_n407), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n458), .A2(new_n343), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n454), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n404), .A2(new_n408), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n655), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n654), .B1(new_n659), .B2(new_n312), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n607), .A2(new_n569), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n613), .A2(new_n639), .A3(new_n642), .A4(new_n643), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n555), .A2(new_n661), .A3(new_n662), .A4(new_n574), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n494), .A2(G169), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(KEYINPUT93), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT93), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n666), .B1(new_n494), .B2(G169), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n566), .A2(new_n499), .A3(new_n665), .A4(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n663), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT26), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n538), .A2(KEYINPUT94), .A3(new_n550), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n671), .A2(new_n569), .A3(new_n668), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n573), .B1(new_n533), .B2(new_n537), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n673), .A2(KEYINPUT94), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n670), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  AND3_X1   g0475(.A1(new_n568), .A2(KEYINPUT89), .A3(new_n569), .ZN(new_n676));
  AOI21_X1  g0476(.A(KEYINPUT89), .B1(new_n568), .B2(new_n569), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n555), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(KEYINPUT26), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n669), .B1(new_n675), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n660), .B1(new_n461), .B2(new_n681), .ZN(G369));
  NAND3_X1  g0482(.A1(new_n297), .A2(new_n276), .A3(G13), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(KEYINPUT27), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT95), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n684), .B(new_n685), .ZN(new_n686));
  OAI211_X1 g0486(.A(new_n686), .B(G213), .C1(KEYINPUT27), .C2(new_n683), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT96), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n687), .A2(new_n688), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(G343), .A3(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(new_n612), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n693), .A2(new_n613), .A3(new_n607), .ZN(new_n694));
  INV_X1    g0494(.A(new_n613), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n692), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n639), .A2(new_n642), .A3(new_n643), .ZN(new_n698));
  INV_X1    g0498(.A(new_n629), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n691), .A2(new_n699), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n652), .A2(new_n700), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AND3_X1   g0503(.A1(new_n703), .A2(KEYINPUT97), .A3(G330), .ZN(new_n704));
  AOI21_X1  g0504(.A(KEYINPUT97), .B1(new_n703), .B2(G330), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n697), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n698), .A2(new_n691), .ZN(new_n708));
  OR2_X1    g0508(.A1(new_n708), .A2(new_n614), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n613), .B2(new_n692), .ZN(new_n710));
  OR2_X1    g0510(.A1(new_n707), .A2(new_n710), .ZN(G399));
  NAND2_X1  g0511(.A1(new_n263), .A2(new_n207), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n472), .A2(G116), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n712), .A2(G1), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(new_n213), .B2(new_n712), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n715), .B(KEYINPUT28), .ZN(new_n716));
  NOR3_X1   g0516(.A1(new_n681), .A2(KEYINPUT29), .A3(new_n692), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT29), .ZN(new_n718));
  INV_X1    g0518(.A(new_n669), .ZN(new_n719));
  OAI21_X1  g0519(.A(KEYINPUT26), .B1(new_n672), .B2(new_n674), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n678), .A2(new_n670), .A3(new_n679), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n719), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n718), .B1(new_n722), .B2(new_n691), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n717), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n652), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n725), .A2(new_n613), .A3(new_n607), .A4(new_n691), .ZN(new_n726));
  OAI21_X1  g0526(.A(KEYINPUT98), .B1(new_n575), .B2(new_n726), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n614), .A2(new_n652), .A3(new_n692), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT98), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n516), .A2(new_n532), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n550), .B1(new_n730), .B2(G200), .ZN(new_n731));
  AOI22_X1  g0531(.A1(new_n571), .A2(new_n731), .B1(new_n538), .B2(new_n554), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n678), .A2(new_n728), .A3(new_n729), .A4(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n727), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n608), .A2(new_n494), .A3(new_n605), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(new_n640), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n736), .A2(new_n516), .A3(new_n532), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT30), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n603), .A2(new_n524), .ZN(new_n740));
  AOI211_X1 g0540(.A(G179), .B(new_n494), .C1(new_n635), .C2(new_n630), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n730), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n736), .A2(new_n516), .A3(KEYINPUT30), .A4(new_n532), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n739), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(new_n692), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT31), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n744), .A2(KEYINPUT31), .A3(new_n692), .ZN(new_n748));
  AND2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n734), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G330), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n724), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n716), .B1(new_n753), .B2(G1), .ZN(G364));
  NOR2_X1   g0554(.A1(new_n704), .A2(new_n705), .ZN(new_n755));
  INV_X1    g0555(.A(new_n712), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n291), .A2(G20), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n297), .B1(new_n757), .B2(G45), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  OAI211_X1 g0561(.A(new_n755), .B(new_n761), .C1(G330), .C2(new_n703), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n210), .B1(G20), .B2(new_n313), .ZN(new_n763));
  OR2_X1    g0563(.A1(new_n763), .A2(KEYINPUT100), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(KEYINPUT100), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n276), .A2(G179), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G190), .A2(G200), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G159), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n767), .A2(new_n495), .A3(G200), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n771), .A2(KEYINPUT32), .B1(G107), .B2(new_n773), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n495), .A2(G179), .A3(G200), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n276), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G97), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n276), .A2(new_n339), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G200), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n495), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n774), .B(new_n778), .C1(new_n202), .C2(new_n782), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n767), .A2(G190), .A3(G200), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G87), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n780), .A2(G190), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n786), .B1(new_n771), .B2(KEYINPUT32), .C1(new_n788), .C2(new_n232), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n779), .A2(new_n768), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n779), .A2(G190), .A3(new_n399), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n253), .B1(new_n790), .B2(new_n255), .C1(new_n370), .C2(new_n791), .ZN(new_n792));
  NOR3_X1   g0592(.A1(new_n783), .A2(new_n789), .A3(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G317), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(KEYINPUT33), .ZN(new_n795));
  OR2_X1    g0595(.A1(new_n794), .A2(KEYINPUT33), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n787), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(G303), .ZN(new_n798));
  INV_X1    g0598(.A(G326), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n797), .B1(new_n798), .B2(new_n784), .C1(new_n799), .C2(new_n782), .ZN(new_n800));
  INV_X1    g0600(.A(new_n791), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n801), .A2(G322), .B1(new_n770), .B2(G329), .ZN(new_n802));
  INV_X1    g0602(.A(G311), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n802), .B(new_n330), .C1(new_n803), .C2(new_n790), .ZN(new_n804));
  INV_X1    g0604(.A(G283), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n776), .A2(new_n601), .B1(new_n772), .B2(new_n805), .ZN(new_n806));
  NOR3_X1   g0606(.A1(new_n800), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n766), .B1(new_n793), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n355), .A2(new_n356), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(new_n207), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT99), .ZN(new_n812));
  INV_X1    g0612(.A(new_n213), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(new_n264), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n812), .B(new_n814), .C1(new_n264), .C2(new_n236), .ZN(new_n815));
  INV_X1    g0615(.A(new_n207), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(new_n330), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n817), .A2(G355), .B1(new_n616), .B2(new_n816), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(G13), .A2(G33), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(G20), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n766), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n808), .B(new_n760), .C1(new_n819), .C2(new_n824), .ZN(new_n825));
  XOR2_X1   g0625(.A(new_n825), .B(KEYINPUT101), .Z(new_n826));
  INV_X1    g0626(.A(new_n822), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n826), .B1(new_n703), .B2(new_n827), .ZN(new_n828));
  AND2_X1   g0628(.A1(new_n762), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(G396));
  NOR2_X1   g0630(.A1(new_n766), .A2(new_n820), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n761), .B1(new_n831), .B2(new_n255), .ZN(new_n832));
  INV_X1    g0632(.A(new_n790), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n781), .A2(G303), .B1(new_n833), .B2(G116), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(new_n805), .B2(new_n788), .ZN(new_n835));
  XOR2_X1   g0635(.A(new_n835), .B(KEYINPUT102), .Z(new_n836));
  OAI221_X1 g0636(.A(new_n330), .B1(new_n769), .B2(new_n803), .C1(new_n791), .C2(new_n601), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n778), .B1(new_n469), .B2(new_n772), .C1(new_n471), .C2(new_n784), .ZN(new_n838));
  NOR3_X1   g0638(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n773), .A2(G68), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n840), .B1(new_n202), .B2(new_n784), .C1(new_n370), .C2(new_n776), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n810), .B(new_n841), .C1(G132), .C2(new_n770), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(KEYINPUT103), .ZN(new_n843));
  OR2_X1    g0643(.A1(new_n842), .A2(KEYINPUT103), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n801), .A2(G143), .B1(new_n833), .B2(G159), .ZN(new_n845));
  INV_X1    g0645(.A(G150), .ZN(new_n846));
  INV_X1    g0646(.A(G137), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n845), .B1(new_n788), .B2(new_n846), .C1(new_n847), .C2(new_n782), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT34), .ZN(new_n849));
  AND2_X1   g0649(.A1(new_n844), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n839), .B1(new_n843), .B2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n766), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n692), .A2(new_n327), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n348), .B(new_n853), .C1(new_n341), .C2(new_n342), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n691), .B1(new_n319), .B2(new_n326), .ZN(new_n855));
  INV_X1    g0655(.A(new_n342), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n855), .A2(new_n856), .A3(new_n340), .A4(new_n338), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  OAI221_X1 g0658(.A(new_n832), .B1(new_n851), .B2(new_n852), .C1(new_n858), .C2(new_n821), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT104), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  AND2_X1   g0661(.A1(new_n854), .A2(new_n857), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n681), .B2(new_n692), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n668), .A2(new_n569), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n864), .B1(KEYINPUT94), .B2(new_n673), .ZN(new_n865));
  INV_X1    g0665(.A(new_n674), .ZN(new_n866));
  AOI21_X1  g0666(.A(KEYINPUT26), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NOR4_X1   g0667(.A1(new_n676), .A2(new_n555), .A3(new_n677), .A4(new_n670), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n719), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n869), .A2(new_n691), .A3(new_n858), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n863), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n751), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n761), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n871), .A2(new_n751), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n861), .B1(new_n873), .B2(new_n874), .ZN(G384));
  NOR2_X1   g0675(.A1(new_n757), .A2(new_n297), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n747), .A2(new_n748), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n877), .B1(new_n733), .B2(new_n727), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT106), .ZN(new_n879));
  AND3_X1   g0679(.A1(new_n692), .A2(new_n879), .A3(new_n422), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n879), .B1(new_n692), .B2(new_n422), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n459), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n454), .A2(new_n458), .A3(new_n882), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n884), .A2(new_n858), .A3(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n878), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n379), .B1(new_n395), .B2(new_n396), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT16), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n353), .B1(new_n890), .B2(new_n375), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n402), .B1(new_n891), .B2(new_n393), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n689), .A2(new_n690), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(KEYINPUT37), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n405), .A2(new_n392), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT37), .ZN(new_n897));
  INV_X1    g0697(.A(new_n893), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n373), .B1(new_n364), .B2(new_n366), .ZN(new_n899));
  NOR3_X1   g0699(.A1(new_n899), .A2(new_n380), .A3(new_n289), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n898), .B1(new_n900), .B2(new_n353), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n896), .A2(new_n897), .A3(new_n901), .A4(new_n402), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n895), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n409), .A2(new_n894), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n903), .A2(new_n904), .A3(KEYINPUT38), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT38), .B1(new_n903), .B2(new_n904), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT107), .ZN(new_n907));
  NOR3_X1   g0707(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n903), .A2(new_n904), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT38), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n903), .A2(new_n904), .A3(KEYINPUT38), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT107), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n887), .B1(new_n908), .B2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT40), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n896), .A2(new_n402), .A3(new_n901), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(KEYINPUT37), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n902), .ZN(new_n919));
  INV_X1    g0719(.A(new_n901), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n409), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n910), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n915), .B1(new_n923), .B2(new_n912), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n887), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n916), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n461), .A2(new_n878), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(G330), .B1(new_n926), .B2(new_n927), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT109), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n931), .B1(new_n930), .B2(new_n929), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT110), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n460), .B1(new_n717), .B2(new_n723), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n660), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT108), .ZN(new_n936));
  AND3_X1   g0736(.A1(new_n454), .A2(new_n458), .A3(new_n882), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n882), .B1(new_n454), .B2(new_n458), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n344), .A2(new_n692), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n940), .B1(new_n870), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n913), .B2(new_n908), .ZN(new_n944));
  AOI21_X1  g0744(.A(KEYINPUT39), .B1(new_n923), .B2(new_n912), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n454), .A2(new_n692), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n911), .A2(KEYINPUT39), .A3(new_n912), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n946), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n655), .A2(new_n898), .ZN(new_n951));
  AND3_X1   g0751(.A1(new_n944), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n936), .B(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n876), .B1(new_n933), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n933), .B2(new_n953), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT35), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n544), .A2(new_n956), .ZN(new_n957));
  AOI211_X1 g0757(.A(new_n616), .B(new_n212), .C1(new_n544), .C2(new_n956), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n957), .B1(new_n959), .B2(KEYINPUT105), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(KEYINPUT105), .B2(new_n959), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT36), .ZN(new_n962));
  OAI21_X1  g0762(.A(G77), .B1(new_n370), .B2(new_n232), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n231), .B1(new_n963), .B2(new_n213), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n964), .A2(G1), .A3(new_n291), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n955), .A2(new_n962), .A3(new_n965), .ZN(G367));
  OAI21_X1  g0766(.A(new_n823), .B1(new_n207), .B2(new_n323), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(new_n812), .B2(new_n229), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n968), .A2(new_n761), .ZN(new_n969));
  OAI22_X1  g0769(.A1(new_n782), .A2(new_n803), .B1(new_n471), .B2(new_n776), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(G294), .B2(new_n787), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n791), .A2(new_n798), .B1(new_n790), .B2(new_n805), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n972), .B1(G317), .B2(new_n770), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n809), .B1(G97), .B2(new_n773), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n971), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n784), .A2(new_n616), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT46), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n772), .A2(new_n255), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(G159), .B2(new_n787), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n370), .B2(new_n784), .ZN(new_n980));
  AOI22_X1  g0780(.A1(G68), .A2(new_n777), .B1(new_n781), .B2(G143), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n330), .B1(new_n770), .B2(G137), .ZN(new_n982));
  AOI22_X1  g0782(.A1(new_n801), .A2(G150), .B1(new_n833), .B2(G50), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n981), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n975), .A2(new_n977), .B1(new_n980), .B2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT47), .ZN(new_n986));
  AND2_X1   g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n766), .B1(new_n985), .B2(new_n986), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n501), .A2(new_n485), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n692), .A2(new_n989), .ZN(new_n990));
  MUX2_X1   g0790(.A(new_n668), .B(new_n864), .S(new_n990), .Z(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n969), .B1(new_n987), .B2(new_n988), .C1(new_n992), .C2(new_n827), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n732), .B1(new_n573), .B2(new_n691), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n673), .A2(new_n692), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT111), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n695), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n692), .B1(new_n998), .B2(new_n555), .ZN(new_n999));
  AND2_X1   g0799(.A1(new_n994), .A2(new_n995), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n1000), .A2(new_n709), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n1001), .B(KEYINPUT42), .Z(new_n1002));
  OR4_X1    g0802(.A1(KEYINPUT43), .A2(new_n999), .A3(new_n1002), .A4(new_n992), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n999), .A2(new_n1002), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT112), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n991), .B(KEYINPUT43), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1003), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1005), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n997), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n1008), .A2(new_n1009), .B1(new_n706), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1009), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1010), .A2(new_n706), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1012), .A2(new_n1013), .A3(new_n1003), .A4(new_n1007), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1011), .A2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1000), .A2(new_n710), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT45), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n707), .A2(KEYINPUT113), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1000), .A2(new_n710), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT44), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1019), .B(new_n1020), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1017), .A2(new_n1018), .A3(new_n1021), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n707), .A2(KEYINPUT113), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1022), .B(new_n1023), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n694), .A2(new_n696), .A3(new_n708), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n709), .A2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n755), .B(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n753), .B1(new_n1024), .B2(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n712), .B(KEYINPUT41), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n759), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n993), .B1(new_n1015), .B2(new_n1031), .ZN(G387));
  NAND2_X1  g0832(.A1(new_n752), .A2(new_n1027), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n1034), .A2(KEYINPUT116), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n752), .A2(new_n1027), .ZN(new_n1036));
  OR3_X1    g0836(.A1(new_n1036), .A2(KEYINPUT115), .A3(new_n712), .ZN(new_n1037));
  OAI21_X1  g0837(.A(KEYINPUT115), .B1(new_n1036), .B2(new_n712), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1034), .A2(KEYINPUT116), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1035), .A2(new_n1037), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1027), .A2(new_n758), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n694), .A2(new_n696), .A3(new_n822), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n817), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n1043), .A2(new_n713), .B1(G107), .B2(new_n207), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n812), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(G45), .B2(new_n226), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n713), .B(new_n264), .C1(new_n232), .C2(new_n255), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT114), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1050));
  OAI21_X1  g0850(.A(KEYINPUT50), .B1(new_n279), .B2(G50), .ZN(new_n1051));
  OR3_X1    g0851(.A1(new_n279), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1044), .B1(new_n1046), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n760), .B1(new_n1054), .B2(new_n824), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n801), .A2(G317), .B1(new_n833), .B2(G303), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n781), .A2(G322), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1056), .B(new_n1057), .C1(new_n803), .C2(new_n788), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT48), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1060), .B1(new_n805), .B2(new_n776), .C1(new_n601), .C2(new_n784), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  AND2_X1   g0863(.A1(new_n1063), .A2(KEYINPUT49), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n810), .B1(new_n616), .B2(new_n772), .C1(new_n799), .C2(new_n769), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(KEYINPUT49), .B2(new_n1063), .ZN(new_n1067));
  INV_X1    g0867(.A(G159), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n1068), .A2(new_n782), .B1(new_n788), .B2(new_n279), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(G77), .B2(new_n785), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n810), .B1(G97), .B2(new_n773), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n463), .A2(new_n777), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n791), .A2(new_n202), .B1(new_n790), .B2(new_n232), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(G150), .B2(new_n770), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1070), .A2(new_n1071), .A3(new_n1072), .A4(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1067), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1055), .B1(new_n1076), .B2(new_n766), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1041), .B1(new_n1042), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1040), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(KEYINPUT117), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT117), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1040), .A2(new_n1081), .A3(new_n1078), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1080), .A2(new_n1082), .ZN(G393));
  INV_X1    g0883(.A(new_n1024), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n712), .B1(new_n1084), .B2(new_n1036), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n1036), .B2(new_n1084), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1010), .A2(new_n822), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n823), .B1(new_n470), .B2(new_n207), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(new_n812), .B2(new_n239), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n782), .A2(new_n794), .B1(new_n803), .B2(new_n791), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT52), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n790), .A2(new_n601), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n253), .B(new_n1092), .C1(G322), .C2(new_n770), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n787), .A2(G303), .B1(new_n773), .B2(G107), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n777), .A2(G116), .B1(new_n785), .B2(G283), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n1091), .A2(new_n1093), .A3(new_n1094), .A4(new_n1095), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n785), .A2(G68), .B1(new_n773), .B2(G87), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n810), .B(new_n1098), .C1(G143), .C2(new_n770), .ZN(new_n1099));
  OR2_X1    g0899(.A1(new_n1099), .A2(KEYINPUT118), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(KEYINPUT118), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n782), .A2(new_n846), .B1(new_n1068), .B2(new_n791), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT51), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1100), .A2(new_n1101), .A3(new_n1103), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n776), .A2(new_n255), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n320), .B2(new_n833), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1106), .B1(new_n202), .B2(new_n788), .ZN(new_n1107));
  XOR2_X1   g0907(.A(new_n1107), .B(KEYINPUT119), .Z(new_n1108));
  OAI21_X1  g0908(.A(new_n1096), .B1(new_n1104), .B2(new_n1108), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n761), .B(new_n1089), .C1(new_n1109), .C2(new_n766), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n1084), .A2(new_n759), .B1(new_n1087), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1086), .A2(new_n1111), .ZN(G390));
  NOR3_X1   g0912(.A1(new_n751), .A2(new_n862), .A3(new_n940), .ZN(new_n1113));
  NOR3_X1   g0913(.A1(new_n681), .A2(new_n692), .A3(new_n862), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n939), .B1(new_n1114), .B2(new_n941), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n1115), .A2(new_n947), .B1(new_n946), .B2(new_n949), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n722), .A2(new_n691), .A3(new_n858), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n940), .B1(new_n1117), .B2(new_n942), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(new_n947), .B(KEYINPUT120), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n923), .A2(new_n912), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1118), .A2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1113), .B1(new_n1116), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n949), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n943), .A2(new_n948), .B1(new_n1124), .B2(new_n945), .ZN(new_n1125));
  INV_X1    g0925(.A(G330), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n878), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1127), .A2(new_n858), .A3(new_n939), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1125), .B(new_n1128), .C1(new_n1118), .C2(new_n1121), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1123), .A2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1130), .A2(new_n758), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n820), .B1(new_n1124), .B2(new_n945), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n788), .A2(new_n471), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n1105), .B(new_n1133), .C1(G283), .C2(new_n781), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n790), .A2(new_n470), .B1(new_n769), .B2(new_n601), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n253), .B(new_n1135), .C1(G116), .C2(new_n801), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1134), .A2(new_n786), .A3(new_n840), .A4(new_n1136), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n784), .A2(new_n846), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(KEYINPUT121), .B(KEYINPUT53), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1138), .B(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(G132), .ZN(new_n1141));
  INV_X1    g0941(.A(G125), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n791), .A2(new_n1141), .B1(new_n769), .B2(new_n1142), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(KEYINPUT54), .B(G143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n253), .B1(new_n790), .B2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n781), .A2(G128), .B1(new_n773), .B2(G50), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(G159), .A2(new_n777), .B1(new_n787), .B2(G137), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1140), .A2(new_n1146), .A3(new_n1147), .A4(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n852), .B1(new_n1137), .B2(new_n1149), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n761), .B(new_n1150), .C1(new_n279), .C2(new_n831), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1131), .B1(new_n1132), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1127), .A2(new_n460), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n934), .A2(new_n660), .A3(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n870), .A2(new_n942), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n939), .B1(new_n1127), .B2(new_n858), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1155), .B1(new_n1113), .B2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n940), .B1(new_n751), .B2(new_n862), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1158), .A2(new_n1128), .A3(new_n942), .A4(new_n1117), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1154), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1130), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1160), .A2(new_n1123), .A3(new_n1129), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1162), .A2(new_n756), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1152), .A2(new_n1164), .ZN(G378));
  NAND3_X1  g0965(.A1(new_n944), .A2(new_n950), .A3(new_n951), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n898), .A2(new_n301), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n316), .B(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1168), .B(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1126), .B1(new_n924), .B2(new_n887), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1170), .B1(new_n916), .B2(new_n1171), .ZN(new_n1172));
  NOR3_X1   g0972(.A1(new_n937), .A2(new_n938), .A3(new_n862), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n750), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n907), .B1(new_n905), .B2(new_n906), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n911), .A2(KEYINPUT107), .A3(new_n912), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1174), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1171), .B(new_n1170), .C1(new_n1177), .C2(KEYINPUT40), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1166), .B1(new_n1172), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1170), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1177), .A2(KEYINPUT40), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1171), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1181), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1184), .A2(new_n952), .A3(new_n1178), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1180), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1181), .A2(new_n820), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n810), .A2(new_n263), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1188), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n772), .A2(new_n370), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n784), .A2(new_n255), .B1(new_n769), .B2(new_n805), .ZN(new_n1191));
  NOR3_X1   g0991(.A1(new_n1188), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1192), .B(KEYINPUT122), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(G97), .A2(new_n787), .B1(new_n781), .B2(G116), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n777), .A2(G68), .B1(new_n801), .B2(G107), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1194), .B(new_n1195), .C1(new_n323), .C2(new_n790), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1193), .A2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1189), .B1(new_n1197), .B2(KEYINPUT58), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT123), .ZN(new_n1199));
  OR2_X1    g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n1142), .A2(new_n782), .B1(new_n788), .B2(new_n1141), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(G150), .B2(new_n777), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n801), .A2(G128), .B1(new_n833), .B2(G137), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1203), .B(new_n1204), .C1(new_n784), .C2(new_n1144), .ZN(new_n1205));
  OR2_X1    g1005(.A1(new_n1205), .A2(KEYINPUT59), .ZN(new_n1206));
  AOI211_X1 g1006(.A(G33), .B(G41), .C1(new_n770), .C2(G124), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n1068), .B2(new_n772), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(new_n1205), .B2(KEYINPUT59), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n1206), .A2(new_n1209), .B1(KEYINPUT58), .B2(new_n1197), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1200), .A2(new_n1201), .A3(new_n1210), .ZN(new_n1211));
  AND2_X1   g1011(.A1(new_n1211), .A2(new_n766), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n761), .B(new_n1212), .C1(new_n202), .C2(new_n831), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n1186), .A2(new_n759), .B1(new_n1187), .B2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1154), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1163), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(new_n1186), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT57), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1218), .B1(new_n1180), .B2(new_n1185), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n712), .B1(new_n1220), .B2(new_n1216), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT124), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1219), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  AOI211_X1 g1023(.A(KEYINPUT124), .B(new_n712), .C1(new_n1220), .C2(new_n1216), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1214), .B1(new_n1223), .B2(new_n1224), .ZN(G375));
  NAND3_X1  g1025(.A1(new_n1157), .A2(new_n1159), .A3(new_n1154), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1161), .A2(new_n1030), .A3(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n759), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n761), .B1(new_n831), .B2(new_n232), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n781), .A2(G132), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(new_n1231), .B(KEYINPUT125), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(G150), .A2(new_n833), .B1(new_n770), .B2(G128), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1233), .B1(new_n847), .B2(new_n791), .ZN(new_n1234));
  NOR4_X1   g1034(.A1(new_n1232), .A2(new_n810), .A3(new_n1234), .A4(new_n1190), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n788), .A2(new_n1144), .B1(new_n1068), .B2(new_n784), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(G50), .B2(new_n777), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n782), .A2(new_n601), .B1(new_n784), .B2(new_n470), .ZN(new_n1238));
  AOI211_X1 g1038(.A(new_n978), .B(new_n1238), .C1(G116), .C2(new_n787), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n330), .B1(new_n769), .B2(new_n798), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n791), .A2(new_n805), .B1(new_n790), .B2(new_n471), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n1240), .B(new_n1241), .C1(new_n463), .C2(new_n777), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n1235), .A2(new_n1237), .B1(new_n1239), .B2(new_n1242), .ZN(new_n1243));
  OAI221_X1 g1043(.A(new_n1230), .B1(new_n852), .B2(new_n1243), .C1(new_n939), .C2(new_n821), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1227), .A2(new_n1229), .A3(new_n1244), .ZN(G381));
  INV_X1    g1045(.A(G375), .ZN(new_n1246));
  NOR4_X1   g1046(.A1(G387), .A2(G390), .A3(G384), .A4(G381), .ZN(new_n1247));
  INV_X1    g1047(.A(G378), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(G393), .A2(G396), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1246), .A2(new_n1247), .A3(new_n1248), .A4(new_n1249), .ZN(G407));
  INV_X1    g1050(.A(G213), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1251), .A2(G343), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1246), .A2(new_n1248), .A3(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(G407), .A2(G213), .A3(new_n1253), .ZN(G409));
  NAND3_X1  g1054(.A1(G387), .A2(new_n1086), .A3(new_n1111), .ZN(new_n1255));
  OAI211_X1 g1055(.A(G390), .B(new_n993), .C1(new_n1031), .C2(new_n1015), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n829), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1257), .B1(new_n1249), .B2(new_n1258), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1249), .A2(new_n1258), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1260), .A2(new_n1256), .A3(new_n1255), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT61), .ZN(new_n1262));
  AND3_X1   g1062(.A1(new_n1259), .A2(new_n1261), .A3(new_n1262), .ZN(new_n1263));
  OAI211_X1 g1063(.A(G378), .B(new_n1214), .C1(new_n1223), .C2(new_n1224), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1214), .B1(new_n1029), .B2(new_n1217), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1248), .A2(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1252), .B1(new_n1264), .B2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1229), .A2(new_n1244), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT60), .ZN(new_n1269));
  NOR3_X1   g1069(.A1(new_n1228), .A2(new_n1269), .A3(new_n1215), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1270), .A2(new_n712), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1226), .B1(new_n1160), .B2(new_n1269), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1268), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(G384), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1273), .A2(G384), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1267), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT63), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1267), .A2(KEYINPUT63), .A3(new_n1277), .ZN(new_n1281));
  OAI211_X1 g1081(.A(G2897), .B(new_n1252), .C1(new_n1275), .C2(new_n1276), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1276), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1252), .A2(G2897), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1283), .A2(new_n1274), .A3(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1282), .A2(new_n1285), .ZN(new_n1286));
  OR2_X1    g1086(.A1(new_n1267), .A2(new_n1286), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1263), .A2(new_n1280), .A3(new_n1281), .A4(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT62), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1267), .A2(new_n1289), .A3(new_n1277), .ZN(new_n1290));
  XNOR2_X1  g1090(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1291), .B1(new_n1267), .B2(new_n1286), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1289), .B1(new_n1267), .B2(new_n1277), .ZN(new_n1293));
  NOR3_X1   g1093(.A1(new_n1290), .A2(new_n1292), .A3(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1259), .A2(new_n1261), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(KEYINPUT127), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT127), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1259), .A2(new_n1261), .A3(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1296), .A2(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1288), .B1(new_n1294), .B2(new_n1299), .ZN(G405));
  NAND2_X1  g1100(.A1(G375), .A2(new_n1248), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n1264), .ZN(new_n1302));
  OR2_X1    g1102(.A1(new_n1302), .A2(new_n1277), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1277), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1295), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1303), .A2(new_n1261), .A3(new_n1259), .A4(new_n1304), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(G402));
endmodule


