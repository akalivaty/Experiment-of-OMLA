

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U556 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U557 ( .A1(n969), .A2(G29), .ZN(n521) );
  OR2_X1 U558 ( .A1(n982), .A2(n713), .ZN(n712) );
  NAND2_X1 U559 ( .A1(n720), .A2(n719), .ZN(n723) );
  NOR2_X1 U560 ( .A1(n735), .A2(n758), .ZN(n736) );
  NAND2_X1 U561 ( .A1(n647), .A2(G54), .ZN(n587) );
  NOR2_X1 U562 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U563 ( .A(KEYINPUT15), .B(n594), .ZN(n595) );
  NOR2_X2 U564 ( .A1(G651), .A2(n630), .ZN(n647) );
  NOR2_X2 U565 ( .A1(n549), .A2(G2105), .ZN(n878) );
  XOR2_X1 U566 ( .A(KEYINPUT1), .B(n522), .Z(n648) );
  NOR2_X2 U567 ( .A1(n552), .A2(n551), .ZN(G160) );
  XOR2_X1 U568 ( .A(G543), .B(KEYINPUT0), .Z(n630) );
  NAND2_X1 U569 ( .A1(G51), .A2(n647), .ZN(n524) );
  INV_X1 U570 ( .A(G651), .ZN(n527) );
  NOR2_X1 U571 ( .A1(G543), .A2(n527), .ZN(n522) );
  NAND2_X1 U572 ( .A1(G63), .A2(n648), .ZN(n523) );
  NAND2_X1 U573 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U574 ( .A(KEYINPUT6), .B(n525), .ZN(n532) );
  NOR2_X1 U575 ( .A1(G543), .A2(G651), .ZN(n651) );
  NAND2_X1 U576 ( .A1(n651), .A2(G89), .ZN(n526) );
  XNOR2_X1 U577 ( .A(n526), .B(KEYINPUT4), .ZN(n529) );
  NOR2_X2 U578 ( .A1(n630), .A2(n527), .ZN(n655) );
  NAND2_X1 U579 ( .A1(G76), .A2(n655), .ZN(n528) );
  NAND2_X1 U580 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U581 ( .A(n530), .B(KEYINPUT5), .Z(n531) );
  NOR2_X1 U582 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U583 ( .A(KEYINPUT7), .B(n533), .Z(n534) );
  XOR2_X1 U584 ( .A(KEYINPUT77), .B(n534), .Z(G168) );
  XOR2_X1 U585 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U586 ( .A1(G91), .A2(n651), .ZN(n536) );
  NAND2_X1 U587 ( .A1(G53), .A2(n647), .ZN(n535) );
  NAND2_X1 U588 ( .A1(n536), .A2(n535), .ZN(n539) );
  NAND2_X1 U589 ( .A1(G78), .A2(n655), .ZN(n537) );
  XNOR2_X1 U590 ( .A(KEYINPUT69), .B(n537), .ZN(n538) );
  NOR2_X1 U591 ( .A1(n539), .A2(n538), .ZN(n541) );
  NAND2_X1 U592 ( .A1(n648), .A2(G65), .ZN(n540) );
  NAND2_X1 U593 ( .A1(n541), .A2(n540), .ZN(G299) );
  XNOR2_X1 U594 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n543) );
  NOR2_X1 U595 ( .A1(G2104), .A2(G2105), .ZN(n542) );
  XNOR2_X2 U596 ( .A(n543), .B(n542), .ZN(n877) );
  NAND2_X1 U597 ( .A1(G137), .A2(n877), .ZN(n545) );
  AND2_X1 U598 ( .A1(G2104), .A2(G2105), .ZN(n881) );
  NAND2_X1 U599 ( .A1(G113), .A2(n881), .ZN(n544) );
  NAND2_X1 U600 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U601 ( .A(KEYINPUT66), .B(n546), .Z(n548) );
  XOR2_X1 U602 ( .A(KEYINPUT64), .B(G2104), .Z(n549) );
  AND2_X1 U603 ( .A1(n549), .A2(G2105), .ZN(n882) );
  NAND2_X1 U604 ( .A1(n882), .A2(G125), .ZN(n547) );
  NAND2_X1 U605 ( .A1(n548), .A2(n547), .ZN(n552) );
  NAND2_X1 U606 ( .A1(G101), .A2(n878), .ZN(n550) );
  XNOR2_X1 U607 ( .A(KEYINPUT23), .B(n550), .ZN(n551) );
  NAND2_X1 U608 ( .A1(G114), .A2(n881), .ZN(n554) );
  NAND2_X1 U609 ( .A1(G126), .A2(n882), .ZN(n553) );
  NAND2_X1 U610 ( .A1(n554), .A2(n553), .ZN(n560) );
  INV_X1 U611 ( .A(KEYINPUT85), .ZN(n558) );
  NAND2_X1 U612 ( .A1(n878), .A2(G102), .ZN(n556) );
  NAND2_X1 U613 ( .A1(n877), .A2(G138), .ZN(n555) );
  NAND2_X1 U614 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U615 ( .A(n558), .B(n557), .ZN(n559) );
  NOR2_X1 U616 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U617 ( .A(KEYINPUT86), .B(n561), .ZN(n699) );
  BUF_X1 U618 ( .A(n699), .Z(G164) );
  AND2_X1 U619 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U620 ( .A(G860), .ZN(n619) );
  NAND2_X1 U621 ( .A1(n651), .A2(G81), .ZN(n562) );
  XNOR2_X1 U622 ( .A(n562), .B(KEYINPUT12), .ZN(n564) );
  NAND2_X1 U623 ( .A1(G68), .A2(n655), .ZN(n563) );
  NAND2_X1 U624 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U625 ( .A(n565), .B(KEYINPUT13), .ZN(n567) );
  NAND2_X1 U626 ( .A1(G43), .A2(n647), .ZN(n566) );
  NAND2_X1 U627 ( .A1(n567), .A2(n566), .ZN(n570) );
  NAND2_X1 U628 ( .A1(n648), .A2(G56), .ZN(n568) );
  XOR2_X1 U629 ( .A(KEYINPUT14), .B(n568), .Z(n569) );
  NOR2_X1 U630 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U631 ( .A(KEYINPUT72), .B(n571), .Z(n977) );
  OR2_X1 U632 ( .A1(n619), .A2(n977), .ZN(G153) );
  INV_X1 U633 ( .A(G132), .ZN(G219) );
  INV_X1 U634 ( .A(G120), .ZN(G236) );
  INV_X1 U635 ( .A(G69), .ZN(G235) );
  INV_X1 U636 ( .A(G108), .ZN(G238) );
  NAND2_X1 U637 ( .A1(G52), .A2(n647), .ZN(n572) );
  XOR2_X1 U638 ( .A(KEYINPUT68), .B(n572), .Z(n579) );
  NAND2_X1 U639 ( .A1(G90), .A2(n651), .ZN(n574) );
  NAND2_X1 U640 ( .A1(G77), .A2(n655), .ZN(n573) );
  NAND2_X1 U641 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n575), .B(KEYINPUT9), .ZN(n577) );
  NAND2_X1 U643 ( .A1(G64), .A2(n648), .ZN(n576) );
  NAND2_X1 U644 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U645 ( .A1(n579), .A2(n578), .ZN(G171) );
  XOR2_X1 U646 ( .A(KEYINPUT10), .B(KEYINPUT71), .Z(n581) );
  NAND2_X1 U647 ( .A1(G7), .A2(G661), .ZN(n580) );
  XNOR2_X1 U648 ( .A(n581), .B(n580), .ZN(G223) );
  INV_X1 U649 ( .A(G223), .ZN(n827) );
  NAND2_X1 U650 ( .A1(n827), .A2(G567), .ZN(n582) );
  XOR2_X1 U651 ( .A(KEYINPUT11), .B(n582), .Z(G234) );
  INV_X1 U652 ( .A(G171), .ZN(G301) );
  NAND2_X1 U653 ( .A1(G92), .A2(n651), .ZN(n584) );
  NAND2_X1 U654 ( .A1(G66), .A2(n648), .ZN(n583) );
  NAND2_X1 U655 ( .A1(n584), .A2(n583), .ZN(n593) );
  INV_X1 U656 ( .A(KEYINPUT73), .ZN(n586) );
  NAND2_X1 U657 ( .A1(n655), .A2(G79), .ZN(n585) );
  XNOR2_X1 U658 ( .A(n586), .B(n585), .ZN(n589) );
  XNOR2_X1 U659 ( .A(KEYINPUT74), .B(n587), .ZN(n588) );
  NAND2_X1 U660 ( .A1(n589), .A2(n588), .ZN(n591) );
  INV_X1 U661 ( .A(KEYINPUT75), .ZN(n590) );
  XNOR2_X1 U662 ( .A(n591), .B(n590), .ZN(n592) );
  INV_X1 U663 ( .A(n595), .ZN(n596) );
  XOR2_X1 U664 ( .A(KEYINPUT76), .B(n596), .Z(n901) );
  NOR2_X1 U665 ( .A1(n901), .A2(G868), .ZN(n598) );
  INV_X1 U666 ( .A(G868), .ZN(n599) );
  NOR2_X1 U667 ( .A1(n599), .A2(G301), .ZN(n597) );
  NOR2_X1 U668 ( .A1(n598), .A2(n597), .ZN(G284) );
  NOR2_X1 U669 ( .A1(G286), .A2(n599), .ZN(n601) );
  NOR2_X1 U670 ( .A1(G868), .A2(G299), .ZN(n600) );
  NOR2_X1 U671 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U672 ( .A(KEYINPUT78), .B(n602), .ZN(G297) );
  NAND2_X1 U673 ( .A1(n619), .A2(G559), .ZN(n603) );
  INV_X1 U674 ( .A(n901), .ZN(n982) );
  NAND2_X1 U675 ( .A1(n603), .A2(n982), .ZN(n604) );
  XNOR2_X1 U676 ( .A(n604), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U677 ( .A1(n977), .A2(G868), .ZN(n607) );
  NAND2_X1 U678 ( .A1(n982), .A2(G868), .ZN(n605) );
  NOR2_X1 U679 ( .A1(G559), .A2(n605), .ZN(n606) );
  NOR2_X1 U680 ( .A1(n607), .A2(n606), .ZN(G282) );
  XOR2_X1 U681 ( .A(G2100), .B(KEYINPUT80), .Z(n617) );
  NAND2_X1 U682 ( .A1(G135), .A2(n877), .ZN(n609) );
  NAND2_X1 U683 ( .A1(G111), .A2(n881), .ZN(n608) );
  NAND2_X1 U684 ( .A1(n609), .A2(n608), .ZN(n612) );
  NAND2_X1 U685 ( .A1(n882), .A2(G123), .ZN(n610) );
  XOR2_X1 U686 ( .A(KEYINPUT18), .B(n610), .Z(n611) );
  NOR2_X1 U687 ( .A1(n612), .A2(n611), .ZN(n614) );
  NAND2_X1 U688 ( .A1(n878), .A2(G99), .ZN(n613) );
  NAND2_X1 U689 ( .A1(n614), .A2(n613), .ZN(n957) );
  XNOR2_X1 U690 ( .A(KEYINPUT79), .B(n957), .ZN(n615) );
  XNOR2_X1 U691 ( .A(n615), .B(G2096), .ZN(n616) );
  NAND2_X1 U692 ( .A1(n617), .A2(n616), .ZN(G156) );
  NAND2_X1 U693 ( .A1(n982), .A2(G559), .ZN(n618) );
  XOR2_X1 U694 ( .A(n977), .B(n618), .Z(n663) );
  NAND2_X1 U695 ( .A1(n619), .A2(n663), .ZN(n626) );
  NAND2_X1 U696 ( .A1(G55), .A2(n647), .ZN(n621) );
  NAND2_X1 U697 ( .A1(G67), .A2(n648), .ZN(n620) );
  NAND2_X1 U698 ( .A1(n621), .A2(n620), .ZN(n625) );
  NAND2_X1 U699 ( .A1(G93), .A2(n651), .ZN(n623) );
  NAND2_X1 U700 ( .A1(G80), .A2(n655), .ZN(n622) );
  NAND2_X1 U701 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U702 ( .A1(n625), .A2(n624), .ZN(n666) );
  XOR2_X1 U703 ( .A(n626), .B(n666), .Z(G145) );
  NAND2_X1 U704 ( .A1(G49), .A2(n647), .ZN(n628) );
  NAND2_X1 U705 ( .A1(G74), .A2(G651), .ZN(n627) );
  NAND2_X1 U706 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U707 ( .A1(n648), .A2(n629), .ZN(n632) );
  NAND2_X1 U708 ( .A1(n630), .A2(G87), .ZN(n631) );
  NAND2_X1 U709 ( .A1(n632), .A2(n631), .ZN(G288) );
  NAND2_X1 U710 ( .A1(G88), .A2(n651), .ZN(n634) );
  NAND2_X1 U711 ( .A1(G75), .A2(n655), .ZN(n633) );
  NAND2_X1 U712 ( .A1(n634), .A2(n633), .ZN(n639) );
  NAND2_X1 U713 ( .A1(G62), .A2(n648), .ZN(n635) );
  XOR2_X1 U714 ( .A(KEYINPUT81), .B(n635), .Z(n637) );
  NAND2_X1 U715 ( .A1(n647), .A2(G50), .ZN(n636) );
  NAND2_X1 U716 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U717 ( .A1(n639), .A2(n638), .ZN(G166) );
  NAND2_X1 U718 ( .A1(G86), .A2(n651), .ZN(n641) );
  NAND2_X1 U719 ( .A1(G48), .A2(n647), .ZN(n640) );
  NAND2_X1 U720 ( .A1(n641), .A2(n640), .ZN(n644) );
  NAND2_X1 U721 ( .A1(n655), .A2(G73), .ZN(n642) );
  XOR2_X1 U722 ( .A(KEYINPUT2), .B(n642), .Z(n643) );
  NOR2_X1 U723 ( .A1(n644), .A2(n643), .ZN(n646) );
  NAND2_X1 U724 ( .A1(n648), .A2(G61), .ZN(n645) );
  NAND2_X1 U725 ( .A1(n646), .A2(n645), .ZN(G305) );
  NAND2_X1 U726 ( .A1(G47), .A2(n647), .ZN(n650) );
  NAND2_X1 U727 ( .A1(G60), .A2(n648), .ZN(n649) );
  NAND2_X1 U728 ( .A1(n650), .A2(n649), .ZN(n654) );
  NAND2_X1 U729 ( .A1(G85), .A2(n651), .ZN(n652) );
  XNOR2_X1 U730 ( .A(KEYINPUT67), .B(n652), .ZN(n653) );
  NOR2_X1 U731 ( .A1(n654), .A2(n653), .ZN(n657) );
  NAND2_X1 U732 ( .A1(n655), .A2(G72), .ZN(n656) );
  NAND2_X1 U733 ( .A1(n657), .A2(n656), .ZN(G290) );
  XNOR2_X1 U734 ( .A(KEYINPUT19), .B(G288), .ZN(n662) );
  XNOR2_X1 U735 ( .A(G166), .B(G299), .ZN(n658) );
  XNOR2_X1 U736 ( .A(n658), .B(G305), .ZN(n659) );
  XNOR2_X1 U737 ( .A(n666), .B(n659), .ZN(n660) );
  XNOR2_X1 U738 ( .A(n660), .B(G290), .ZN(n661) );
  XNOR2_X1 U739 ( .A(n662), .B(n661), .ZN(n898) );
  XNOR2_X1 U740 ( .A(KEYINPUT82), .B(n663), .ZN(n664) );
  XNOR2_X1 U741 ( .A(n898), .B(n664), .ZN(n665) );
  NAND2_X1 U742 ( .A1(n665), .A2(G868), .ZN(n668) );
  OR2_X1 U743 ( .A1(G868), .A2(n666), .ZN(n667) );
  NAND2_X1 U744 ( .A1(n668), .A2(n667), .ZN(G295) );
  NAND2_X1 U745 ( .A1(G2078), .A2(G2084), .ZN(n669) );
  XNOR2_X1 U746 ( .A(n669), .B(KEYINPUT20), .ZN(n670) );
  XNOR2_X1 U747 ( .A(n670), .B(KEYINPUT83), .ZN(n671) );
  NAND2_X1 U748 ( .A1(n671), .A2(G2090), .ZN(n672) );
  XNOR2_X1 U749 ( .A(KEYINPUT21), .B(n672), .ZN(n673) );
  NAND2_X1 U750 ( .A1(n673), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U751 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U752 ( .A(KEYINPUT70), .B(G82), .Z(G220) );
  NOR2_X1 U753 ( .A1(G235), .A2(G236), .ZN(n674) );
  XOR2_X1 U754 ( .A(KEYINPUT84), .B(n674), .Z(n675) );
  NOR2_X1 U755 ( .A1(G238), .A2(n675), .ZN(n676) );
  NAND2_X1 U756 ( .A1(G57), .A2(n676), .ZN(n833) );
  NAND2_X1 U757 ( .A1(n833), .A2(G567), .ZN(n681) );
  NOR2_X1 U758 ( .A1(G220), .A2(G219), .ZN(n677) );
  XOR2_X1 U759 ( .A(KEYINPUT22), .B(n677), .Z(n678) );
  NOR2_X1 U760 ( .A1(G218), .A2(n678), .ZN(n679) );
  NAND2_X1 U761 ( .A1(G96), .A2(n679), .ZN(n834) );
  NAND2_X1 U762 ( .A1(n834), .A2(G2106), .ZN(n680) );
  NAND2_X1 U763 ( .A1(n681), .A2(n680), .ZN(n835) );
  NAND2_X1 U764 ( .A1(G483), .A2(G661), .ZN(n682) );
  NOR2_X1 U765 ( .A1(n835), .A2(n682), .ZN(n832) );
  NAND2_X1 U766 ( .A1(n832), .A2(G36), .ZN(G176) );
  XNOR2_X1 U767 ( .A(KEYINPUT87), .B(G166), .ZN(G303) );
  NAND2_X1 U768 ( .A1(G131), .A2(n877), .ZN(n684) );
  NAND2_X1 U769 ( .A1(G95), .A2(n878), .ZN(n683) );
  NAND2_X1 U770 ( .A1(n684), .A2(n683), .ZN(n688) );
  NAND2_X1 U771 ( .A1(G107), .A2(n881), .ZN(n686) );
  NAND2_X1 U772 ( .A1(G119), .A2(n882), .ZN(n685) );
  NAND2_X1 U773 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U774 ( .A1(n688), .A2(n687), .ZN(n864) );
  INV_X1 U775 ( .A(G1991), .ZN(n925) );
  NOR2_X1 U776 ( .A1(n864), .A2(n925), .ZN(n698) );
  XOR2_X1 U777 ( .A(KEYINPUT92), .B(KEYINPUT38), .Z(n690) );
  NAND2_X1 U778 ( .A1(G105), .A2(n878), .ZN(n689) );
  XNOR2_X1 U779 ( .A(n690), .B(n689), .ZN(n694) );
  NAND2_X1 U780 ( .A1(G141), .A2(n877), .ZN(n692) );
  NAND2_X1 U781 ( .A1(G117), .A2(n881), .ZN(n691) );
  NAND2_X1 U782 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U783 ( .A1(n694), .A2(n693), .ZN(n696) );
  NAND2_X1 U784 ( .A1(n882), .A2(G129), .ZN(n695) );
  NAND2_X1 U785 ( .A1(n696), .A2(n695), .ZN(n891) );
  AND2_X1 U786 ( .A1(n891), .A2(G1996), .ZN(n697) );
  NOR2_X1 U787 ( .A1(n698), .A2(n697), .ZN(n949) );
  NOR2_X2 U788 ( .A1(G1384), .A2(n699), .ZN(n703) );
  NAND2_X1 U789 ( .A1(G160), .A2(G40), .ZN(n701) );
  NOR2_X1 U790 ( .A1(n703), .A2(n701), .ZN(n821) );
  INV_X1 U791 ( .A(n821), .ZN(n700) );
  NOR2_X1 U792 ( .A1(n949), .A2(n700), .ZN(n815) );
  INV_X1 U793 ( .A(n815), .ZN(n794) );
  INV_X1 U794 ( .A(n701), .ZN(n702) );
  NAND2_X2 U795 ( .A1(n703), .A2(n702), .ZN(n746) );
  NAND2_X1 U796 ( .A1(G1348), .A2(n746), .ZN(n705) );
  INV_X1 U797 ( .A(n746), .ZN(n729) );
  NAND2_X1 U798 ( .A1(G2067), .A2(n729), .ZN(n704) );
  NAND2_X1 U799 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U800 ( .A(KEYINPUT97), .B(n706), .ZN(n713) );
  INV_X1 U801 ( .A(G1996), .ZN(n922) );
  NOR2_X1 U802 ( .A1(n746), .A2(n922), .ZN(n707) );
  XOR2_X1 U803 ( .A(n707), .B(KEYINPUT26), .Z(n709) );
  NAND2_X1 U804 ( .A1(n746), .A2(G1341), .ZN(n708) );
  NAND2_X1 U805 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U806 ( .A1(n977), .A2(n710), .ZN(n711) );
  NAND2_X1 U807 ( .A1(n712), .A2(n711), .ZN(n715) );
  NAND2_X1 U808 ( .A1(n982), .A2(n713), .ZN(n714) );
  NAND2_X1 U809 ( .A1(n715), .A2(n714), .ZN(n722) );
  INV_X1 U810 ( .A(KEYINPUT27), .ZN(n717) );
  NAND2_X1 U811 ( .A1(n729), .A2(G2072), .ZN(n716) );
  XNOR2_X1 U812 ( .A(n717), .B(n716), .ZN(n720) );
  NAND2_X1 U813 ( .A1(G1956), .A2(n746), .ZN(n718) );
  XNOR2_X1 U814 ( .A(KEYINPUT96), .B(n718), .ZN(n719) );
  NOR2_X1 U815 ( .A1(G299), .A2(n723), .ZN(n721) );
  NOR2_X1 U816 ( .A1(n722), .A2(n721), .ZN(n726) );
  NAND2_X1 U817 ( .A1(n723), .A2(G299), .ZN(n724) );
  XOR2_X1 U818 ( .A(KEYINPUT28), .B(n724), .Z(n725) );
  NOR2_X1 U819 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U820 ( .A(n727), .B(KEYINPUT29), .ZN(n733) );
  XNOR2_X1 U821 ( .A(G1961), .B(KEYINPUT94), .ZN(n1008) );
  NOR2_X1 U822 ( .A1(n729), .A2(n1008), .ZN(n728) );
  XNOR2_X1 U823 ( .A(n728), .B(KEYINPUT95), .ZN(n731) );
  XNOR2_X1 U824 ( .A(KEYINPUT25), .B(G2078), .ZN(n927) );
  NAND2_X1 U825 ( .A1(n729), .A2(n927), .ZN(n730) );
  NAND2_X1 U826 ( .A1(n731), .A2(n730), .ZN(n738) );
  NAND2_X1 U827 ( .A1(G171), .A2(n738), .ZN(n732) );
  NAND2_X1 U828 ( .A1(n733), .A2(n732), .ZN(n743) );
  NOR2_X1 U829 ( .A1(n746), .A2(G2084), .ZN(n734) );
  XNOR2_X1 U830 ( .A(n734), .B(KEYINPUT93), .ZN(n754) );
  NAND2_X1 U831 ( .A1(G8), .A2(n754), .ZN(n735) );
  NAND2_X1 U832 ( .A1(G8), .A2(n746), .ZN(n787) );
  NOR2_X1 U833 ( .A1(G1966), .A2(n787), .ZN(n758) );
  XOR2_X1 U834 ( .A(KEYINPUT30), .B(n736), .Z(n737) );
  NOR2_X1 U835 ( .A1(G168), .A2(n737), .ZN(n740) );
  NOR2_X1 U836 ( .A1(G171), .A2(n738), .ZN(n739) );
  NOR2_X1 U837 ( .A1(n740), .A2(n739), .ZN(n741) );
  XOR2_X1 U838 ( .A(KEYINPUT31), .B(n741), .Z(n742) );
  NAND2_X1 U839 ( .A1(n743), .A2(n742), .ZN(n756) );
  NAND2_X1 U840 ( .A1(n756), .A2(G286), .ZN(n744) );
  XNOR2_X1 U841 ( .A(n744), .B(KEYINPUT98), .ZN(n751) );
  NOR2_X1 U842 ( .A1(G1971), .A2(n787), .ZN(n745) );
  XOR2_X1 U843 ( .A(KEYINPUT99), .B(n745), .Z(n748) );
  NOR2_X1 U844 ( .A1(G2090), .A2(n746), .ZN(n747) );
  NOR2_X1 U845 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U846 ( .A1(n749), .A2(G303), .ZN(n750) );
  NAND2_X1 U847 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U848 ( .A1(n752), .A2(G8), .ZN(n753) );
  XNOR2_X1 U849 ( .A(n753), .B(KEYINPUT32), .ZN(n782) );
  INV_X1 U850 ( .A(n754), .ZN(n755) );
  NAND2_X1 U851 ( .A1(G8), .A2(n755), .ZN(n760) );
  INV_X1 U852 ( .A(n756), .ZN(n757) );
  NOR2_X1 U853 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U854 ( .A1(n760), .A2(n759), .ZN(n783) );
  NAND2_X1 U855 ( .A1(G1976), .A2(G288), .ZN(n980) );
  AND2_X1 U856 ( .A1(n783), .A2(n980), .ZN(n761) );
  NAND2_X1 U857 ( .A1(n782), .A2(n761), .ZN(n765) );
  INV_X1 U858 ( .A(n980), .ZN(n763) );
  NOR2_X1 U859 ( .A1(G1976), .A2(G288), .ZN(n770) );
  NOR2_X1 U860 ( .A1(G1971), .A2(G303), .ZN(n762) );
  NOR2_X1 U861 ( .A1(n770), .A2(n762), .ZN(n984) );
  OR2_X1 U862 ( .A1(n763), .A2(n984), .ZN(n764) );
  AND2_X1 U863 ( .A1(n765), .A2(n764), .ZN(n767) );
  INV_X1 U864 ( .A(KEYINPUT100), .ZN(n769) );
  OR2_X1 U865 ( .A1(n787), .A2(n769), .ZN(n766) );
  NOR2_X1 U866 ( .A1(KEYINPUT33), .A2(n768), .ZN(n776) );
  NAND2_X1 U867 ( .A1(n769), .A2(n770), .ZN(n773) );
  NAND2_X1 U868 ( .A1(n770), .A2(KEYINPUT33), .ZN(n771) );
  NAND2_X1 U869 ( .A1(n771), .A2(KEYINPUT100), .ZN(n772) );
  NAND2_X1 U870 ( .A1(n773), .A2(n772), .ZN(n774) );
  NOR2_X1 U871 ( .A1(n787), .A2(n774), .ZN(n775) );
  NOR2_X1 U872 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U873 ( .A(G1981), .B(G305), .Z(n971) );
  NAND2_X1 U874 ( .A1(n777), .A2(n971), .ZN(n792) );
  NOR2_X1 U875 ( .A1(G1981), .A2(G305), .ZN(n778) );
  XOR2_X1 U876 ( .A(n778), .B(KEYINPUT24), .Z(n779) );
  OR2_X1 U877 ( .A1(n787), .A2(n779), .ZN(n790) );
  NOR2_X1 U878 ( .A1(G2090), .A2(G303), .ZN(n780) );
  NAND2_X1 U879 ( .A1(G8), .A2(n780), .ZN(n781) );
  XOR2_X1 U880 ( .A(KEYINPUT101), .B(n781), .Z(n785) );
  NAND2_X1 U881 ( .A1(n783), .A2(n782), .ZN(n784) );
  NAND2_X1 U882 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U883 ( .A(n786), .B(KEYINPUT102), .ZN(n788) );
  NAND2_X1 U884 ( .A1(n788), .A2(n787), .ZN(n789) );
  AND2_X1 U885 ( .A1(n790), .A2(n789), .ZN(n791) );
  NAND2_X1 U886 ( .A1(n792), .A2(n791), .ZN(n793) );
  AND2_X1 U887 ( .A1(n794), .A2(n793), .ZN(n810) );
  XOR2_X1 U888 ( .A(G2067), .B(KEYINPUT37), .Z(n795) );
  XNOR2_X1 U889 ( .A(KEYINPUT89), .B(n795), .ZN(n811) );
  NAND2_X1 U890 ( .A1(G140), .A2(n877), .ZN(n797) );
  NAND2_X1 U891 ( .A1(G104), .A2(n878), .ZN(n796) );
  NAND2_X1 U892 ( .A1(n797), .A2(n796), .ZN(n798) );
  XNOR2_X1 U893 ( .A(KEYINPUT34), .B(n798), .ZN(n803) );
  NAND2_X1 U894 ( .A1(G116), .A2(n881), .ZN(n800) );
  NAND2_X1 U895 ( .A1(G128), .A2(n882), .ZN(n799) );
  NAND2_X1 U896 ( .A1(n800), .A2(n799), .ZN(n801) );
  XOR2_X1 U897 ( .A(n801), .B(KEYINPUT35), .Z(n802) );
  NOR2_X1 U898 ( .A1(n803), .A2(n802), .ZN(n804) );
  XOR2_X1 U899 ( .A(KEYINPUT36), .B(n804), .Z(n805) );
  XOR2_X1 U900 ( .A(KEYINPUT90), .B(n805), .Z(n895) );
  NOR2_X1 U901 ( .A1(n811), .A2(n895), .ZN(n806) );
  XNOR2_X1 U902 ( .A(n806), .B(KEYINPUT91), .ZN(n964) );
  XOR2_X1 U903 ( .A(G1986), .B(KEYINPUT88), .Z(n807) );
  XNOR2_X1 U904 ( .A(G290), .B(n807), .ZN(n975) );
  NAND2_X1 U905 ( .A1(n964), .A2(n975), .ZN(n808) );
  NAND2_X1 U906 ( .A1(n808), .A2(n821), .ZN(n809) );
  NAND2_X1 U907 ( .A1(n810), .A2(n809), .ZN(n824) );
  NAND2_X1 U908 ( .A1(n895), .A2(n811), .ZN(n948) );
  NOR2_X1 U909 ( .A1(G1996), .A2(n891), .ZN(n812) );
  XOR2_X1 U910 ( .A(KEYINPUT103), .B(n812), .Z(n951) );
  NOR2_X1 U911 ( .A1(G1986), .A2(G290), .ZN(n813) );
  AND2_X1 U912 ( .A1(n925), .A2(n864), .ZN(n960) );
  NOR2_X1 U913 ( .A1(n813), .A2(n960), .ZN(n814) );
  NOR2_X1 U914 ( .A1(n815), .A2(n814), .ZN(n816) );
  NOR2_X1 U915 ( .A1(n951), .A2(n816), .ZN(n817) );
  XNOR2_X1 U916 ( .A(KEYINPUT104), .B(n817), .ZN(n818) );
  XNOR2_X1 U917 ( .A(n818), .B(KEYINPUT39), .ZN(n819) );
  NAND2_X1 U918 ( .A1(n819), .A2(n964), .ZN(n820) );
  NAND2_X1 U919 ( .A1(n948), .A2(n820), .ZN(n822) );
  NAND2_X1 U920 ( .A1(n822), .A2(n821), .ZN(n823) );
  NAND2_X1 U921 ( .A1(n824), .A2(n823), .ZN(n826) );
  XOR2_X1 U922 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n825) );
  XNOR2_X1 U923 ( .A(n826), .B(n825), .ZN(G329) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n827), .ZN(G217) );
  NAND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n828) );
  XOR2_X1 U926 ( .A(KEYINPUT108), .B(n828), .Z(n829) );
  NAND2_X1 U927 ( .A1(n829), .A2(G661), .ZN(n830) );
  XOR2_X1 U928 ( .A(KEYINPUT109), .B(n830), .Z(G259) );
  NAND2_X1 U929 ( .A1(G3), .A2(G1), .ZN(n831) );
  NAND2_X1 U930 ( .A1(n832), .A2(n831), .ZN(G188) );
  XOR2_X1 U931 ( .A(G96), .B(KEYINPUT110), .Z(G221) );
  NOR2_X1 U933 ( .A1(n834), .A2(n833), .ZN(G325) );
  INV_X1 U934 ( .A(G325), .ZN(G261) );
  INV_X1 U935 ( .A(n835), .ZN(G319) );
  XOR2_X1 U936 ( .A(KEYINPUT112), .B(KEYINPUT111), .Z(n837) );
  XNOR2_X1 U937 ( .A(G2678), .B(KEYINPUT43), .ZN(n836) );
  XNOR2_X1 U938 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U939 ( .A(KEYINPUT42), .B(G2090), .Z(n839) );
  XNOR2_X1 U940 ( .A(G2067), .B(G2072), .ZN(n838) );
  XNOR2_X1 U941 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U942 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U943 ( .A(G2100), .B(G2096), .ZN(n842) );
  XNOR2_X1 U944 ( .A(n843), .B(n842), .ZN(n845) );
  XOR2_X1 U945 ( .A(G2078), .B(G2084), .Z(n844) );
  XNOR2_X1 U946 ( .A(n845), .B(n844), .ZN(G227) );
  XOR2_X1 U947 ( .A(G1981), .B(G1956), .Z(n847) );
  XNOR2_X1 U948 ( .A(G1996), .B(G1966), .ZN(n846) );
  XNOR2_X1 U949 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U950 ( .A(G1976), .B(G1971), .Z(n849) );
  XNOR2_X1 U951 ( .A(G1986), .B(G1961), .ZN(n848) );
  XNOR2_X1 U952 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U953 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U954 ( .A(KEYINPUT113), .B(G2474), .ZN(n852) );
  XNOR2_X1 U955 ( .A(n853), .B(n852), .ZN(n854) );
  XNOR2_X1 U956 ( .A(KEYINPUT41), .B(n854), .ZN(n855) );
  XNOR2_X1 U957 ( .A(n855), .B(n925), .ZN(G229) );
  NAND2_X1 U958 ( .A1(G100), .A2(n878), .ZN(n857) );
  NAND2_X1 U959 ( .A1(G112), .A2(n881), .ZN(n856) );
  NAND2_X1 U960 ( .A1(n857), .A2(n856), .ZN(n863) );
  NAND2_X1 U961 ( .A1(G124), .A2(n882), .ZN(n858) );
  XNOR2_X1 U962 ( .A(n858), .B(KEYINPUT44), .ZN(n861) );
  NAND2_X1 U963 ( .A1(G136), .A2(n877), .ZN(n859) );
  XNOR2_X1 U964 ( .A(n859), .B(KEYINPUT114), .ZN(n860) );
  NAND2_X1 U965 ( .A1(n861), .A2(n860), .ZN(n862) );
  NOR2_X1 U966 ( .A1(n863), .A2(n862), .ZN(G162) );
  XOR2_X1 U967 ( .A(KEYINPUT48), .B(KEYINPUT116), .Z(n866) );
  XNOR2_X1 U968 ( .A(n864), .B(KEYINPUT46), .ZN(n865) );
  XNOR2_X1 U969 ( .A(n866), .B(n865), .ZN(n876) );
  NAND2_X1 U970 ( .A1(G118), .A2(n881), .ZN(n868) );
  NAND2_X1 U971 ( .A1(G130), .A2(n882), .ZN(n867) );
  NAND2_X1 U972 ( .A1(n868), .A2(n867), .ZN(n874) );
  NAND2_X1 U973 ( .A1(G142), .A2(n877), .ZN(n870) );
  NAND2_X1 U974 ( .A1(G106), .A2(n878), .ZN(n869) );
  NAND2_X1 U975 ( .A1(n870), .A2(n869), .ZN(n871) );
  XNOR2_X1 U976 ( .A(KEYINPUT115), .B(n871), .ZN(n872) );
  XNOR2_X1 U977 ( .A(KEYINPUT45), .B(n872), .ZN(n873) );
  NOR2_X1 U978 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U979 ( .A(n876), .B(n875), .Z(n889) );
  NAND2_X1 U980 ( .A1(G139), .A2(n877), .ZN(n880) );
  NAND2_X1 U981 ( .A1(G103), .A2(n878), .ZN(n879) );
  NAND2_X1 U982 ( .A1(n880), .A2(n879), .ZN(n887) );
  NAND2_X1 U983 ( .A1(G115), .A2(n881), .ZN(n884) );
  NAND2_X1 U984 ( .A1(G127), .A2(n882), .ZN(n883) );
  NAND2_X1 U985 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U986 ( .A(KEYINPUT47), .B(n885), .Z(n886) );
  NOR2_X1 U987 ( .A1(n887), .A2(n886), .ZN(n944) );
  XNOR2_X1 U988 ( .A(n944), .B(G162), .ZN(n888) );
  XNOR2_X1 U989 ( .A(n889), .B(n888), .ZN(n890) );
  XNOR2_X1 U990 ( .A(n957), .B(n890), .ZN(n893) );
  XOR2_X1 U991 ( .A(G160), .B(n891), .Z(n892) );
  XNOR2_X1 U992 ( .A(n893), .B(n892), .ZN(n894) );
  XOR2_X1 U993 ( .A(n895), .B(n894), .Z(n896) );
  XNOR2_X1 U994 ( .A(G164), .B(n896), .ZN(n897) );
  NOR2_X1 U995 ( .A1(G37), .A2(n897), .ZN(G395) );
  XOR2_X1 U996 ( .A(n898), .B(G286), .Z(n900) );
  XNOR2_X1 U997 ( .A(G171), .B(n977), .ZN(n899) );
  XNOR2_X1 U998 ( .A(n900), .B(n899), .ZN(n902) );
  XNOR2_X1 U999 ( .A(n902), .B(n901), .ZN(n903) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n903), .ZN(G397) );
  XNOR2_X1 U1001 ( .A(G2427), .B(KEYINPUT106), .ZN(n913) );
  XOR2_X1 U1002 ( .A(G2430), .B(G2446), .Z(n905) );
  XNOR2_X1 U1003 ( .A(G2435), .B(G2438), .ZN(n904) );
  XNOR2_X1 U1004 ( .A(n905), .B(n904), .ZN(n909) );
  XOR2_X1 U1005 ( .A(G2454), .B(KEYINPUT107), .Z(n907) );
  XNOR2_X1 U1006 ( .A(G1341), .B(G1348), .ZN(n906) );
  XNOR2_X1 U1007 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1008 ( .A(n909), .B(n908), .Z(n911) );
  XNOR2_X1 U1009 ( .A(G2451), .B(G2443), .ZN(n910) );
  XNOR2_X1 U1010 ( .A(n911), .B(n910), .ZN(n912) );
  XNOR2_X1 U1011 ( .A(n913), .B(n912), .ZN(n914) );
  NAND2_X1 U1012 ( .A1(n914), .A2(G14), .ZN(n920) );
  NAND2_X1 U1013 ( .A1(G319), .A2(n920), .ZN(n917) );
  NOR2_X1 U1014 ( .A1(G227), .A2(G229), .ZN(n915) );
  XNOR2_X1 U1015 ( .A(KEYINPUT49), .B(n915), .ZN(n916) );
  NOR2_X1 U1016 ( .A1(n917), .A2(n916), .ZN(n919) );
  NOR2_X1 U1017 ( .A1(G395), .A2(G397), .ZN(n918) );
  NAND2_X1 U1018 ( .A1(n919), .A2(n918), .ZN(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  INV_X1 U1020 ( .A(G57), .ZN(G237) );
  INV_X1 U1021 ( .A(n920), .ZN(G401) );
  XOR2_X1 U1022 ( .A(KEYINPUT55), .B(KEYINPUT120), .Z(n943) );
  XOR2_X1 U1023 ( .A(KEYINPUT54), .B(G34), .Z(n921) );
  XNOR2_X1 U1024 ( .A(n921), .B(G2084), .ZN(n939) );
  XNOR2_X1 U1025 ( .A(G2090), .B(G35), .ZN(n937) );
  XOR2_X1 U1026 ( .A(G2067), .B(G26), .Z(n924) );
  XNOR2_X1 U1027 ( .A(n922), .B(G32), .ZN(n923) );
  NAND2_X1 U1028 ( .A1(n924), .A2(n923), .ZN(n934) );
  XNOR2_X1 U1029 ( .A(G25), .B(n925), .ZN(n932) );
  XOR2_X1 U1030 ( .A(G2072), .B(G33), .Z(n926) );
  NAND2_X1 U1031 ( .A1(n926), .A2(G28), .ZN(n930) );
  XNOR2_X1 U1032 ( .A(G27), .B(n927), .ZN(n928) );
  XNOR2_X1 U1033 ( .A(KEYINPUT121), .B(n928), .ZN(n929) );
  NOR2_X1 U1034 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1035 ( .A1(n932), .A2(n931), .ZN(n933) );
  NOR2_X1 U1036 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1037 ( .A(KEYINPUT53), .B(n935), .ZN(n936) );
  NOR2_X1 U1038 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1039 ( .A1(n939), .A2(n938), .ZN(n941) );
  INV_X1 U1040 ( .A(G29), .ZN(n940) );
  NAND2_X1 U1041 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1042 ( .A(n943), .B(n942), .ZN(n970) );
  XOR2_X1 U1043 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n967) );
  XOR2_X1 U1044 ( .A(G2072), .B(n944), .Z(n946) );
  XOR2_X1 U1045 ( .A(G164), .B(G2078), .Z(n945) );
  NOR2_X1 U1046 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1047 ( .A(KEYINPUT50), .B(n947), .ZN(n956) );
  NAND2_X1 U1048 ( .A1(n949), .A2(n948), .ZN(n954) );
  XOR2_X1 U1049 ( .A(G2090), .B(G162), .Z(n950) );
  NOR2_X1 U1050 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1051 ( .A(n952), .B(KEYINPUT51), .ZN(n953) );
  NOR2_X1 U1052 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n963) );
  XNOR2_X1 U1054 ( .A(G160), .B(G2084), .ZN(n958) );
  NAND2_X1 U1055 ( .A1(n958), .A2(n957), .ZN(n959) );
  NOR2_X1 U1056 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1057 ( .A(KEYINPUT117), .B(n961), .ZN(n962) );
  NOR2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n965) );
  NAND2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1060 ( .A(n967), .B(n966), .ZN(n968) );
  XNOR2_X1 U1061 ( .A(KEYINPUT52), .B(n968), .ZN(n969) );
  NAND2_X1 U1062 ( .A1(n970), .A2(n521), .ZN(n1025) );
  XNOR2_X1 U1063 ( .A(KEYINPUT56), .B(G16), .ZN(n994) );
  XNOR2_X1 U1064 ( .A(G1966), .B(G168), .ZN(n972) );
  NAND2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1066 ( .A(n973), .B(KEYINPUT57), .ZN(n992) );
  XOR2_X1 U1067 ( .A(G1956), .B(KEYINPUT122), .Z(n974) );
  XNOR2_X1 U1068 ( .A(G299), .B(n974), .ZN(n976) );
  NAND2_X1 U1069 ( .A1(n976), .A2(n975), .ZN(n979) );
  XNOR2_X1 U1070 ( .A(G1341), .B(n977), .ZN(n978) );
  NOR2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n981) );
  NAND2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n990) );
  XNOR2_X1 U1073 ( .A(G1348), .B(n982), .ZN(n988) );
  NAND2_X1 U1074 ( .A1(G1971), .A2(G303), .ZN(n983) );
  NAND2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n986) );
  XNOR2_X1 U1076 ( .A(G1961), .B(G301), .ZN(n985) );
  NOR2_X1 U1077 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1078 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1079 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1080 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1081 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1082 ( .A(n995), .B(KEYINPUT123), .ZN(n1022) );
  XOR2_X1 U1083 ( .A(KEYINPUT125), .B(G4), .Z(n997) );
  XNOR2_X1 U1084 ( .A(G1348), .B(KEYINPUT59), .ZN(n996) );
  XNOR2_X1 U1085 ( .A(n997), .B(n996), .ZN(n1001) );
  XNOR2_X1 U1086 ( .A(G1341), .B(G19), .ZN(n999) );
  XNOR2_X1 U1087 ( .A(G1981), .B(G6), .ZN(n998) );
  NOR2_X1 U1088 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1089 ( .A1(n1001), .A2(n1000), .ZN(n1004) );
  XNOR2_X1 U1090 ( .A(G20), .B(G1956), .ZN(n1002) );
  XNOR2_X1 U1091 ( .A(KEYINPUT124), .B(n1002), .ZN(n1003) );
  NOR2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1093 ( .A(KEYINPUT60), .B(n1005), .Z(n1007) );
  XNOR2_X1 U1094 ( .A(G1966), .B(G21), .ZN(n1006) );
  NOR2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1018) );
  XNOR2_X1 U1096 ( .A(n1008), .B(G5), .ZN(n1016) );
  XOR2_X1 U1097 ( .A(G1986), .B(G24), .Z(n1013) );
  XNOR2_X1 U1098 ( .A(G1971), .B(G22), .ZN(n1010) );
  XNOR2_X1 U1099 ( .A(G23), .B(G1976), .ZN(n1009) );
  NOR2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1101 ( .A(n1011), .B(KEYINPUT126), .ZN(n1012) );
  NAND2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1103 ( .A(n1014), .B(KEYINPUT58), .ZN(n1015) );
  NOR2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1106 ( .A(KEYINPUT61), .B(n1019), .ZN(n1020) );
  NOR2_X1 U1107 ( .A1(n1020), .A2(G16), .ZN(n1021) );
  NOR2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1109 ( .A(n1023), .B(KEYINPUT127), .ZN(n1024) );
  NOR2_X1 U1110 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1111 ( .A1(n1026), .A2(G11), .ZN(n1027) );
  XOR2_X1 U1112 ( .A(KEYINPUT62), .B(n1027), .Z(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
endmodule

