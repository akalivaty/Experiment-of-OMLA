

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U560 ( .A(n716), .B(KEYINPUT64), .ZN(n742) );
  BUF_X1 U561 ( .A(n742), .Z(n526) );
  NOR2_X1 U562 ( .A1(KEYINPUT33), .A2(n528), .ZN(n803) );
  XNOR2_X1 U563 ( .A(n731), .B(n730), .ZN(n778) );
  NOR2_X1 U564 ( .A1(n721), .A2(G168), .ZN(n723) );
  NOR2_X1 U565 ( .A1(n534), .A2(n1007), .ZN(n741) );
  AND2_X1 U566 ( .A1(n739), .A2(n738), .ZN(n534) );
  INV_X1 U567 ( .A(G164), .ZN(n535) );
  NOR2_X1 U568 ( .A1(n540), .A2(n578), .ZN(n536) );
  NOR2_X4 U569 ( .A1(G2105), .A2(n564), .ZN(n569) );
  NAND2_X1 U570 ( .A1(n529), .A2(n541), .ZN(n540) );
  INV_X1 U571 ( .A(G1384), .ZN(n541) );
  INV_X1 U572 ( .A(KEYINPUT101), .ZN(n552) );
  AND2_X1 U573 ( .A1(n558), .A2(KEYINPUT101), .ZN(n555) );
  NAND2_X1 U574 ( .A1(n550), .A2(n549), .ZN(n548) );
  OR2_X1 U575 ( .A1(n531), .A2(KEYINPUT101), .ZN(n549) );
  NAND2_X1 U576 ( .A1(n551), .A2(n531), .ZN(n550) );
  NAND2_X1 U577 ( .A1(n553), .A2(n552), .ZN(n551) );
  INV_X1 U578 ( .A(KEYINPUT84), .ZN(n544) );
  NOR2_X1 U579 ( .A1(n1013), .A2(n746), .ZN(n747) );
  INV_X1 U580 ( .A(KEYINPUT93), .ZN(n717) );
  XNOR2_X1 U581 ( .A(KEYINPUT31), .B(KEYINPUT96), .ZN(n730) );
  XNOR2_X1 U582 ( .A(KEYINPUT32), .B(KEYINPUT97), .ZN(n775) );
  INV_X1 U583 ( .A(n558), .ZN(n553) );
  INV_X1 U584 ( .A(G40), .ZN(n543) );
  NOR2_X1 U585 ( .A1(G2105), .A2(G2104), .ZN(n561) );
  NAND2_X1 U586 ( .A1(n546), .A2(n532), .ZN(n545) );
  NOR2_X1 U587 ( .A1(n527), .A2(n530), .ZN(n537) );
  OR2_X1 U588 ( .A1(n567), .A2(n544), .ZN(n539) );
  NOR2_X1 U589 ( .A1(n578), .A2(n577), .ZN(G160) );
  AND2_X1 U590 ( .A1(n568), .A2(n544), .ZN(n527) );
  NAND2_X1 U591 ( .A1(n542), .A2(n529), .ZN(n820) );
  AND2_X1 U592 ( .A1(n796), .A2(n795), .ZN(n528) );
  NOR2_X1 U593 ( .A1(n577), .A2(n543), .ZN(n529) );
  AND2_X1 U594 ( .A1(n567), .A2(n544), .ZN(n530) );
  NOR2_X1 U595 ( .A1(n840), .A2(n844), .ZN(n531) );
  AND2_X1 U596 ( .A1(n531), .A2(n552), .ZN(n532) );
  NOR2_X1 U597 ( .A1(G164), .A2(G1384), .ZN(n533) );
  NAND2_X1 U598 ( .A1(n534), .A2(n1007), .ZN(n756) );
  NAND2_X1 U599 ( .A1(n536), .A2(n535), .ZN(n716) );
  NAND2_X2 U600 ( .A1(n537), .A2(n538), .ZN(G164) );
  OR2_X1 U601 ( .A1(n539), .A2(n568), .ZN(n538) );
  INV_X1 U602 ( .A(n578), .ZN(n542) );
  NAND2_X1 U603 ( .A1(n547), .A2(n545), .ZN(n556) );
  INV_X1 U604 ( .A(n559), .ZN(n546) );
  AND2_X1 U605 ( .A1(n554), .A2(n548), .ZN(n547) );
  NAND2_X1 U606 ( .A1(n559), .A2(n555), .ZN(n554) );
  NAND2_X1 U607 ( .A1(n556), .A2(n841), .ZN(n854) );
  AND2_X1 U608 ( .A1(G2105), .A2(G2104), .ZN(n914) );
  XNOR2_X1 U609 ( .A(n735), .B(KEYINPUT89), .ZN(n732) );
  OR2_X1 U610 ( .A1(n1018), .A2(n791), .ZN(n557) );
  XOR2_X1 U611 ( .A(n810), .B(KEYINPUT88), .Z(n558) );
  AND2_X1 U612 ( .A1(n806), .A2(n805), .ZN(n559) );
  INV_X1 U613 ( .A(G2104), .ZN(n564) );
  INV_X1 U614 ( .A(KEYINPUT89), .ZN(n734) );
  XNOR2_X1 U615 ( .A(n735), .B(n734), .ZN(n748) );
  INV_X1 U616 ( .A(KEYINPUT27), .ZN(n736) );
  INV_X1 U617 ( .A(KEYINPUT94), .ZN(n722) );
  INV_X1 U618 ( .A(n1021), .ZN(n793) );
  NOR2_X1 U619 ( .A1(n794), .A2(n793), .ZN(n795) );
  XNOR2_X1 U620 ( .A(n776), .B(n775), .ZN(n785) );
  INV_X1 U621 ( .A(KEYINPUT17), .ZN(n560) );
  AND2_X1 U622 ( .A1(n564), .A2(G2105), .ZN(n915) );
  NOR2_X1 U623 ( .A1(G651), .A2(n672), .ZN(n683) );
  XNOR2_X2 U624 ( .A(n561), .B(n560), .ZN(n911) );
  NAND2_X1 U625 ( .A1(G138), .A2(n911), .ZN(n563) );
  NAND2_X1 U626 ( .A1(G126), .A2(n915), .ZN(n562) );
  NAND2_X1 U627 ( .A1(n563), .A2(n562), .ZN(n568) );
  NAND2_X1 U628 ( .A1(G102), .A2(n569), .ZN(n566) );
  NAND2_X1 U629 ( .A1(G114), .A2(n914), .ZN(n565) );
  NAND2_X1 U630 ( .A1(n566), .A2(n565), .ZN(n567) );
  NAND2_X1 U631 ( .A1(G101), .A2(n569), .ZN(n570) );
  XNOR2_X1 U632 ( .A(n570), .B(KEYINPUT65), .ZN(n571) );
  XNOR2_X1 U633 ( .A(KEYINPUT23), .B(n571), .ZN(n574) );
  NAND2_X1 U634 ( .A1(G137), .A2(n911), .ZN(n572) );
  XNOR2_X1 U635 ( .A(n572), .B(KEYINPUT66), .ZN(n573) );
  NAND2_X1 U636 ( .A1(n574), .A2(n573), .ZN(n578) );
  NAND2_X1 U637 ( .A1(G113), .A2(n914), .ZN(n576) );
  NAND2_X1 U638 ( .A1(G125), .A2(n915), .ZN(n575) );
  NAND2_X1 U639 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U640 ( .A1(G651), .A2(G543), .ZN(n676) );
  NAND2_X1 U641 ( .A1(n676), .A2(G89), .ZN(n579) );
  XNOR2_X1 U642 ( .A(n579), .B(KEYINPUT4), .ZN(n581) );
  XOR2_X1 U643 ( .A(KEYINPUT0), .B(G543), .Z(n672) );
  INV_X1 U644 ( .A(G651), .ZN(n583) );
  NOR2_X1 U645 ( .A1(n672), .A2(n583), .ZN(n679) );
  NAND2_X1 U646 ( .A1(G76), .A2(n679), .ZN(n580) );
  NAND2_X1 U647 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n582), .B(KEYINPUT5), .ZN(n589) );
  NOR2_X1 U649 ( .A1(G543), .A2(n583), .ZN(n584) );
  XOR2_X1 U650 ( .A(KEYINPUT1), .B(n584), .Z(n675) );
  NAND2_X1 U651 ( .A1(G63), .A2(n675), .ZN(n586) );
  NAND2_X1 U652 ( .A1(G51), .A2(n683), .ZN(n585) );
  NAND2_X1 U653 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U654 ( .A(KEYINPUT6), .B(n587), .Z(n588) );
  NAND2_X1 U655 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U656 ( .A(n590), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U657 ( .A1(G72), .A2(n679), .ZN(n592) );
  NAND2_X1 U658 ( .A1(G85), .A2(n676), .ZN(n591) );
  NAND2_X1 U659 ( .A1(n592), .A2(n591), .ZN(n596) );
  NAND2_X1 U660 ( .A1(G60), .A2(n675), .ZN(n594) );
  NAND2_X1 U661 ( .A1(G47), .A2(n683), .ZN(n593) );
  NAND2_X1 U662 ( .A1(n594), .A2(n593), .ZN(n595) );
  OR2_X1 U663 ( .A1(n596), .A2(n595), .ZN(G290) );
  NAND2_X1 U664 ( .A1(n676), .A2(G90), .ZN(n597) );
  XNOR2_X1 U665 ( .A(n597), .B(KEYINPUT68), .ZN(n599) );
  NAND2_X1 U666 ( .A1(G77), .A2(n679), .ZN(n598) );
  NAND2_X1 U667 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U668 ( .A(n600), .B(KEYINPUT9), .ZN(n602) );
  NAND2_X1 U669 ( .A1(G64), .A2(n675), .ZN(n601) );
  NAND2_X1 U670 ( .A1(n602), .A2(n601), .ZN(n605) );
  NAND2_X1 U671 ( .A1(G52), .A2(n683), .ZN(n603) );
  XNOR2_X1 U672 ( .A(KEYINPUT67), .B(n603), .ZN(n604) );
  NOR2_X1 U673 ( .A1(n605), .A2(n604), .ZN(G171) );
  AND2_X1 U674 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U675 ( .A1(G123), .A2(n915), .ZN(n606) );
  XNOR2_X1 U676 ( .A(n606), .B(KEYINPUT18), .ZN(n613) );
  NAND2_X1 U677 ( .A1(G99), .A2(n569), .ZN(n608) );
  NAND2_X1 U678 ( .A1(G135), .A2(n911), .ZN(n607) );
  NAND2_X1 U679 ( .A1(n608), .A2(n607), .ZN(n611) );
  NAND2_X1 U680 ( .A1(n914), .A2(G111), .ZN(n609) );
  XOR2_X1 U681 ( .A(KEYINPUT74), .B(n609), .Z(n610) );
  NOR2_X1 U682 ( .A1(n611), .A2(n610), .ZN(n612) );
  NAND2_X1 U683 ( .A1(n613), .A2(n612), .ZN(n956) );
  XNOR2_X1 U684 ( .A(G2096), .B(n956), .ZN(n614) );
  OR2_X1 U685 ( .A1(G2100), .A2(n614), .ZN(G156) );
  INV_X1 U686 ( .A(G132), .ZN(G219) );
  INV_X1 U687 ( .A(G82), .ZN(G220) );
  INV_X1 U688 ( .A(G57), .ZN(G237) );
  NAND2_X1 U689 ( .A1(G88), .A2(n676), .ZN(n615) );
  XNOR2_X1 U690 ( .A(n615), .B(KEYINPUT76), .ZN(n617) );
  NAND2_X1 U691 ( .A1(n675), .A2(G62), .ZN(n616) );
  NAND2_X1 U692 ( .A1(n617), .A2(n616), .ZN(n621) );
  NAND2_X1 U693 ( .A1(G75), .A2(n679), .ZN(n619) );
  NAND2_X1 U694 ( .A1(G50), .A2(n683), .ZN(n618) );
  NAND2_X1 U695 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U696 ( .A1(n621), .A2(n620), .ZN(G166) );
  XOR2_X1 U697 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U698 ( .A1(G7), .A2(G661), .ZN(n622) );
  XNOR2_X1 U699 ( .A(n622), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U700 ( .A(G223), .ZN(n856) );
  NAND2_X1 U701 ( .A1(n856), .A2(G567), .ZN(n623) );
  XOR2_X1 U702 ( .A(KEYINPUT11), .B(n623), .Z(G234) );
  NAND2_X1 U703 ( .A1(n675), .A2(G56), .ZN(n624) );
  XNOR2_X1 U704 ( .A(n624), .B(KEYINPUT14), .ZN(n632) );
  NAND2_X1 U705 ( .A1(G68), .A2(n679), .ZN(n628) );
  XOR2_X1 U706 ( .A(KEYINPUT12), .B(KEYINPUT69), .Z(n626) );
  NAND2_X1 U707 ( .A1(G81), .A2(n676), .ZN(n625) );
  XNOR2_X1 U708 ( .A(n626), .B(n625), .ZN(n627) );
  NAND2_X1 U709 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U710 ( .A(n629), .B(KEYINPUT13), .ZN(n630) );
  XNOR2_X1 U711 ( .A(KEYINPUT70), .B(n630), .ZN(n631) );
  NAND2_X1 U712 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U713 ( .A(n633), .B(KEYINPUT71), .ZN(n635) );
  NAND2_X1 U714 ( .A1(G43), .A2(n683), .ZN(n634) );
  NAND2_X1 U715 ( .A1(n635), .A2(n634), .ZN(n1013) );
  INV_X1 U716 ( .A(G860), .ZN(n654) );
  OR2_X1 U717 ( .A1(n1013), .A2(n654), .ZN(G153) );
  XOR2_X1 U718 ( .A(G171), .B(KEYINPUT72), .Z(G301) );
  NAND2_X1 U719 ( .A1(G868), .A2(G301), .ZN(n645) );
  NAND2_X1 U720 ( .A1(G66), .A2(n675), .ZN(n637) );
  NAND2_X1 U721 ( .A1(G79), .A2(n679), .ZN(n636) );
  NAND2_X1 U722 ( .A1(n637), .A2(n636), .ZN(n641) );
  NAND2_X1 U723 ( .A1(G92), .A2(n676), .ZN(n639) );
  NAND2_X1 U724 ( .A1(G54), .A2(n683), .ZN(n638) );
  NAND2_X1 U725 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U726 ( .A1(n641), .A2(n640), .ZN(n643) );
  XNOR2_X1 U727 ( .A(KEYINPUT73), .B(KEYINPUT15), .ZN(n642) );
  XNOR2_X1 U728 ( .A(n643), .B(n642), .ZN(n1008) );
  OR2_X1 U729 ( .A1(n1008), .A2(G868), .ZN(n644) );
  NAND2_X1 U730 ( .A1(n645), .A2(n644), .ZN(G284) );
  NAND2_X1 U731 ( .A1(G65), .A2(n675), .ZN(n647) );
  NAND2_X1 U732 ( .A1(G53), .A2(n683), .ZN(n646) );
  NAND2_X1 U733 ( .A1(n647), .A2(n646), .ZN(n651) );
  NAND2_X1 U734 ( .A1(G78), .A2(n679), .ZN(n649) );
  NAND2_X1 U735 ( .A1(G91), .A2(n676), .ZN(n648) );
  NAND2_X1 U736 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U737 ( .A1(n651), .A2(n650), .ZN(n1007) );
  INV_X1 U738 ( .A(n1007), .ZN(G299) );
  INV_X1 U739 ( .A(G868), .ZN(n686) );
  NOR2_X1 U740 ( .A1(G286), .A2(n686), .ZN(n653) );
  NOR2_X1 U741 ( .A1(G868), .A2(G299), .ZN(n652) );
  NOR2_X1 U742 ( .A1(n653), .A2(n652), .ZN(G297) );
  NAND2_X1 U743 ( .A1(n654), .A2(G559), .ZN(n655) );
  NAND2_X1 U744 ( .A1(n655), .A2(n1008), .ZN(n656) );
  XNOR2_X1 U745 ( .A(n656), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U746 ( .A1(G868), .A2(n1013), .ZN(n659) );
  NAND2_X1 U747 ( .A1(n1008), .A2(G868), .ZN(n657) );
  NOR2_X1 U748 ( .A1(G559), .A2(n657), .ZN(n658) );
  NOR2_X1 U749 ( .A1(n659), .A2(n658), .ZN(G282) );
  NAND2_X1 U750 ( .A1(G67), .A2(n675), .ZN(n661) );
  NAND2_X1 U751 ( .A1(G80), .A2(n679), .ZN(n660) );
  NAND2_X1 U752 ( .A1(n661), .A2(n660), .ZN(n664) );
  NAND2_X1 U753 ( .A1(G93), .A2(n676), .ZN(n662) );
  XNOR2_X1 U754 ( .A(KEYINPUT75), .B(n662), .ZN(n663) );
  NOR2_X1 U755 ( .A1(n664), .A2(n663), .ZN(n666) );
  NAND2_X1 U756 ( .A1(n683), .A2(G55), .ZN(n665) );
  NAND2_X1 U757 ( .A1(n666), .A2(n665), .ZN(n694) );
  NAND2_X1 U758 ( .A1(G559), .A2(n1008), .ZN(n667) );
  XNOR2_X1 U759 ( .A(n667), .B(n1013), .ZN(n697) );
  NOR2_X1 U760 ( .A1(G860), .A2(n697), .ZN(n668) );
  XOR2_X1 U761 ( .A(n694), .B(n668), .Z(G145) );
  NAND2_X1 U762 ( .A1(G49), .A2(n683), .ZN(n670) );
  NAND2_X1 U763 ( .A1(G74), .A2(G651), .ZN(n669) );
  NAND2_X1 U764 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U765 ( .A1(n675), .A2(n671), .ZN(n674) );
  NAND2_X1 U766 ( .A1(n672), .A2(G87), .ZN(n673) );
  NAND2_X1 U767 ( .A1(n674), .A2(n673), .ZN(G288) );
  NAND2_X1 U768 ( .A1(G61), .A2(n675), .ZN(n678) );
  NAND2_X1 U769 ( .A1(G86), .A2(n676), .ZN(n677) );
  NAND2_X1 U770 ( .A1(n678), .A2(n677), .ZN(n682) );
  NAND2_X1 U771 ( .A1(n679), .A2(G73), .ZN(n680) );
  XOR2_X1 U772 ( .A(KEYINPUT2), .B(n680), .Z(n681) );
  NOR2_X1 U773 ( .A1(n682), .A2(n681), .ZN(n685) );
  NAND2_X1 U774 ( .A1(n683), .A2(G48), .ZN(n684) );
  NAND2_X1 U775 ( .A1(n685), .A2(n684), .ZN(G305) );
  NAND2_X1 U776 ( .A1(n686), .A2(n694), .ZN(n687) );
  XNOR2_X1 U777 ( .A(n687), .B(KEYINPUT80), .ZN(n700) );
  XOR2_X1 U778 ( .A(KEYINPUT78), .B(KEYINPUT77), .Z(n689) );
  XNOR2_X1 U779 ( .A(KEYINPUT19), .B(KEYINPUT79), .ZN(n688) );
  XNOR2_X1 U780 ( .A(n689), .B(n688), .ZN(n690) );
  XNOR2_X1 U781 ( .A(n1007), .B(n690), .ZN(n692) );
  XNOR2_X1 U782 ( .A(G288), .B(G166), .ZN(n691) );
  XNOR2_X1 U783 ( .A(n692), .B(n691), .ZN(n693) );
  XNOR2_X1 U784 ( .A(n693), .B(G290), .ZN(n695) );
  XNOR2_X1 U785 ( .A(n695), .B(n694), .ZN(n696) );
  XNOR2_X1 U786 ( .A(n696), .B(G305), .ZN(n929) );
  XNOR2_X1 U787 ( .A(n929), .B(n697), .ZN(n698) );
  NAND2_X1 U788 ( .A1(G868), .A2(n698), .ZN(n699) );
  NAND2_X1 U789 ( .A1(n700), .A2(n699), .ZN(G295) );
  NAND2_X1 U790 ( .A1(G2078), .A2(G2084), .ZN(n701) );
  XOR2_X1 U791 ( .A(KEYINPUT20), .B(n701), .Z(n702) );
  NAND2_X1 U792 ( .A1(G2090), .A2(n702), .ZN(n704) );
  XOR2_X1 U793 ( .A(KEYINPUT81), .B(KEYINPUT21), .Z(n703) );
  XNOR2_X1 U794 ( .A(n704), .B(n703), .ZN(n705) );
  NAND2_X1 U795 ( .A1(G2072), .A2(n705), .ZN(G158) );
  XNOR2_X1 U796 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U797 ( .A1(G120), .A2(G69), .ZN(n706) );
  NOR2_X1 U798 ( .A1(G237), .A2(n706), .ZN(n707) );
  XNOR2_X1 U799 ( .A(KEYINPUT82), .B(n707), .ZN(n708) );
  NAND2_X1 U800 ( .A1(n708), .A2(G108), .ZN(n860) );
  NAND2_X1 U801 ( .A1(n860), .A2(G567), .ZN(n713) );
  NOR2_X1 U802 ( .A1(G220), .A2(G219), .ZN(n709) );
  XOR2_X1 U803 ( .A(KEYINPUT22), .B(n709), .Z(n710) );
  NOR2_X1 U804 ( .A1(G218), .A2(n710), .ZN(n711) );
  NAND2_X1 U805 ( .A1(G96), .A2(n711), .ZN(n861) );
  NAND2_X1 U806 ( .A1(n861), .A2(G2106), .ZN(n712) );
  NAND2_X1 U807 ( .A1(n713), .A2(n712), .ZN(n885) );
  NAND2_X1 U808 ( .A1(G661), .A2(G483), .ZN(n714) );
  XOR2_X1 U809 ( .A(KEYINPUT83), .B(n714), .Z(n715) );
  NOR2_X1 U810 ( .A1(n885), .A2(n715), .ZN(n859) );
  NAND2_X1 U811 ( .A1(n859), .A2(G36), .ZN(G176) );
  INV_X1 U812 ( .A(G166), .ZN(G303) );
  NAND2_X1 U813 ( .A1(n742), .A2(G8), .ZN(n809) );
  NOR2_X1 U814 ( .A1(G1966), .A2(n809), .ZN(n782) );
  NOR2_X1 U815 ( .A1(n742), .A2(G2084), .ZN(n779) );
  NOR2_X1 U816 ( .A1(n782), .A2(n779), .ZN(n718) );
  XNOR2_X1 U817 ( .A(n718), .B(n717), .ZN(n719) );
  NAND2_X1 U818 ( .A1(n719), .A2(G8), .ZN(n720) );
  XNOR2_X1 U819 ( .A(KEYINPUT30), .B(n720), .ZN(n721) );
  XNOR2_X1 U820 ( .A(n723), .B(n722), .ZN(n729) );
  INV_X1 U821 ( .A(n742), .ZN(n735) );
  XOR2_X1 U822 ( .A(KEYINPUT25), .B(G2078), .Z(n987) );
  NOR2_X1 U823 ( .A1(n732), .A2(n987), .ZN(n725) );
  NOR2_X1 U824 ( .A1(G1961), .A2(n735), .ZN(n724) );
  NOR2_X1 U825 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U826 ( .A(KEYINPUT90), .B(n726), .Z(n761) );
  NOR2_X1 U827 ( .A1(G171), .A2(n761), .ZN(n727) );
  XNOR2_X1 U828 ( .A(KEYINPUT95), .B(n727), .ZN(n728) );
  NAND2_X1 U829 ( .A1(n729), .A2(n728), .ZN(n731) );
  NAND2_X1 U830 ( .A1(n732), .A2(G1956), .ZN(n733) );
  XNOR2_X1 U831 ( .A(KEYINPUT92), .B(n733), .ZN(n739) );
  NAND2_X1 U832 ( .A1(n748), .A2(G2072), .ZN(n737) );
  XNOR2_X1 U833 ( .A(n737), .B(n736), .ZN(n738) );
  INV_X1 U834 ( .A(KEYINPUT28), .ZN(n740) );
  XNOR2_X1 U835 ( .A(n741), .B(n740), .ZN(n758) );
  INV_X1 U836 ( .A(G1996), .ZN(n983) );
  NOR2_X1 U837 ( .A1(n526), .A2(n983), .ZN(n743) );
  XOR2_X1 U838 ( .A(n743), .B(KEYINPUT26), .Z(n745) );
  NAND2_X1 U839 ( .A1(n526), .A2(G1341), .ZN(n744) );
  NAND2_X1 U840 ( .A1(n745), .A2(n744), .ZN(n746) );
  OR2_X1 U841 ( .A1(n1008), .A2(n747), .ZN(n754) );
  NAND2_X1 U842 ( .A1(n1008), .A2(n747), .ZN(n752) );
  NAND2_X1 U843 ( .A1(G1348), .A2(n526), .ZN(n750) );
  NAND2_X1 U844 ( .A1(G2067), .A2(n748), .ZN(n749) );
  NAND2_X1 U845 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U846 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U847 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U848 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U849 ( .A1(n758), .A2(n757), .ZN(n760) );
  INV_X1 U850 ( .A(KEYINPUT29), .ZN(n759) );
  XNOR2_X1 U851 ( .A(n760), .B(n759), .ZN(n764) );
  NAND2_X1 U852 ( .A1(G171), .A2(n761), .ZN(n762) );
  XOR2_X1 U853 ( .A(KEYINPUT91), .B(n762), .Z(n763) );
  NAND2_X1 U854 ( .A1(n764), .A2(n763), .ZN(n777) );
  INV_X1 U855 ( .A(G8), .ZN(n769) );
  NOR2_X1 U856 ( .A1(n526), .A2(G2090), .ZN(n766) );
  NOR2_X1 U857 ( .A1(G1971), .A2(n809), .ZN(n765) );
  NOR2_X1 U858 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U859 ( .A1(n767), .A2(G303), .ZN(n768) );
  OR2_X1 U860 ( .A1(n769), .A2(n768), .ZN(n771) );
  AND2_X1 U861 ( .A1(n777), .A2(n771), .ZN(n770) );
  NAND2_X1 U862 ( .A1(n778), .A2(n770), .ZN(n774) );
  INV_X1 U863 ( .A(n771), .ZN(n772) );
  OR2_X1 U864 ( .A1(n772), .A2(G286), .ZN(n773) );
  NAND2_X1 U865 ( .A1(n774), .A2(n773), .ZN(n776) );
  NAND2_X1 U866 ( .A1(n778), .A2(n777), .ZN(n781) );
  NAND2_X1 U867 ( .A1(G8), .A2(n779), .ZN(n780) );
  NAND2_X1 U868 ( .A1(n781), .A2(n780), .ZN(n783) );
  NOR2_X1 U869 ( .A1(n783), .A2(n782), .ZN(n784) );
  NOR2_X1 U870 ( .A1(n785), .A2(n784), .ZN(n792) );
  NAND2_X1 U871 ( .A1(G166), .A2(G8), .ZN(n786) );
  NOR2_X1 U872 ( .A1(G2090), .A2(n786), .ZN(n787) );
  NOR2_X1 U873 ( .A1(n792), .A2(n787), .ZN(n788) );
  XNOR2_X1 U874 ( .A(n788), .B(KEYINPUT99), .ZN(n789) );
  NAND2_X1 U875 ( .A1(n789), .A2(n809), .ZN(n790) );
  XNOR2_X1 U876 ( .A(n790), .B(KEYINPUT100), .ZN(n806) );
  NOR2_X1 U877 ( .A1(G1976), .A2(G288), .ZN(n1018) );
  NOR2_X1 U878 ( .A1(G1971), .A2(G303), .ZN(n791) );
  OR2_X2 U879 ( .A1(n792), .A2(n557), .ZN(n796) );
  INV_X1 U880 ( .A(KEYINPUT98), .ZN(n797) );
  OR2_X1 U881 ( .A1(n809), .A2(n797), .ZN(n794) );
  NAND2_X1 U882 ( .A1(G1976), .A2(G288), .ZN(n1021) );
  NAND2_X1 U883 ( .A1(n797), .A2(n1018), .ZN(n800) );
  NAND2_X1 U884 ( .A1(n1018), .A2(KEYINPUT33), .ZN(n798) );
  NAND2_X1 U885 ( .A1(n798), .A2(KEYINPUT98), .ZN(n799) );
  NAND2_X1 U886 ( .A1(n800), .A2(n799), .ZN(n801) );
  NOR2_X1 U887 ( .A1(n809), .A2(n801), .ZN(n802) );
  NOR2_X1 U888 ( .A1(n803), .A2(n802), .ZN(n804) );
  XOR2_X1 U889 ( .A(G1981), .B(G305), .Z(n1004) );
  NAND2_X1 U890 ( .A1(n804), .A2(n1004), .ZN(n805) );
  NOR2_X1 U891 ( .A1(G1981), .A2(G305), .ZN(n807) );
  XOR2_X1 U892 ( .A(n807), .B(KEYINPUT24), .Z(n808) );
  NOR2_X1 U893 ( .A1(n809), .A2(n808), .ZN(n810) );
  XNOR2_X1 U894 ( .A(G2067), .B(KEYINPUT37), .ZN(n849) );
  NAND2_X1 U895 ( .A1(G104), .A2(n569), .ZN(n812) );
  NAND2_X1 U896 ( .A1(G140), .A2(n911), .ZN(n811) );
  NAND2_X1 U897 ( .A1(n812), .A2(n811), .ZN(n813) );
  XNOR2_X1 U898 ( .A(KEYINPUT34), .B(n813), .ZN(n818) );
  NAND2_X1 U899 ( .A1(G116), .A2(n914), .ZN(n815) );
  NAND2_X1 U900 ( .A1(G128), .A2(n915), .ZN(n814) );
  NAND2_X1 U901 ( .A1(n815), .A2(n814), .ZN(n816) );
  XOR2_X1 U902 ( .A(KEYINPUT35), .B(n816), .Z(n817) );
  NOR2_X1 U903 ( .A1(n818), .A2(n817), .ZN(n819) );
  XNOR2_X1 U904 ( .A(KEYINPUT36), .B(n819), .ZN(n926) );
  NOR2_X1 U905 ( .A1(n849), .A2(n926), .ZN(n962) );
  NOR2_X1 U906 ( .A1(n533), .A2(n820), .ZN(n851) );
  NAND2_X1 U907 ( .A1(n962), .A2(n851), .ZN(n821) );
  XOR2_X1 U908 ( .A(KEYINPUT85), .B(n821), .Z(n847) );
  INV_X1 U909 ( .A(n847), .ZN(n840) );
  NAND2_X1 U910 ( .A1(n911), .A2(G131), .ZN(n828) );
  NAND2_X1 U911 ( .A1(G107), .A2(n914), .ZN(n823) );
  NAND2_X1 U912 ( .A1(G95), .A2(n569), .ZN(n822) );
  NAND2_X1 U913 ( .A1(n823), .A2(n822), .ZN(n826) );
  NAND2_X1 U914 ( .A1(n915), .A2(G119), .ZN(n824) );
  XOR2_X1 U915 ( .A(KEYINPUT86), .B(n824), .Z(n825) );
  NOR2_X1 U916 ( .A1(n826), .A2(n825), .ZN(n827) );
  NAND2_X1 U917 ( .A1(n828), .A2(n827), .ZN(n829) );
  XOR2_X1 U918 ( .A(KEYINPUT87), .B(n829), .Z(n923) );
  AND2_X1 U919 ( .A1(n923), .A2(G1991), .ZN(n838) );
  NAND2_X1 U920 ( .A1(G117), .A2(n914), .ZN(n831) );
  NAND2_X1 U921 ( .A1(G141), .A2(n911), .ZN(n830) );
  NAND2_X1 U922 ( .A1(n831), .A2(n830), .ZN(n834) );
  NAND2_X1 U923 ( .A1(n569), .A2(G105), .ZN(n832) );
  XOR2_X1 U924 ( .A(KEYINPUT38), .B(n832), .Z(n833) );
  NOR2_X1 U925 ( .A1(n834), .A2(n833), .ZN(n836) );
  NAND2_X1 U926 ( .A1(n915), .A2(G129), .ZN(n835) );
  NAND2_X1 U927 ( .A1(n836), .A2(n835), .ZN(n895) );
  AND2_X1 U928 ( .A1(G1996), .A2(n895), .ZN(n837) );
  NOR2_X1 U929 ( .A1(n838), .A2(n837), .ZN(n970) );
  INV_X1 U930 ( .A(n851), .ZN(n839) );
  NOR2_X1 U931 ( .A1(n970), .A2(n839), .ZN(n844) );
  XNOR2_X1 U932 ( .A(G1986), .B(G290), .ZN(n1012) );
  NAND2_X1 U933 ( .A1(n1012), .A2(n851), .ZN(n841) );
  NOR2_X1 U934 ( .A1(G1996), .A2(n895), .ZN(n965) );
  NOR2_X1 U935 ( .A1(G1986), .A2(G290), .ZN(n842) );
  NOR2_X1 U936 ( .A1(G1991), .A2(n923), .ZN(n959) );
  NOR2_X1 U937 ( .A1(n842), .A2(n959), .ZN(n843) );
  NOR2_X1 U938 ( .A1(n844), .A2(n843), .ZN(n845) );
  NOR2_X1 U939 ( .A1(n965), .A2(n845), .ZN(n846) );
  XNOR2_X1 U940 ( .A(KEYINPUT39), .B(n846), .ZN(n848) );
  NAND2_X1 U941 ( .A1(n848), .A2(n847), .ZN(n850) );
  NAND2_X1 U942 ( .A1(n849), .A2(n926), .ZN(n972) );
  NAND2_X1 U943 ( .A1(n850), .A2(n972), .ZN(n852) );
  NAND2_X1 U944 ( .A1(n852), .A2(n851), .ZN(n853) );
  NAND2_X1 U945 ( .A1(n854), .A2(n853), .ZN(n855) );
  XNOR2_X1 U946 ( .A(KEYINPUT40), .B(n855), .ZN(G329) );
  NAND2_X1 U947 ( .A1(G2106), .A2(n856), .ZN(G217) );
  AND2_X1 U948 ( .A1(G15), .A2(G2), .ZN(n857) );
  NAND2_X1 U949 ( .A1(G661), .A2(n857), .ZN(G259) );
  NAND2_X1 U950 ( .A1(G3), .A2(G1), .ZN(n858) );
  NAND2_X1 U951 ( .A1(n859), .A2(n858), .ZN(G188) );
  INV_X1 U953 ( .A(G120), .ZN(G236) );
  INV_X1 U954 ( .A(G108), .ZN(G238) );
  INV_X1 U955 ( .A(G96), .ZN(G221) );
  INV_X1 U956 ( .A(G69), .ZN(G235) );
  NOR2_X1 U957 ( .A1(n861), .A2(n860), .ZN(G325) );
  INV_X1 U958 ( .A(G325), .ZN(G261) );
  XOR2_X1 U959 ( .A(G1966), .B(G1971), .Z(n863) );
  XNOR2_X1 U960 ( .A(G1981), .B(G1976), .ZN(n862) );
  XNOR2_X1 U961 ( .A(n863), .B(n862), .ZN(n876) );
  XOR2_X1 U962 ( .A(KEYINPUT104), .B(KEYINPUT103), .Z(n865) );
  XNOR2_X1 U963 ( .A(G1996), .B(G1991), .ZN(n864) );
  XNOR2_X1 U964 ( .A(n865), .B(n864), .ZN(n866) );
  XOR2_X1 U965 ( .A(n866), .B(KEYINPUT108), .Z(n874) );
  XOR2_X1 U966 ( .A(G2474), .B(G1956), .Z(n868) );
  XNOR2_X1 U967 ( .A(G1986), .B(G1961), .ZN(n867) );
  XNOR2_X1 U968 ( .A(n868), .B(n867), .ZN(n872) );
  XOR2_X1 U969 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n870) );
  XNOR2_X1 U970 ( .A(KEYINPUT107), .B(KEYINPUT41), .ZN(n869) );
  XNOR2_X1 U971 ( .A(n870), .B(n869), .ZN(n871) );
  XNOR2_X1 U972 ( .A(n872), .B(n871), .ZN(n873) );
  XNOR2_X1 U973 ( .A(n874), .B(n873), .ZN(n875) );
  XOR2_X1 U974 ( .A(n876), .B(n875), .Z(G229) );
  XOR2_X1 U975 ( .A(G2100), .B(G2096), .Z(n878) );
  XNOR2_X1 U976 ( .A(KEYINPUT42), .B(G2678), .ZN(n877) );
  XNOR2_X1 U977 ( .A(n878), .B(n877), .ZN(n882) );
  XOR2_X1 U978 ( .A(KEYINPUT43), .B(G2090), .Z(n880) );
  XNOR2_X1 U979 ( .A(G2067), .B(G2072), .ZN(n879) );
  XNOR2_X1 U980 ( .A(n880), .B(n879), .ZN(n881) );
  XOR2_X1 U981 ( .A(n882), .B(n881), .Z(n884) );
  XNOR2_X1 U982 ( .A(G2078), .B(G2084), .ZN(n883) );
  XNOR2_X1 U983 ( .A(n884), .B(n883), .ZN(G227) );
  INV_X1 U984 ( .A(n885), .ZN(G319) );
  NAND2_X1 U985 ( .A1(G112), .A2(n914), .ZN(n887) );
  NAND2_X1 U986 ( .A1(G100), .A2(n569), .ZN(n886) );
  NAND2_X1 U987 ( .A1(n887), .A2(n886), .ZN(n888) );
  XNOR2_X1 U988 ( .A(KEYINPUT110), .B(n888), .ZN(n894) );
  NAND2_X1 U989 ( .A1(G124), .A2(n915), .ZN(n889) );
  XOR2_X1 U990 ( .A(KEYINPUT44), .B(n889), .Z(n890) );
  XNOR2_X1 U991 ( .A(n890), .B(KEYINPUT109), .ZN(n892) );
  NAND2_X1 U992 ( .A1(G136), .A2(n911), .ZN(n891) );
  NAND2_X1 U993 ( .A1(n892), .A2(n891), .ZN(n893) );
  NOR2_X1 U994 ( .A1(n894), .A2(n893), .ZN(G162) );
  XOR2_X1 U995 ( .A(n895), .B(G162), .Z(n897) );
  XNOR2_X1 U996 ( .A(G160), .B(G164), .ZN(n896) );
  XNOR2_X1 U997 ( .A(n897), .B(n896), .ZN(n910) );
  XNOR2_X1 U998 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n908) );
  NAND2_X1 U999 ( .A1(G118), .A2(n914), .ZN(n899) );
  NAND2_X1 U1000 ( .A1(G130), .A2(n915), .ZN(n898) );
  NAND2_X1 U1001 ( .A1(n899), .A2(n898), .ZN(n905) );
  NAND2_X1 U1002 ( .A1(G106), .A2(n569), .ZN(n901) );
  NAND2_X1 U1003 ( .A1(G142), .A2(n911), .ZN(n900) );
  NAND2_X1 U1004 ( .A1(n901), .A2(n900), .ZN(n902) );
  XNOR2_X1 U1005 ( .A(KEYINPUT45), .B(n902), .ZN(n903) );
  XNOR2_X1 U1006 ( .A(KEYINPUT111), .B(n903), .ZN(n904) );
  NOR2_X1 U1007 ( .A1(n905), .A2(n904), .ZN(n906) );
  XNOR2_X1 U1008 ( .A(n956), .B(n906), .ZN(n907) );
  XNOR2_X1 U1009 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1010 ( .A(n910), .B(n909), .Z(n925) );
  NAND2_X1 U1011 ( .A1(G103), .A2(n569), .ZN(n913) );
  NAND2_X1 U1012 ( .A1(G139), .A2(n911), .ZN(n912) );
  NAND2_X1 U1013 ( .A1(n913), .A2(n912), .ZN(n921) );
  NAND2_X1 U1014 ( .A1(G115), .A2(n914), .ZN(n917) );
  NAND2_X1 U1015 ( .A1(G127), .A2(n915), .ZN(n916) );
  NAND2_X1 U1016 ( .A1(n917), .A2(n916), .ZN(n918) );
  XOR2_X1 U1017 ( .A(KEYINPUT47), .B(n918), .Z(n919) );
  XNOR2_X1 U1018 ( .A(KEYINPUT112), .B(n919), .ZN(n920) );
  NOR2_X1 U1019 ( .A1(n921), .A2(n920), .ZN(n922) );
  XOR2_X1 U1020 ( .A(KEYINPUT113), .B(n922), .Z(n951) );
  XOR2_X1 U1021 ( .A(n923), .B(n951), .Z(n924) );
  XNOR2_X1 U1022 ( .A(n925), .B(n924), .ZN(n927) );
  XNOR2_X1 U1023 ( .A(n927), .B(n926), .ZN(n928) );
  NOR2_X1 U1024 ( .A1(G37), .A2(n928), .ZN(G395) );
  XOR2_X1 U1025 ( .A(n929), .B(G286), .Z(n931) );
  XNOR2_X1 U1026 ( .A(G171), .B(n1008), .ZN(n930) );
  XNOR2_X1 U1027 ( .A(n931), .B(n930), .ZN(n932) );
  XNOR2_X1 U1028 ( .A(n932), .B(n1013), .ZN(n933) );
  NOR2_X1 U1029 ( .A1(G37), .A2(n933), .ZN(G397) );
  XNOR2_X1 U1030 ( .A(KEYINPUT49), .B(KEYINPUT114), .ZN(n935) );
  NOR2_X1 U1031 ( .A1(G229), .A2(G227), .ZN(n934) );
  XNOR2_X1 U1032 ( .A(n935), .B(n934), .ZN(n947) );
  XOR2_X1 U1033 ( .A(KEYINPUT102), .B(G2446), .Z(n937) );
  XNOR2_X1 U1034 ( .A(G2443), .B(G2454), .ZN(n936) );
  XNOR2_X1 U1035 ( .A(n937), .B(n936), .ZN(n938) );
  XOR2_X1 U1036 ( .A(n938), .B(G2451), .Z(n940) );
  XNOR2_X1 U1037 ( .A(G1341), .B(G1348), .ZN(n939) );
  XNOR2_X1 U1038 ( .A(n940), .B(n939), .ZN(n944) );
  XOR2_X1 U1039 ( .A(G2435), .B(G2427), .Z(n942) );
  XNOR2_X1 U1040 ( .A(G2430), .B(G2438), .ZN(n941) );
  XNOR2_X1 U1041 ( .A(n942), .B(n941), .ZN(n943) );
  XOR2_X1 U1042 ( .A(n944), .B(n943), .Z(n945) );
  NAND2_X1 U1043 ( .A1(G14), .A2(n945), .ZN(n950) );
  NAND2_X1 U1044 ( .A1(G319), .A2(n950), .ZN(n946) );
  NOR2_X1 U1045 ( .A1(n947), .A2(n946), .ZN(n949) );
  NOR2_X1 U1046 ( .A1(G395), .A2(G397), .ZN(n948) );
  NAND2_X1 U1047 ( .A1(n949), .A2(n948), .ZN(G225) );
  INV_X1 U1048 ( .A(G225), .ZN(G308) );
  INV_X1 U1049 ( .A(n950), .ZN(G401) );
  XNOR2_X1 U1050 ( .A(G164), .B(G2078), .ZN(n954) );
  XNOR2_X1 U1051 ( .A(G2072), .B(n951), .ZN(n952) );
  XNOR2_X1 U1052 ( .A(n952), .B(KEYINPUT118), .ZN(n953) );
  NAND2_X1 U1053 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1054 ( .A(n955), .B(KEYINPUT50), .ZN(n975) );
  XNOR2_X1 U1055 ( .A(G160), .B(G2084), .ZN(n957) );
  NAND2_X1 U1056 ( .A1(n957), .A2(n956), .ZN(n958) );
  NOR2_X1 U1057 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1058 ( .A(n960), .B(KEYINPUT115), .ZN(n961) );
  NOR2_X1 U1059 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1060 ( .A(KEYINPUT116), .B(n963), .Z(n968) );
  XOR2_X1 U1061 ( .A(G2090), .B(G162), .Z(n964) );
  NOR2_X1 U1062 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1063 ( .A(KEYINPUT51), .B(n966), .ZN(n967) );
  NOR2_X1 U1064 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1065 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1066 ( .A(n971), .B(KEYINPUT117), .ZN(n973) );
  NAND2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n974) );
  NOR2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1069 ( .A(KEYINPUT52), .B(n976), .ZN(n978) );
  INV_X1 U1070 ( .A(KEYINPUT55), .ZN(n977) );
  NAND2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1072 ( .A1(n979), .A2(G29), .ZN(n980) );
  XOR2_X1 U1073 ( .A(KEYINPUT119), .B(n980), .Z(n1059) );
  XOR2_X1 U1074 ( .A(G29), .B(KEYINPUT122), .Z(n1002) );
  XNOR2_X1 U1075 ( .A(G1991), .B(G25), .ZN(n992) );
  XNOR2_X1 U1076 ( .A(G2067), .B(G26), .ZN(n982) );
  XNOR2_X1 U1077 ( .A(G33), .B(G2072), .ZN(n981) );
  NOR2_X1 U1078 ( .A1(n982), .A2(n981), .ZN(n986) );
  XNOR2_X1 U1079 ( .A(G32), .B(KEYINPUT120), .ZN(n984) );
  XNOR2_X1 U1080 ( .A(n984), .B(n983), .ZN(n985) );
  NAND2_X1 U1081 ( .A1(n986), .A2(n985), .ZN(n989) );
  XNOR2_X1 U1082 ( .A(G27), .B(n987), .ZN(n988) );
  NOR2_X1 U1083 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1084 ( .A(KEYINPUT121), .B(n990), .ZN(n991) );
  NOR2_X1 U1085 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1086 ( .A1(G28), .A2(n993), .ZN(n994) );
  XNOR2_X1 U1087 ( .A(n994), .B(KEYINPUT53), .ZN(n997) );
  XOR2_X1 U1088 ( .A(G2084), .B(G34), .Z(n995) );
  XNOR2_X1 U1089 ( .A(KEYINPUT54), .B(n995), .ZN(n996) );
  NAND2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n999) );
  XNOR2_X1 U1091 ( .A(G35), .B(G2090), .ZN(n998) );
  NOR2_X1 U1092 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1093 ( .A(n1000), .B(KEYINPUT55), .ZN(n1001) );
  NAND2_X1 U1094 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1095 ( .A1(G11), .A2(n1003), .ZN(n1057) );
  XNOR2_X1 U1096 ( .A(G16), .B(KEYINPUT56), .ZN(n1030) );
  XNOR2_X1 U1097 ( .A(G1966), .B(G168), .ZN(n1005) );
  NAND2_X1 U1098 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1099 ( .A(KEYINPUT57), .B(n1006), .ZN(n1028) );
  XNOR2_X1 U1100 ( .A(n1007), .B(G1956), .ZN(n1010) );
  XNOR2_X1 U1101 ( .A(n1008), .B(G1348), .ZN(n1009) );
  NAND2_X1 U1102 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NOR2_X1 U1103 ( .A1(n1012), .A2(n1011), .ZN(n1017) );
  XOR2_X1 U1104 ( .A(G171), .B(G1961), .Z(n1015) );
  XNOR2_X1 U1105 ( .A(n1013), .B(G1341), .ZN(n1014) );
  NOR2_X1 U1106 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1107 ( .A1(n1017), .A2(n1016), .ZN(n1025) );
  XOR2_X1 U1108 ( .A(n1018), .B(KEYINPUT123), .Z(n1020) );
  XOR2_X1 U1109 ( .A(G1971), .B(G166), .Z(n1019) );
  NOR2_X1 U1110 ( .A1(n1020), .A2(n1019), .ZN(n1022) );
  NAND2_X1 U1111 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1112 ( .A(KEYINPUT124), .B(n1023), .ZN(n1024) );
  NOR2_X1 U1113 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1114 ( .A(KEYINPUT125), .B(n1026), .Z(n1027) );
  NAND2_X1 U1115 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1116 ( .A1(n1030), .A2(n1029), .ZN(n1055) );
  INV_X1 U1117 ( .A(G16), .ZN(n1053) );
  XNOR2_X1 U1118 ( .A(G1348), .B(KEYINPUT59), .ZN(n1031) );
  XNOR2_X1 U1119 ( .A(n1031), .B(G4), .ZN(n1035) );
  XNOR2_X1 U1120 ( .A(G1341), .B(G19), .ZN(n1033) );
  XNOR2_X1 U1121 ( .A(G1956), .B(G20), .ZN(n1032) );
  NOR2_X1 U1122 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NAND2_X1 U1123 ( .A1(n1035), .A2(n1034), .ZN(n1038) );
  XNOR2_X1 U1124 ( .A(KEYINPUT126), .B(G1981), .ZN(n1036) );
  XNOR2_X1 U1125 ( .A(G6), .B(n1036), .ZN(n1037) );
  NOR2_X1 U1126 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  XNOR2_X1 U1127 ( .A(KEYINPUT60), .B(n1039), .ZN(n1043) );
  XNOR2_X1 U1128 ( .A(G1966), .B(G21), .ZN(n1041) );
  XNOR2_X1 U1129 ( .A(G5), .B(G1961), .ZN(n1040) );
  NOR2_X1 U1130 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  NAND2_X1 U1131 ( .A1(n1043), .A2(n1042), .ZN(n1050) );
  XNOR2_X1 U1132 ( .A(G1976), .B(G23), .ZN(n1045) );
  XNOR2_X1 U1133 ( .A(G1971), .B(G22), .ZN(n1044) );
  NOR2_X1 U1134 ( .A1(n1045), .A2(n1044), .ZN(n1047) );
  XOR2_X1 U1135 ( .A(G1986), .B(G24), .Z(n1046) );
  NAND2_X1 U1136 ( .A1(n1047), .A2(n1046), .ZN(n1048) );
  XNOR2_X1 U1137 ( .A(KEYINPUT58), .B(n1048), .ZN(n1049) );
  NOR2_X1 U1138 ( .A1(n1050), .A2(n1049), .ZN(n1051) );
  XNOR2_X1 U1139 ( .A(KEYINPUT61), .B(n1051), .ZN(n1052) );
  NAND2_X1 U1140 ( .A1(n1053), .A2(n1052), .ZN(n1054) );
  NAND2_X1 U1141 ( .A1(n1055), .A2(n1054), .ZN(n1056) );
  NOR2_X1 U1142 ( .A1(n1057), .A2(n1056), .ZN(n1058) );
  NAND2_X1 U1143 ( .A1(n1059), .A2(n1058), .ZN(n1060) );
  XNOR2_X1 U1144 ( .A(n1060), .B(KEYINPUT62), .ZN(n1061) );
  XNOR2_X1 U1145 ( .A(KEYINPUT127), .B(n1061), .ZN(G311) );
  INV_X1 U1146 ( .A(G311), .ZN(G150) );
endmodule

