

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764;

  XNOR2_X1 U375 ( .A(n530), .B(n529), .ZN(n565) );
  AND2_X1 U376 ( .A1(n553), .A2(n711), .ZN(n530) );
  AND2_X1 U377 ( .A1(n399), .A2(n397), .ZN(n553) );
  NOR2_X1 U378 ( .A1(n590), .A2(n414), .ZN(n611) );
  INV_X1 U379 ( .A(n584), .ZN(n604) );
  BUF_X1 U380 ( .A(n598), .Z(n702) );
  NAND2_X1 U381 ( .A1(n697), .A2(n698), .ZN(n693) );
  XNOR2_X1 U382 ( .A(n542), .B(n541), .ZN(n572) );
  OR2_X1 U383 ( .A1(n627), .A2(n410), .ZN(n409) );
  BUF_X1 U384 ( .A(G143), .Z(n357) );
  XNOR2_X1 U385 ( .A(n511), .B(n446), .ZN(n499) );
  XNOR2_X1 U386 ( .A(n373), .B(G146), .ZN(n513) );
  INV_X1 U387 ( .A(G125), .ZN(n373) );
  INV_X2 U388 ( .A(G143), .ZN(n445) );
  XNOR2_X1 U389 ( .A(G101), .B(KEYINPUT3), .ZN(n394) );
  INV_X4 U390 ( .A(G953), .ZN(n749) );
  NOR2_X2 U391 ( .A1(n762), .A2(n764), .ZN(n369) );
  XNOR2_X2 U392 ( .A(n371), .B(n370), .ZN(n762) );
  NAND2_X1 U393 ( .A1(n356), .A2(n383), .ZN(n381) );
  NOR2_X1 U394 ( .A1(n428), .A2(n430), .ZN(n356) );
  XNOR2_X2 U395 ( .A(n499), .B(n435), .ZN(n747) );
  XNOR2_X1 U396 ( .A(G113), .B(n357), .ZN(n483) );
  XNOR2_X1 U397 ( .A(G119), .B(G128), .ZN(n461) );
  XNOR2_X2 U398 ( .A(n389), .B(n366), .ZN(n597) );
  AND2_X1 U399 ( .A1(n378), .A2(n614), .ZN(n387) );
  INV_X1 U400 ( .A(n548), .ZN(n677) );
  AND2_X1 U401 ( .A1(n553), .A2(n552), .ZN(n555) );
  NAND2_X1 U402 ( .A1(n407), .A2(n413), .ZN(n562) );
  NOR2_X1 U403 ( .A1(n537), .A2(n536), .ZN(n538) );
  AND2_X1 U404 ( .A1(n400), .A2(n527), .ZN(n399) );
  XNOR2_X1 U405 ( .A(n398), .B(n528), .ZN(n397) );
  NAND2_X1 U406 ( .A1(n711), .A2(n710), .ZN(n715) );
  AND2_X1 U407 ( .A1(n409), .A2(n412), .ZN(n407) );
  AND2_X1 U408 ( .A1(n409), .A2(n365), .ZN(n408) );
  XNOR2_X2 U409 ( .A(n747), .B(G146), .ZN(n469) );
  XNOR2_X1 U410 ( .A(n513), .B(n372), .ZN(n482) );
  INV_X1 U411 ( .A(KEYINPUT10), .ZN(n372) );
  XNOR2_X1 U412 ( .A(G113), .B(KEYINPUT72), .ZN(n438) );
  NAND2_X1 U413 ( .A1(n411), .A2(n517), .ZN(n410) );
  NAND2_X1 U414 ( .A1(n597), .A2(n360), .ZN(n379) );
  INV_X1 U415 ( .A(n639), .ZN(n401) );
  NAND2_X1 U416 ( .A1(n431), .A2(n426), .ZN(n425) );
  XNOR2_X1 U417 ( .A(n369), .B(n531), .ZN(n383) );
  XNOR2_X1 U418 ( .A(G137), .B(G116), .ZN(n442) );
  XOR2_X1 U419 ( .A(KEYINPUT5), .B(KEYINPUT89), .Z(n443) );
  XOR2_X1 U420 ( .A(G131), .B(KEYINPUT4), .Z(n435) );
  XNOR2_X1 U421 ( .A(G131), .B(KEYINPUT91), .ZN(n477) );
  XNOR2_X1 U422 ( .A(G137), .B(G140), .ZN(n470) );
  XNOR2_X1 U423 ( .A(G104), .B(KEYINPUT86), .ZN(n393) );
  XNOR2_X1 U424 ( .A(G101), .B(G110), .ZN(n471) );
  XNOR2_X1 U425 ( .A(n375), .B(n391), .ZN(n390) );
  INV_X1 U426 ( .A(KEYINPUT34), .ZN(n391) );
  INV_X1 U427 ( .A(G469), .ZN(n388) );
  XNOR2_X1 U428 ( .A(KEYINPUT85), .B(KEYINPUT4), .ZN(n512) );
  XNOR2_X1 U429 ( .A(n507), .B(n506), .ZN(n646) );
  INV_X1 U430 ( .A(KEYINPUT2), .ZN(n406) );
  NOR2_X1 U431 ( .A1(n741), .A2(G902), .ZN(n465) );
  XNOR2_X1 U432 ( .A(n491), .B(n490), .ZN(n576) );
  XNOR2_X1 U433 ( .A(n489), .B(G475), .ZN(n490) );
  NAND2_X1 U434 ( .A1(n385), .A2(n414), .ZN(n539) );
  XNOR2_X1 U435 ( .A(n386), .B(KEYINPUT36), .ZN(n385) );
  NOR2_X1 U436 ( .A1(n559), .A2(n562), .ZN(n386) );
  XNOR2_X1 U437 ( .A(n558), .B(n429), .ZN(n428) );
  INV_X1 U438 ( .A(KEYINPUT79), .ZN(n429) );
  XOR2_X1 U439 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n478) );
  INV_X1 U440 ( .A(G237), .ZN(n518) );
  INV_X1 U441 ( .A(G902), .ZN(n519) );
  INV_X1 U442 ( .A(G122), .ZN(n476) );
  NAND2_X1 U443 ( .A1(n619), .A2(KEYINPUT66), .ZN(n422) );
  NOR2_X1 U444 ( .A1(n377), .A2(n425), .ZN(n424) );
  NAND2_X1 U445 ( .A1(n520), .A2(n617), .ZN(n412) );
  XOR2_X1 U446 ( .A(KEYINPUT20), .B(KEYINPUT87), .Z(n449) );
  XNOR2_X1 U447 ( .A(n603), .B(n526), .ZN(n400) );
  NAND2_X1 U448 ( .A1(n591), .A2(n710), .ZN(n398) );
  XNOR2_X1 U449 ( .A(n441), .B(n396), .ZN(n395) );
  XNOR2_X1 U450 ( .A(n440), .B(n444), .ZN(n396) );
  XNOR2_X1 U451 ( .A(n461), .B(n460), .ZN(n462) );
  INV_X1 U452 ( .A(KEYINPUT23), .ZN(n460) );
  XOR2_X1 U453 ( .A(G110), .B(KEYINPUT24), .Z(n459) );
  XNOR2_X1 U454 ( .A(n458), .B(n433), .ZN(n492) );
  INV_X1 U455 ( .A(KEYINPUT8), .ZN(n433) );
  INV_X1 U456 ( .A(G134), .ZN(n446) );
  XOR2_X1 U457 ( .A(KEYINPUT95), .B(G122), .Z(n494) );
  XNOR2_X1 U458 ( .A(n488), .B(n487), .ZN(n651) );
  XNOR2_X1 U459 ( .A(n486), .B(n437), .ZN(n487) );
  XNOR2_X1 U460 ( .A(n474), .B(G107), .ZN(n427) );
  XNOR2_X1 U461 ( .A(n473), .B(n392), .ZN(n474) );
  XNOR2_X1 U462 ( .A(n470), .B(n393), .ZN(n392) );
  XNOR2_X1 U463 ( .A(n376), .B(n417), .ZN(n416) );
  NOR2_X1 U464 ( .A1(n599), .A2(n581), .ZN(n376) );
  INV_X1 U465 ( .A(n727), .ZN(n415) );
  NAND2_X1 U466 ( .A1(n390), .A2(n362), .ZN(n389) );
  XNOR2_X1 U467 ( .A(n745), .B(n463), .ZN(n741) );
  XNOR2_X1 U468 ( .A(n434), .B(n432), .ZN(n463) );
  NAND2_X1 U469 ( .A1(n492), .A2(G221), .ZN(n432) );
  XNOR2_X1 U470 ( .A(n462), .B(n459), .ZN(n434) );
  XNOR2_X1 U471 ( .A(n646), .B(n516), .ZN(n627) );
  AND2_X1 U472 ( .A1(n630), .A2(n754), .ZN(n744) );
  XNOR2_X1 U473 ( .A(n404), .B(n403), .ZN(n402) );
  INV_X1 U474 ( .A(KEYINPUT81), .ZN(n403) );
  NAND2_X1 U475 ( .A1(n405), .A2(n691), .ZN(n404) );
  BUF_X1 U476 ( .A(G953), .Z(n754) );
  INV_X1 U477 ( .A(KEYINPUT40), .ZN(n370) );
  INV_X1 U478 ( .A(n581), .ZN(n609) );
  INV_X1 U479 ( .A(n539), .ZN(n686) );
  XNOR2_X1 U480 ( .A(n532), .B(KEYINPUT1), .ZN(n694) );
  AND2_X1 U481 ( .A1(n596), .A2(KEYINPUT70), .ZN(n358) );
  XOR2_X1 U482 ( .A(KEYINPUT25), .B(n436), .Z(n359) );
  AND2_X1 U483 ( .A1(n401), .A2(n358), .ZN(n360) );
  OR2_X1 U484 ( .A1(n719), .A2(n718), .ZN(n361) );
  AND2_X1 U485 ( .A1(n576), .A2(n575), .ZN(n362) );
  XNOR2_X1 U486 ( .A(n598), .B(KEYINPUT99), .ZN(n591) );
  OR2_X1 U487 ( .A1(n548), .A2(n547), .ZN(n363) );
  OR2_X1 U488 ( .A1(n620), .A2(n690), .ZN(n364) );
  INV_X1 U489 ( .A(n694), .ZN(n414) );
  AND2_X1 U490 ( .A1(n710), .A2(n412), .ZN(n365) );
  XOR2_X1 U491 ( .A(KEYINPUT76), .B(KEYINPUT35), .Z(n366) );
  XNOR2_X1 U492 ( .A(n469), .B(n395), .ZN(n633) );
  XNOR2_X1 U493 ( .A(n469), .B(n427), .ZN(n657) );
  XNOR2_X1 U494 ( .A(KEYINPUT48), .B(KEYINPUT71), .ZN(n367) );
  NOR2_X1 U495 ( .A1(n581), .A2(n534), .ZN(n535) );
  INV_X1 U496 ( .A(n597), .ZN(n757) );
  NAND2_X1 U497 ( .A1(n615), .A2(n387), .ZN(n368) );
  XNOR2_X2 U498 ( .A(n368), .B(n616), .ZN(n620) );
  NAND2_X1 U499 ( .A1(n379), .A2(KEYINPUT44), .ZN(n378) );
  XOR2_X2 U500 ( .A(n521), .B(n562), .Z(n711) );
  NAND2_X1 U501 ( .A1(n565), .A2(n544), .ZN(n371) );
  XNOR2_X2 U502 ( .A(n374), .B(n388), .ZN(n532) );
  NAND2_X1 U503 ( .A1(n657), .A2(n519), .ZN(n374) );
  NAND2_X1 U504 ( .A1(n416), .A2(n604), .ZN(n375) );
  NAND2_X1 U505 ( .A1(n419), .A2(n377), .ZN(n418) );
  NOR2_X2 U506 ( .A1(n620), .A2(n517), .ZN(n377) );
  NAND2_X2 U507 ( .A1(n380), .A2(n566), .ZN(n621) );
  XNOR2_X2 U508 ( .A(n381), .B(n367), .ZN(n380) );
  XNOR2_X2 U509 ( .A(n384), .B(n447), .ZN(n598) );
  NAND2_X1 U510 ( .A1(n633), .A2(n519), .ZN(n384) );
  XNOR2_X2 U511 ( .A(n621), .B(n567), .ZN(n748) );
  XNOR2_X2 U512 ( .A(n702), .B(n533), .ZN(n581) );
  XNOR2_X1 U513 ( .A(n394), .B(G119), .ZN(n439) );
  NOR2_X2 U514 ( .A1(n532), .A2(n693), .ZN(n603) );
  AND2_X2 U515 ( .A1(n593), .A2(n608), .ZN(n639) );
  NAND2_X1 U516 ( .A1(n402), .A2(n732), .ZN(n733) );
  NAND2_X1 U517 ( .A1(n364), .A2(n406), .ZN(n405) );
  NAND2_X1 U518 ( .A1(n408), .A2(n413), .ZN(n542) );
  NAND2_X1 U519 ( .A1(n627), .A2(n520), .ZN(n413) );
  INV_X1 U520 ( .A(n520), .ZN(n411) );
  NAND2_X1 U521 ( .A1(n611), .A2(n467), .ZN(n592) );
  AND2_X1 U522 ( .A1(n416), .A2(n361), .ZN(n720) );
  AND2_X1 U523 ( .A1(n416), .A2(n415), .ZN(n728) );
  INV_X1 U524 ( .A(KEYINPUT33), .ZN(n417) );
  NAND2_X1 U525 ( .A1(n420), .A2(n418), .ZN(n624) );
  AND2_X1 U526 ( .A1(n748), .A2(KEYINPUT66), .ZN(n419) );
  NOR2_X1 U527 ( .A1(n424), .A2(n421), .ZN(n420) );
  NAND2_X1 U528 ( .A1(n423), .A2(n422), .ZN(n421) );
  OR2_X2 U529 ( .A1(n748), .A2(n425), .ZN(n423) );
  INV_X1 U530 ( .A(KEYINPUT66), .ZN(n426) );
  NAND2_X1 U531 ( .A1(n539), .A2(n363), .ZN(n430) );
  INV_X1 U532 ( .A(n619), .ZN(n431) );
  BUF_X1 U533 ( .A(n735), .Z(n740) );
  AND2_X1 U534 ( .A1(n464), .A2(G217), .ZN(n436) );
  AND2_X1 U535 ( .A1(G214), .A2(n485), .ZN(n437) );
  XNOR2_X1 U536 ( .A(n763), .B(KEYINPUT80), .ZN(n556) );
  INV_X1 U537 ( .A(KEYINPUT103), .ZN(n526) );
  INV_X1 U538 ( .A(KEYINPUT39), .ZN(n529) );
  INV_X1 U539 ( .A(KEYINPUT104), .ZN(n554) );
  XNOR2_X1 U540 ( .A(n439), .B(n438), .ZN(n506) );
  INV_X1 U541 ( .A(n506), .ZN(n441) );
  NOR2_X1 U542 ( .A1(n754), .A2(G237), .ZN(n485) );
  AND2_X1 U543 ( .A1(G210), .A2(n485), .ZN(n440) );
  XNOR2_X1 U544 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X2 U545 ( .A(n445), .B(G128), .ZN(n511) );
  INV_X1 U546 ( .A(G472), .ZN(n447) );
  INV_X1 U547 ( .A(n591), .ZN(n467) );
  XNOR2_X2 U548 ( .A(G902), .B(KEYINPUT15), .ZN(n517) );
  NAND2_X1 U549 ( .A1(G234), .A2(n517), .ZN(n448) );
  XNOR2_X1 U550 ( .A(n449), .B(n448), .ZN(n464) );
  AND2_X1 U551 ( .A1(n464), .A2(G221), .ZN(n451) );
  XNOR2_X1 U552 ( .A(KEYINPUT88), .B(KEYINPUT21), .ZN(n450) );
  XNOR2_X1 U553 ( .A(n451), .B(n450), .ZN(n698) );
  NAND2_X1 U554 ( .A1(G234), .A2(G237), .ZN(n452) );
  XNOR2_X1 U555 ( .A(n452), .B(KEYINPUT14), .ZN(n692) );
  INV_X1 U556 ( .A(G952), .ZN(n630) );
  NAND2_X1 U557 ( .A1(n749), .A2(n630), .ZN(n454) );
  OR2_X1 U558 ( .A1(n749), .A2(G902), .ZN(n453) );
  AND2_X1 U559 ( .A1(n454), .A2(n453), .ZN(n455) );
  AND2_X1 U560 ( .A1(n692), .A2(n455), .ZN(n570) );
  NAND2_X1 U561 ( .A1(n754), .A2(G900), .ZN(n456) );
  NAND2_X1 U562 ( .A1(n570), .A2(n456), .ZN(n457) );
  XOR2_X1 U563 ( .A(KEYINPUT78), .B(n457), .Z(n527) );
  XNOR2_X1 U564 ( .A(n482), .B(n470), .ZN(n745) );
  NAND2_X1 U565 ( .A1(n749), .A2(G234), .ZN(n458) );
  XNOR2_X2 U566 ( .A(n465), .B(n359), .ZN(n697) );
  INV_X1 U567 ( .A(n697), .ZN(n608) );
  AND2_X1 U568 ( .A1(n527), .A2(n608), .ZN(n466) );
  NAND2_X1 U569 ( .A1(n698), .A2(n466), .ZN(n534) );
  NOR2_X1 U570 ( .A1(n467), .A2(n534), .ZN(n468) );
  XOR2_X1 U571 ( .A(KEYINPUT28), .B(n468), .Z(n475) );
  NAND2_X1 U572 ( .A1(G227), .A2(n749), .ZN(n472) );
  XOR2_X1 U573 ( .A(n472), .B(n471), .Z(n473) );
  NOR2_X1 U574 ( .A1(n475), .A2(n532), .ZN(n543) );
  INV_X1 U575 ( .A(n543), .ZN(n524) );
  XNOR2_X1 U576 ( .A(n476), .B(G104), .ZN(n504) );
  XNOR2_X1 U577 ( .A(n504), .B(KEYINPUT93), .ZN(n480) );
  XNOR2_X1 U578 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U579 ( .A(n480), .B(n479), .ZN(n481) );
  XOR2_X1 U580 ( .A(n482), .B(n481), .Z(n488) );
  XOR2_X1 U581 ( .A(G140), .B(KEYINPUT92), .Z(n484) );
  XNOR2_X1 U582 ( .A(n484), .B(n483), .ZN(n486) );
  NOR2_X1 U583 ( .A1(G902), .A2(n651), .ZN(n491) );
  XNOR2_X1 U584 ( .A(KEYINPUT13), .B(KEYINPUT94), .ZN(n489) );
  NAND2_X1 U585 ( .A1(G217), .A2(n492), .ZN(n493) );
  XNOR2_X1 U586 ( .A(n494), .B(n493), .ZN(n497) );
  XNOR2_X1 U587 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n495) );
  XNOR2_X2 U588 ( .A(G116), .B(G107), .ZN(n503) );
  XNOR2_X1 U589 ( .A(n495), .B(n503), .ZN(n496) );
  XNOR2_X1 U590 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U591 ( .A(n499), .B(n498), .ZN(n736) );
  NOR2_X1 U592 ( .A1(G902), .A2(n736), .ZN(n501) );
  XOR2_X1 U593 ( .A(KEYINPUT96), .B(G478), .Z(n500) );
  XNOR2_X1 U594 ( .A(n501), .B(n500), .ZN(n575) );
  OR2_X1 U595 ( .A1(n576), .A2(n575), .ZN(n713) );
  XOR2_X1 U596 ( .A(KEYINPUT74), .B(KEYINPUT38), .Z(n521) );
  XNOR2_X1 U597 ( .A(G110), .B(KEYINPUT16), .ZN(n502) );
  XNOR2_X1 U598 ( .A(n503), .B(n502), .ZN(n505) );
  XNOR2_X1 U599 ( .A(n505), .B(n504), .ZN(n507) );
  XNOR2_X1 U600 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n509) );
  NAND2_X1 U601 ( .A1(n749), .A2(G224), .ZN(n508) );
  XNOR2_X1 U602 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U603 ( .A(n511), .B(n510), .ZN(n515) );
  XNOR2_X1 U604 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U605 ( .A(n515), .B(n514), .ZN(n516) );
  INV_X1 U606 ( .A(n517), .ZN(n617) );
  NAND2_X1 U607 ( .A1(n519), .A2(n518), .ZN(n522) );
  NAND2_X1 U608 ( .A1(n522), .A2(G210), .ZN(n520) );
  NAND2_X1 U609 ( .A1(n522), .A2(G214), .ZN(n710) );
  NOR2_X1 U610 ( .A1(n713), .A2(n715), .ZN(n523) );
  XNOR2_X1 U611 ( .A(KEYINPUT41), .B(n523), .ZN(n727) );
  NOR2_X1 U612 ( .A1(n524), .A2(n727), .ZN(n525) );
  XNOR2_X1 U613 ( .A(n525), .B(KEYINPUT42), .ZN(n764) );
  INV_X1 U614 ( .A(KEYINPUT30), .ZN(n528) );
  INV_X1 U615 ( .A(n575), .ZN(n550) );
  AND2_X1 U616 ( .A1(n576), .A2(n550), .ZN(n544) );
  XNOR2_X1 U617 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n531) );
  XNOR2_X1 U618 ( .A(KEYINPUT100), .B(n544), .ZN(n680) );
  INV_X1 U619 ( .A(n680), .ZN(n537) );
  XNOR2_X1 U620 ( .A(KEYINPUT6), .B(KEYINPUT97), .ZN(n533) );
  XNOR2_X1 U621 ( .A(n535), .B(KEYINPUT101), .ZN(n536) );
  NAND2_X1 U622 ( .A1(n538), .A2(n710), .ZN(n559) );
  INV_X1 U623 ( .A(KEYINPUT69), .ZN(n540) );
  XNOR2_X1 U624 ( .A(n540), .B(KEYINPUT19), .ZN(n541) );
  NAND2_X1 U625 ( .A1(n543), .A2(n572), .ZN(n548) );
  INV_X1 U626 ( .A(n544), .ZN(n545) );
  OR2_X1 U627 ( .A1(n576), .A2(n550), .ZN(n564) );
  AND2_X1 U628 ( .A1(n545), .A2(n564), .ZN(n716) );
  NOR2_X1 U629 ( .A1(n716), .A2(KEYINPUT47), .ZN(n546) );
  XNOR2_X1 U630 ( .A(n546), .B(KEYINPUT73), .ZN(n547) );
  INV_X1 U631 ( .A(n716), .ZN(n606) );
  NAND2_X1 U632 ( .A1(n677), .A2(n606), .ZN(n549) );
  NAND2_X1 U633 ( .A1(n549), .A2(KEYINPUT47), .ZN(n557) );
  NOR2_X1 U634 ( .A1(n550), .A2(n562), .ZN(n551) );
  AND2_X1 U635 ( .A1(n576), .A2(n551), .ZN(n552) );
  XNOR2_X2 U636 ( .A(n555), .B(n554), .ZN(n763) );
  NAND2_X1 U637 ( .A1(n557), .A2(n556), .ZN(n558) );
  NOR2_X1 U638 ( .A1(n414), .A2(n559), .ZN(n560) );
  XNOR2_X1 U639 ( .A(n560), .B(KEYINPUT43), .ZN(n561) );
  XOR2_X1 U640 ( .A(n561), .B(KEYINPUT102), .Z(n563) );
  NAND2_X1 U641 ( .A1(n563), .A2(n562), .ZN(n640) );
  INV_X1 U642 ( .A(n564), .ZN(n682) );
  NAND2_X1 U643 ( .A1(n565), .A2(n682), .ZN(n689) );
  AND2_X1 U644 ( .A1(n640), .A2(n689), .ZN(n566) );
  INV_X1 U645 ( .A(KEYINPUT82), .ZN(n567) );
  NOR2_X1 U646 ( .A1(n693), .A2(n694), .ZN(n568) );
  XNOR2_X1 U647 ( .A(n568), .B(KEYINPUT75), .ZN(n599) );
  NAND2_X1 U648 ( .A1(n754), .A2(G898), .ZN(n569) );
  AND2_X1 U649 ( .A1(n570), .A2(n569), .ZN(n571) );
  NAND2_X1 U650 ( .A1(n572), .A2(n571), .ZN(n574) );
  XNOR2_X1 U651 ( .A(KEYINPUT84), .B(KEYINPUT0), .ZN(n573) );
  XNOR2_X1 U652 ( .A(n574), .B(n573), .ZN(n584) );
  INV_X1 U653 ( .A(KEYINPUT70), .ZN(n578) );
  NOR2_X1 U654 ( .A1(n578), .A2(KEYINPUT44), .ZN(n577) );
  NAND2_X1 U655 ( .A1(n597), .A2(n577), .ZN(n580) );
  NAND2_X1 U656 ( .A1(n757), .A2(n578), .ZN(n579) );
  NAND2_X1 U657 ( .A1(n580), .A2(n579), .ZN(n595) );
  XNOR2_X1 U658 ( .A(KEYINPUT77), .B(n581), .ZN(n582) );
  NOR2_X1 U659 ( .A1(n582), .A2(n697), .ZN(n583) );
  NAND2_X1 U660 ( .A1(n583), .A2(n414), .ZN(n588) );
  INV_X1 U661 ( .A(n698), .ZN(n585) );
  NOR2_X1 U662 ( .A1(n713), .A2(n585), .ZN(n586) );
  NAND2_X1 U663 ( .A1(n604), .A2(n586), .ZN(n587) );
  XNOR2_X1 U664 ( .A(n587), .B(KEYINPUT22), .ZN(n590) );
  NOR2_X1 U665 ( .A1(n588), .A2(n590), .ZN(n589) );
  XNOR2_X1 U666 ( .A(n589), .B(KEYINPUT32), .ZN(n760) );
  XNOR2_X1 U667 ( .A(n592), .B(KEYINPUT67), .ZN(n593) );
  NOR2_X1 U668 ( .A1(n760), .A2(n639), .ZN(n594) );
  NAND2_X1 U669 ( .A1(n595), .A2(n594), .ZN(n615) );
  INV_X1 U670 ( .A(n760), .ZN(n596) );
  NOR2_X1 U671 ( .A1(n702), .A2(n599), .ZN(n600) );
  XNOR2_X1 U672 ( .A(KEYINPUT90), .B(n600), .ZN(n707) );
  AND2_X1 U673 ( .A1(n707), .A2(n604), .ZN(n602) );
  INV_X1 U674 ( .A(KEYINPUT31), .ZN(n601) );
  XNOR2_X1 U675 ( .A(n602), .B(n601), .ZN(n683) );
  AND2_X1 U676 ( .A1(n603), .A2(n702), .ZN(n605) );
  AND2_X1 U677 ( .A1(n605), .A2(n604), .ZN(n671) );
  OR2_X1 U678 ( .A1(n683), .A2(n671), .ZN(n607) );
  NAND2_X1 U679 ( .A1(n607), .A2(n606), .ZN(n613) );
  NOR2_X1 U680 ( .A1(n609), .A2(n608), .ZN(n610) );
  NAND2_X1 U681 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U682 ( .A(n612), .B(KEYINPUT98), .ZN(n758) );
  AND2_X1 U683 ( .A1(n613), .A2(n758), .ZN(n614) );
  XNOR2_X1 U684 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n616) );
  NAND2_X1 U685 ( .A1(n617), .A2(KEYINPUT2), .ZN(n618) );
  XOR2_X1 U686 ( .A(n618), .B(KEYINPUT68), .Z(n619) );
  INV_X1 U687 ( .A(n621), .ZN(n622) );
  NAND2_X1 U688 ( .A1(n622), .A2(KEYINPUT2), .ZN(n623) );
  OR2_X1 U689 ( .A1(n620), .A2(n623), .ZN(n691) );
  AND2_X2 U690 ( .A1(n624), .A2(n691), .ZN(n735) );
  NAND2_X1 U691 ( .A1(n735), .A2(G210), .ZN(n629) );
  XOR2_X1 U692 ( .A(KEYINPUT121), .B(KEYINPUT54), .Z(n625) );
  XOR2_X1 U693 ( .A(n625), .B(KEYINPUT55), .Z(n626) );
  XNOR2_X1 U694 ( .A(n627), .B(n626), .ZN(n628) );
  XNOR2_X1 U695 ( .A(n629), .B(n628), .ZN(n631) );
  NOR2_X2 U696 ( .A1(n631), .A2(n744), .ZN(n632) );
  XNOR2_X1 U697 ( .A(n632), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U698 ( .A1(n735), .A2(G472), .ZN(n635) );
  XOR2_X1 U699 ( .A(KEYINPUT62), .B(n633), .Z(n634) );
  XNOR2_X1 U700 ( .A(n635), .B(n634), .ZN(n636) );
  NOR2_X2 U701 ( .A1(n636), .A2(n744), .ZN(n638) );
  XNOR2_X1 U702 ( .A(KEYINPUT63), .B(KEYINPUT83), .ZN(n637) );
  XNOR2_X1 U703 ( .A(n638), .B(n637), .ZN(G57) );
  XOR2_X1 U704 ( .A(n639), .B(G110), .Z(G12) );
  XNOR2_X1 U705 ( .A(n640), .B(G140), .ZN(G42) );
  INV_X1 U706 ( .A(n620), .ZN(n641) );
  NAND2_X1 U707 ( .A1(n641), .A2(n749), .ZN(n645) );
  NAND2_X1 U708 ( .A1(n754), .A2(G224), .ZN(n642) );
  XNOR2_X1 U709 ( .A(KEYINPUT61), .B(n642), .ZN(n643) );
  NAND2_X1 U710 ( .A1(n643), .A2(G898), .ZN(n644) );
  NAND2_X1 U711 ( .A1(n645), .A2(n644), .ZN(n650) );
  INV_X1 U712 ( .A(n646), .ZN(n648) );
  NOR2_X1 U713 ( .A1(G898), .A2(n749), .ZN(n647) );
  NOR2_X1 U714 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U715 ( .A(n650), .B(n649), .ZN(G69) );
  NAND2_X1 U716 ( .A1(n735), .A2(G475), .ZN(n653) );
  XNOR2_X1 U717 ( .A(n651), .B(KEYINPUT59), .ZN(n652) );
  XNOR2_X1 U718 ( .A(n653), .B(n652), .ZN(n654) );
  INV_X1 U719 ( .A(n744), .ZN(n663) );
  NAND2_X1 U720 ( .A1(n654), .A2(n663), .ZN(n656) );
  XNOR2_X1 U721 ( .A(KEYINPUT125), .B(KEYINPUT60), .ZN(n655) );
  XNOR2_X1 U722 ( .A(n656), .B(n655), .ZN(G60) );
  NAND2_X1 U723 ( .A1(n735), .A2(G469), .ZN(n662) );
  XNOR2_X1 U724 ( .A(KEYINPUT123), .B(KEYINPUT57), .ZN(n659) );
  XNOR2_X1 U725 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n658) );
  XNOR2_X1 U726 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U727 ( .A(n657), .B(n660), .ZN(n661) );
  XNOR2_X1 U728 ( .A(n662), .B(n661), .ZN(n664) );
  NAND2_X1 U729 ( .A1(n664), .A2(n663), .ZN(n666) );
  INV_X1 U730 ( .A(KEYINPUT124), .ZN(n665) );
  XNOR2_X1 U731 ( .A(n666), .B(n665), .ZN(G54) );
  NAND2_X1 U732 ( .A1(n680), .A2(n671), .ZN(n667) );
  XNOR2_X1 U733 ( .A(n667), .B(G104), .ZN(G6) );
  XOR2_X1 U734 ( .A(KEYINPUT27), .B(KEYINPUT107), .Z(n669) );
  XNOR2_X1 U735 ( .A(G107), .B(KEYINPUT106), .ZN(n668) );
  XNOR2_X1 U736 ( .A(n669), .B(n668), .ZN(n670) );
  XOR2_X1 U737 ( .A(KEYINPUT26), .B(n670), .Z(n673) );
  NAND2_X1 U738 ( .A1(n671), .A2(n682), .ZN(n672) );
  XNOR2_X1 U739 ( .A(n673), .B(n672), .ZN(G9) );
  XOR2_X1 U740 ( .A(KEYINPUT108), .B(KEYINPUT29), .Z(n675) );
  NAND2_X1 U741 ( .A1(n677), .A2(n682), .ZN(n674) );
  XNOR2_X1 U742 ( .A(n675), .B(n674), .ZN(n676) );
  XNOR2_X1 U743 ( .A(G128), .B(n676), .ZN(G30) );
  XOR2_X1 U744 ( .A(G146), .B(KEYINPUT109), .Z(n679) );
  NAND2_X1 U745 ( .A1(n677), .A2(n680), .ZN(n678) );
  XNOR2_X1 U746 ( .A(n679), .B(n678), .ZN(G48) );
  NAND2_X1 U747 ( .A1(n680), .A2(n683), .ZN(n681) );
  XNOR2_X1 U748 ( .A(n681), .B(G113), .ZN(G15) );
  NAND2_X1 U749 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U750 ( .A(n684), .B(KEYINPUT110), .ZN(n685) );
  XNOR2_X1 U751 ( .A(G116), .B(n685), .ZN(G18) );
  XOR2_X1 U752 ( .A(KEYINPUT111), .B(KEYINPUT37), .Z(n688) );
  XNOR2_X1 U753 ( .A(n686), .B(G125), .ZN(n687) );
  XNOR2_X1 U754 ( .A(n688), .B(n687), .ZN(G27) );
  XNOR2_X1 U755 ( .A(G134), .B(n689), .ZN(G36) );
  INV_X1 U756 ( .A(n748), .ZN(n690) );
  NAND2_X1 U757 ( .A1(G952), .A2(n692), .ZN(n726) );
  XOR2_X1 U758 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n696) );
  NAND2_X1 U759 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U760 ( .A(n696), .B(n695), .ZN(n705) );
  OR2_X1 U761 ( .A1(n698), .A2(n697), .ZN(n701) );
  XNOR2_X1 U762 ( .A(KEYINPUT112), .B(KEYINPUT49), .ZN(n699) );
  XNOR2_X1 U763 ( .A(n699), .B(KEYINPUT113), .ZN(n700) );
  XNOR2_X1 U764 ( .A(n701), .B(n700), .ZN(n703) );
  NAND2_X1 U765 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U766 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U767 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U768 ( .A(KEYINPUT51), .B(n708), .Z(n709) );
  NOR2_X1 U769 ( .A1(n727), .A2(n709), .ZN(n722) );
  NOR2_X1 U770 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U771 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U772 ( .A(KEYINPUT115), .B(n714), .Z(n719) );
  NOR2_X1 U773 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U774 ( .A(KEYINPUT116), .B(n717), .ZN(n718) );
  XOR2_X1 U775 ( .A(KEYINPUT117), .B(n720), .Z(n721) );
  NOR2_X1 U776 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U777 ( .A(KEYINPUT52), .B(n723), .Z(n724) );
  XOR2_X1 U778 ( .A(KEYINPUT118), .B(n724), .Z(n725) );
  NOR2_X1 U779 ( .A1(n726), .A2(n725), .ZN(n730) );
  XOR2_X1 U780 ( .A(KEYINPUT119), .B(n728), .Z(n729) );
  NOR2_X1 U781 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U782 ( .A(KEYINPUT120), .B(n731), .ZN(n732) );
  NOR2_X1 U783 ( .A1(n733), .A2(n754), .ZN(n734) );
  XNOR2_X1 U784 ( .A(n734), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U785 ( .A1(n740), .A2(G478), .ZN(n738) );
  XNOR2_X1 U786 ( .A(n736), .B(KEYINPUT126), .ZN(n737) );
  XNOR2_X1 U787 ( .A(n738), .B(n737), .ZN(n739) );
  NOR2_X1 U788 ( .A1(n744), .A2(n739), .ZN(G63) );
  NAND2_X1 U789 ( .A1(n740), .A2(G217), .ZN(n742) );
  XNOR2_X1 U790 ( .A(n741), .B(n742), .ZN(n743) );
  NOR2_X1 U791 ( .A1(n744), .A2(n743), .ZN(G66) );
  XOR2_X1 U792 ( .A(n745), .B(KEYINPUT86), .Z(n746) );
  XOR2_X1 U793 ( .A(n747), .B(n746), .Z(n751) );
  XOR2_X1 U794 ( .A(n748), .B(n751), .Z(n750) );
  NAND2_X1 U795 ( .A1(n750), .A2(n749), .ZN(n756) );
  XNOR2_X1 U796 ( .A(G227), .B(n751), .ZN(n752) );
  NAND2_X1 U797 ( .A1(n752), .A2(G900), .ZN(n753) );
  NAND2_X1 U798 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U799 ( .A1(n756), .A2(n755), .ZN(G72) );
  XOR2_X1 U800 ( .A(G122), .B(n757), .Z(G24) );
  XOR2_X1 U801 ( .A(G101), .B(n758), .Z(n759) );
  XNOR2_X1 U802 ( .A(KEYINPUT105), .B(n759), .ZN(G3) );
  XNOR2_X1 U803 ( .A(G119), .B(KEYINPUT127), .ZN(n761) );
  XNOR2_X1 U804 ( .A(n761), .B(n760), .ZN(G21) );
  XOR2_X1 U805 ( .A(n762), .B(G131), .Z(G33) );
  XNOR2_X1 U806 ( .A(n357), .B(n763), .ZN(G45) );
  XOR2_X1 U807 ( .A(n764), .B(G137), .Z(G39) );
endmodule

