//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 0 1 1 0 0 0 0 1 0 1 0 0 1 0 0 1 1 1 0 1 1 0 0 1 1 0 1 0 0 1 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:55 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n561, new_n562, new_n563, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n575, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n612, new_n615, new_n617, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1208,
    new_n1209;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT66), .ZN(G234));
  NAND2_X1  g026(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT67), .Z(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n454), .ZN(new_n461));
  AOI21_X1  g036(.A(new_n460), .B1(new_n461), .B2(G2106), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n462), .B(KEYINPUT68), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  OAI211_X1 g041(.A(G137), .B(new_n464), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g046(.A(G125), .B1(new_n465), .B2(new_n466), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g049(.A(KEYINPUT3), .B(G2104), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(KEYINPUT69), .A3(G125), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n474), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n471), .B1(new_n478), .B2(G2105), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT70), .ZN(G160));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n482));
  XOR2_X1   g057(.A(new_n482), .B(KEYINPUT73), .Z(new_n483));
  XNOR2_X1  g058(.A(new_n475), .B(KEYINPUT71), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(new_n464), .ZN(new_n485));
  INV_X1    g060(.A(G136), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n483), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n484), .A2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(G124), .ZN(new_n489));
  OR3_X1    g064(.A1(new_n488), .A2(KEYINPUT72), .A3(new_n489), .ZN(new_n490));
  OAI21_X1  g065(.A(KEYINPUT72), .B1(new_n488), .B2(new_n489), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n487), .B1(new_n490), .B2(new_n491), .ZN(G162));
  AND2_X1   g067(.A1(G126), .A2(G2105), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(G114), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  AOI22_X1  g072(.A1(new_n475), .A2(new_n493), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G138), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n499), .A2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  OAI211_X1 g076(.A(new_n500), .B(new_n501), .C1(new_n466), .C2(new_n465), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n501), .B1(new_n475), .B2(new_n500), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n498), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT74), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI211_X1 g082(.A(KEYINPUT74), .B(new_n498), .C1(new_n503), .C2(new_n504), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(G164));
  OR2_X1    g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  OR2_X1    g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G50), .ZN(new_n521));
  INV_X1    g096(.A(G88), .ZN(new_n522));
  NOR2_X1   g097(.A1(KEYINPUT5), .A2(G543), .ZN(new_n523));
  AND2_X1   g098(.A1(KEYINPUT5), .A2(G543), .ZN(new_n524));
  AND2_X1   g099(.A1(KEYINPUT6), .A2(G651), .ZN(new_n525));
  NOR2_X1   g100(.A1(KEYINPUT6), .A2(G651), .ZN(new_n526));
  OAI22_X1  g101(.A1(new_n523), .A2(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n521), .B1(new_n522), .B2(new_n527), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n516), .A2(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT75), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT7), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n532), .B(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n520), .A2(G51), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n518), .A2(new_n519), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n536), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n524), .A2(new_n523), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n535), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n534), .A2(new_n539), .ZN(G168));
  NAND2_X1  g115(.A1(G77), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G64), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n538), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G651), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT76), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n543), .A2(KEYINPUT76), .A3(G651), .ZN(new_n547));
  INV_X1    g122(.A(new_n527), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n548), .A2(G90), .B1(G52), .B2(new_n520), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n546), .A2(new_n547), .A3(new_n549), .ZN(G301));
  INV_X1    g125(.A(G301), .ZN(G171));
  AOI22_X1  g126(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n552), .A2(new_n515), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n520), .A2(G43), .ZN(new_n554));
  INV_X1    g129(.A(G81), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n555), .B2(new_n527), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(new_n558));
  XOR2_X1   g133(.A(new_n558), .B(KEYINPUT77), .Z(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g135(.A(KEYINPUT78), .B(KEYINPUT8), .Z(new_n561));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n561), .B(new_n562), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(G188));
  NAND2_X1  g139(.A1(new_n520), .A2(G53), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT9), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n527), .A2(KEYINPUT79), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT79), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n513), .A2(new_n536), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n567), .A2(G91), .A3(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n513), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n571));
  OR2_X1    g146(.A1(new_n571), .A2(new_n515), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n566), .A2(new_n570), .A3(new_n572), .ZN(G299));
  INV_X1    g148(.A(G168), .ZN(G286));
  NAND3_X1  g149(.A1(new_n567), .A2(G87), .A3(new_n569), .ZN(new_n575));
  INV_X1    g150(.A(G74), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n511), .A2(new_n576), .A3(new_n512), .ZN(new_n577));
  AOI22_X1  g152(.A1(G49), .A2(new_n520), .B1(new_n577), .B2(G651), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n575), .A2(new_n578), .ZN(G288));
  OAI211_X1 g154(.A(G48), .B(G543), .C1(new_n525), .C2(new_n526), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(KEYINPUT80), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT80), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n536), .A2(new_n582), .A3(G48), .A4(G543), .ZN(new_n583));
  OAI21_X1  g158(.A(G61), .B1(new_n524), .B2(new_n523), .ZN(new_n584));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n581), .A2(new_n583), .B1(new_n586), .B2(G651), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n567), .A2(G86), .A3(new_n569), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(G305));
  AOI22_X1  g164(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n590), .A2(new_n515), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n520), .A2(G47), .ZN(new_n592));
  INV_X1    g167(.A(G85), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n593), .B2(new_n527), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT81), .ZN(new_n595));
  OR3_X1    g170(.A1(new_n591), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n591), .B2(new_n594), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(G290));
  NAND2_X1  g173(.A1(G301), .A2(G868), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n567), .A2(G92), .A3(new_n569), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT10), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n600), .B(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(G79), .A2(G543), .ZN(new_n603));
  INV_X1    g178(.A(G66), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n538), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n605), .A2(G651), .B1(G54), .B2(new_n520), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n599), .B1(new_n608), .B2(G868), .ZN(G284));
  OAI21_X1  g184(.A(new_n599), .B1(new_n608), .B2(G868), .ZN(G321));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(G299), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(new_n611), .B2(G168), .ZN(G297));
  OAI21_X1  g188(.A(new_n612), .B1(new_n611), .B2(G168), .ZN(G280));
  XOR2_X1   g189(.A(KEYINPUT82), .B(G559), .Z(new_n615));
  OAI21_X1  g190(.A(new_n608), .B1(G860), .B2(new_n615), .ZN(G148));
  INV_X1    g191(.A(new_n557), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(new_n611), .ZN(new_n618));
  AND2_X1   g193(.A1(new_n608), .A2(new_n615), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(new_n611), .ZN(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g196(.A(new_n485), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G135), .ZN(new_n623));
  INV_X1    g198(.A(new_n488), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(G123), .ZN(new_n625));
  OR2_X1    g200(.A1(G99), .A2(G2105), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n626), .B(G2104), .C1(G111), .C2(new_n464), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n623), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT83), .B(G2096), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n475), .A2(new_n469), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT12), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT13), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2100), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n631), .A2(new_n632), .A3(new_n636), .ZN(G156));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2435), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT85), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2427), .B(G2430), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(KEYINPUT14), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2451), .B(G2454), .Z(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n646), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT86), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT87), .ZN(new_n654));
  INV_X1    g229(.A(G14), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n655), .B1(new_n650), .B2(new_n652), .ZN(new_n656));
  AND2_X1   g231(.A1(new_n654), .A2(new_n656), .ZN(G401));
  XNOR2_X1  g232(.A(G2067), .B(G2678), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT88), .ZN(new_n659));
  NOR2_X1   g234(.A1(G2072), .A2(G2078), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n442), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2084), .B(G2090), .ZN(new_n662));
  NOR3_X1   g237(.A1(new_n659), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT18), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n659), .A2(new_n661), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n661), .B(KEYINPUT17), .ZN(new_n666));
  OAI211_X1 g241(.A(new_n665), .B(new_n662), .C1(new_n659), .C2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n662), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n666), .A2(new_n659), .A3(new_n668), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n664), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(G2100), .Z(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT89), .B(G2096), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(G227));
  XNOR2_X1  g249(.A(G1956), .B(G2474), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1961), .B(G1966), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1971), .B(G1976), .ZN(new_n678));
  INV_X1    g253(.A(KEYINPUT19), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n675), .A2(new_n676), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n677), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n680), .A2(KEYINPUT90), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n683), .B(new_n684), .Z(new_n685));
  NAND2_X1  g260(.A1(new_n680), .A2(new_n681), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n686), .B(KEYINPUT20), .Z(new_n687));
  OR3_X1    g262(.A1(new_n685), .A2(G1981), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g263(.A(G1981), .B1(new_n685), .B2(new_n687), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(G1986), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT91), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n690), .A2(new_n691), .ZN(new_n697));
  AND3_X1   g272(.A1(new_n693), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n696), .B1(new_n693), .B2(new_n697), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1991), .B(G1996), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n701), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(new_n698), .B2(new_n699), .ZN(new_n704));
  AND2_X1   g279(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(G229));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G24), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n596), .A2(new_n597), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n708), .B1(new_n709), .B2(new_n707), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(G1986), .ZN(new_n711));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G25), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n622), .A2(G131), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n624), .A2(G119), .ZN(new_n715));
  OR2_X1    g290(.A1(G95), .A2(G2105), .ZN(new_n716));
  OAI211_X1 g291(.A(new_n716), .B(G2104), .C1(G107), .C2(new_n464), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n714), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n713), .B1(new_n719), .B2(new_n712), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT92), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT35), .B(G1991), .Z(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT93), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT92), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n720), .B(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(new_n723), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n711), .B1(new_n725), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n707), .A2(G6), .ZN(new_n730));
  INV_X1    g305(.A(G305), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(new_n731), .B2(new_n707), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT32), .B(G1981), .Z(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT94), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n707), .A2(G22), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G166), .B2(new_n707), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT95), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n735), .B1(new_n739), .B2(G1971), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n707), .A2(G23), .ZN(new_n741));
  INV_X1    g316(.A(G288), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n741), .B1(new_n742), .B2(new_n707), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT33), .B(G1976), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(G1971), .ZN(new_n746));
  AOI22_X1  g321(.A1(new_n738), .A2(new_n746), .B1(new_n734), .B2(new_n732), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n740), .A2(new_n745), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(KEYINPUT34), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT34), .ZN(new_n750));
  NAND4_X1  g325(.A1(new_n740), .A2(new_n750), .A3(new_n745), .A4(new_n747), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n729), .A2(new_n749), .A3(new_n751), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT96), .B(KEYINPUT36), .Z(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n622), .A2(G139), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT101), .Z(new_n756));
  NAND2_X1  g331(.A1(new_n475), .A2(G127), .ZN(new_n757));
  INV_X1    g332(.A(G115), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n757), .B1(new_n758), .B2(new_n468), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT25), .ZN(new_n760));
  NAND2_X1  g335(.A1(G103), .A2(G2104), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n760), .B1(new_n761), .B2(G2105), .ZN(new_n762));
  NAND4_X1  g337(.A1(new_n464), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n763));
  AOI22_X1  g338(.A1(new_n759), .A2(G2105), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n756), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n765), .A2(G29), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n712), .A2(G33), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G2072), .ZN(new_n769));
  NOR2_X1   g344(.A1(G29), .A2(G35), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G162), .B2(G29), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT29), .B(G2090), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n622), .A2(G141), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n624), .A2(G129), .ZN(new_n775));
  NAND3_X1  g350(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT26), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n776), .A2(new_n777), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n778), .A2(new_n779), .B1(G105), .B2(new_n469), .ZN(new_n780));
  AND3_X1   g355(.A1(new_n774), .A2(new_n775), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n781), .A2(G29), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT103), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G29), .B2(G32), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(KEYINPUT103), .B2(new_n782), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT27), .B(G1996), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n707), .A2(G20), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT23), .ZN(new_n790));
  INV_X1    g365(.A(G299), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n790), .B1(new_n791), .B2(new_n707), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(G1956), .Z(new_n793));
  NAND2_X1  g368(.A1(new_n707), .A2(G5), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G171), .B2(new_n707), .ZN(new_n795));
  INV_X1    g370(.A(G1961), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n793), .A2(new_n797), .ZN(new_n798));
  NOR4_X1   g373(.A1(new_n769), .A2(new_n773), .A3(new_n788), .A4(new_n798), .ZN(new_n799));
  OAI21_X1  g374(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n800));
  INV_X1    g375(.A(G116), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n800), .B1(new_n801), .B2(G2105), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n622), .B2(G140), .ZN(new_n803));
  AND3_X1   g378(.A1(new_n624), .A2(KEYINPUT98), .A3(G128), .ZN(new_n804));
  AOI21_X1  g379(.A(KEYINPUT98), .B1(new_n624), .B2(G128), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(G29), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT99), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n712), .A2(G26), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT28), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(G2067), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(G16), .A2(G19), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(new_n557), .B2(G16), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT97), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(G1341), .Z(new_n817));
  NOR2_X1   g392(.A1(G4), .A2(G16), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(new_n608), .B2(G16), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(G1348), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n819), .A2(G1348), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n817), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n813), .A2(KEYINPUT100), .A3(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(G27), .A2(G29), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(G164), .B2(G29), .ZN(new_n826));
  INV_X1    g401(.A(G2078), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT30), .B(G28), .ZN(new_n829));
  OR2_X1    g404(.A1(KEYINPUT31), .A2(G11), .ZN(new_n830));
  NAND2_X1  g405(.A1(KEYINPUT31), .A2(G11), .ZN(new_n831));
  AOI22_X1  g406(.A1(new_n829), .A2(new_n712), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(new_n628), .B2(new_n712), .ZN(new_n833));
  INV_X1    g408(.A(G1966), .ZN(new_n834));
  NOR2_X1   g409(.A1(G168), .A2(new_n707), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(new_n707), .B2(G21), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n833), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n828), .B(new_n837), .C1(new_n834), .C2(new_n836), .ZN(new_n838));
  NAND2_X1  g413(.A1(G160), .A2(G29), .ZN(new_n839));
  XOR2_X1   g414(.A(KEYINPUT102), .B(KEYINPUT24), .Z(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(G34), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n839), .B1(G29), .B2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(G2084), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n842), .A2(new_n843), .ZN(new_n845));
  NOR3_X1   g420(.A1(new_n838), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  AND3_X1   g421(.A1(new_n799), .A2(new_n824), .A3(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT100), .ZN(new_n848));
  INV_X1    g423(.A(new_n813), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n848), .B1(new_n849), .B2(new_n822), .ZN(new_n850));
  AND3_X1   g425(.A1(new_n754), .A2(new_n847), .A3(new_n850), .ZN(G311));
  NAND3_X1  g426(.A1(new_n754), .A2(new_n847), .A3(new_n850), .ZN(G150));
  AOI22_X1  g427(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n853), .A2(new_n515), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n520), .A2(G55), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n513), .A2(new_n536), .A3(G93), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT104), .ZN(new_n857));
  AND3_X1   g432(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n857), .B1(new_n855), .B2(new_n856), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n854), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT105), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n557), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n862), .B1(new_n861), .B2(new_n860), .ZN(new_n863));
  INV_X1    g438(.A(new_n860), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n864), .A2(KEYINPUT105), .A3(new_n557), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT38), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n608), .A2(G559), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT39), .ZN(new_n870));
  AOI21_X1  g445(.A(G860), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n871), .B1(new_n870), .B2(new_n869), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n860), .A2(G860), .ZN(new_n873));
  XOR2_X1   g448(.A(KEYINPUT106), .B(KEYINPUT37), .Z(new_n874));
  XNOR2_X1  g449(.A(new_n873), .B(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n872), .A2(new_n875), .ZN(G145));
  NAND2_X1  g451(.A1(new_n622), .A2(G142), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n624), .A2(G130), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n464), .A2(G118), .ZN(new_n879));
  OAI21_X1  g454(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n877), .B(new_n878), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(new_n634), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n756), .A2(new_n781), .A3(new_n764), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n781), .B1(new_n756), .B2(new_n764), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n885), .ZN(new_n887));
  INV_X1    g462(.A(new_n882), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n887), .A2(new_n888), .A3(new_n883), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n806), .B(new_n505), .ZN(new_n891));
  OR2_X1    g466(.A1(new_n891), .A2(new_n719), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n719), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n889), .A2(new_n886), .A3(new_n892), .A4(new_n893), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  XOR2_X1   g472(.A(G162), .B(G160), .Z(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(new_n629), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(G37), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n895), .A2(new_n899), .A3(new_n896), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g480(.A1(new_n709), .A2(G305), .ZN(new_n906));
  XNOR2_X1  g481(.A(G303), .B(new_n742), .ZN(new_n907));
  NOR2_X1   g482(.A1(G290), .A2(new_n731), .ZN(new_n908));
  OR3_X1    g483(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n907), .B1(new_n906), .B2(new_n908), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(KEYINPUT107), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n619), .B(new_n866), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n607), .A2(G299), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n607), .A2(G299), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n917), .A2(KEYINPUT41), .A3(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT41), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n791), .B1(new_n602), .B2(new_n606), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n920), .B1(new_n921), .B2(new_n916), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n919), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n915), .A2(new_n923), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n619), .A2(new_n865), .A3(new_n863), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n619), .B1(new_n865), .B2(new_n863), .ZN(new_n926));
  OAI22_X1  g501(.A1(new_n925), .A2(new_n926), .B1(new_n921), .B2(new_n916), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT42), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n924), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n928), .B1(new_n924), .B2(new_n927), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n914), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n924), .A2(new_n927), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(KEYINPUT42), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n924), .A2(new_n927), .A3(new_n928), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n933), .A2(new_n913), .A3(new_n934), .ZN(new_n935));
  AND4_X1   g510(.A1(KEYINPUT108), .A2(new_n931), .A3(new_n935), .A4(G868), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n931), .A2(new_n935), .A3(G868), .ZN(new_n937));
  AOI21_X1  g512(.A(KEYINPUT108), .B1(new_n860), .B2(new_n611), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(G295));
  AOI21_X1  g514(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(G331));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n941));
  XNOR2_X1  g516(.A(G168), .B(G301), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n863), .A2(new_n942), .A3(new_n865), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n942), .B1(new_n863), .B2(new_n865), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n922), .B(new_n919), .C1(new_n944), .C2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n942), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n866), .A2(new_n947), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n948), .A2(new_n918), .A3(new_n917), .A4(new_n943), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n946), .A2(new_n949), .A3(KEYINPUT109), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n948), .A2(new_n943), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT109), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n951), .A2(new_n952), .A3(new_n922), .A4(new_n919), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n950), .A2(new_n912), .A3(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n946), .A2(new_n911), .A3(new_n949), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n954), .A2(KEYINPUT43), .A3(new_n902), .A4(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n955), .A2(new_n902), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n911), .B1(new_n946), .B2(new_n949), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n957), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n941), .B1(new_n956), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n954), .A2(new_n957), .A3(new_n902), .A4(new_n955), .ZN(new_n963));
  OAI21_X1  g538(.A(KEYINPUT43), .B1(new_n958), .B2(new_n959), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(new_n941), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT110), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n962), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(KEYINPUT44), .B1(new_n963), .B2(new_n964), .ZN(new_n969));
  OAI21_X1  g544(.A(KEYINPUT110), .B1(new_n961), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n968), .A2(new_n970), .ZN(G397));
  XNOR2_X1  g546(.A(new_n806), .B(G2067), .ZN(new_n972));
  INV_X1    g547(.A(G1996), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n781), .A2(new_n973), .ZN(new_n974));
  OR2_X1    g549(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g550(.A(KEYINPUT111), .B(G1384), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n505), .A2(new_n976), .ZN(new_n977));
  OR2_X1    g552(.A1(new_n977), .A2(KEYINPUT112), .ZN(new_n978));
  INV_X1    g553(.A(G40), .ZN(new_n979));
  AOI211_X1 g554(.A(new_n979), .B(new_n471), .C1(new_n478), .C2(G2105), .ZN(new_n980));
  AOI21_X1  g555(.A(KEYINPUT45), .B1(new_n977), .B2(KEYINPUT112), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n978), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  XOR2_X1   g557(.A(new_n982), .B(KEYINPUT113), .Z(new_n983));
  NOR2_X1   g558(.A1(new_n982), .A2(G1996), .ZN(new_n984));
  AOI22_X1  g559(.A1(new_n975), .A2(new_n983), .B1(new_n781), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n983), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n718), .B(new_n722), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n985), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n709), .A2(new_n691), .ZN(new_n989));
  NAND2_X1  g564(.A1(G290), .A2(G1986), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n982), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n988), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT50), .ZN(new_n993));
  INV_X1    g568(.A(G1384), .ZN(new_n994));
  INV_X1    g569(.A(new_n508), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n500), .B1(new_n465), .B2(new_n466), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT4), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(new_n502), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT74), .B1(new_n998), .B2(new_n498), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n993), .B(new_n994), .C1(new_n995), .C2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT114), .ZN(new_n1001));
  OR2_X1    g576(.A1(G102), .A2(G2105), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1002), .A2(new_n497), .A3(G2104), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n493), .B1(new_n465), .B2(new_n466), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1005), .B1(new_n997), .B2(new_n502), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1001), .B1(new_n1006), .B2(G1384), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n505), .A2(KEYINPUT114), .A3(new_n994), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1007), .A2(KEYINPUT50), .A3(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1000), .A2(new_n1009), .A3(new_n980), .ZN(new_n1010));
  XOR2_X1   g585(.A(KEYINPUT121), .B(G1956), .Z(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n994), .B1(new_n995), .B2(new_n999), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT45), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n977), .A2(new_n1014), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n479), .A2(G40), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g593(.A(KEYINPUT56), .B(G2072), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1015), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1012), .A2(new_n1020), .ZN(new_n1021));
  XOR2_X1   g596(.A(G299), .B(KEYINPUT57), .Z(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G1348), .ZN(new_n1025));
  NOR3_X1   g600(.A1(new_n1006), .A2(new_n1001), .A3(G1384), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT114), .B1(new_n505), .B2(new_n994), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n980), .B1(new_n1028), .B2(KEYINPUT50), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n993), .B1(new_n509), .B2(new_n994), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1025), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1032), .A2(new_n812), .A3(new_n980), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT122), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1017), .B1(new_n1032), .B2(new_n993), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1013), .A2(KEYINPUT50), .ZN(new_n1037));
  AOI21_X1  g612(.A(G1348), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT122), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1033), .ZN(new_n1040));
  NOR3_X1   g615(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1035), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1022), .A2(new_n1012), .A3(new_n1020), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(new_n608), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1024), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT60), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1047), .B1(new_n608), .B2(KEYINPUT123), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1048), .B1(new_n1034), .B2(new_n1041), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n608), .A2(KEYINPUT123), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  OAI221_X1 g626(.A(new_n1048), .B1(KEYINPUT123), .B2(new_n608), .C1(new_n1034), .C2(new_n1041), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1035), .A2(new_n1047), .A3(new_n1042), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1044), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1022), .B1(new_n1020), .B2(new_n1012), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT61), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1015), .A2(new_n1018), .A3(new_n973), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n980), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1060));
  XOR2_X1   g635(.A(KEYINPUT58), .B(G1341), .Z(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n617), .B1(new_n1059), .B2(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g638(.A(new_n1063), .B(KEYINPUT59), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT61), .B1(new_n1024), .B2(new_n1044), .ZN(new_n1065));
  NOR3_X1   g640(.A1(new_n1058), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1046), .B1(new_n1054), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT50), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1068));
  NOR3_X1   g643(.A1(new_n1030), .A2(new_n1068), .A3(new_n1017), .ZN(new_n1069));
  OAI21_X1  g644(.A(KEYINPUT126), .B1(new_n1069), .B2(G1961), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1015), .A2(new_n1018), .A3(new_n827), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT53), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1072), .A2(G2078), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1074), .B1(new_n978), .B2(new_n981), .ZN(new_n1075));
  AOI22_X1  g650(.A1(new_n1071), .A2(new_n1072), .B1(new_n1075), .B2(new_n1018), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT126), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(new_n1078), .A3(new_n796), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1070), .A2(new_n1076), .A3(G301), .A4(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT127), .ZN(new_n1081));
  XNOR2_X1  g656(.A(new_n1080), .B(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT125), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1007), .A2(new_n1014), .A3(new_n1008), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1085), .B(new_n980), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1086), .A2(new_n1074), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(G1961), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1084), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1091));
  NOR3_X1   g666(.A1(new_n1087), .A2(new_n1089), .A3(KEYINPUT125), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1083), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(G171), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT54), .B1(new_n1082), .B2(new_n1094), .ZN(new_n1095));
  OAI211_X1 g670(.A(G301), .B(new_n1083), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT54), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1070), .A2(new_n1076), .A3(new_n1079), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1097), .B1(new_n1098), .B2(G171), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1096), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1086), .A2(new_n834), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1101), .B(G168), .C1(new_n1077), .C2(G2084), .ZN(new_n1102));
  OAI21_X1  g677(.A(G8), .B1(KEYINPUT124), .B2(KEYINPUT51), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(KEYINPUT124), .A2(KEYINPUT51), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1101), .B1(new_n1077), .B2(G2084), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1109), .A2(G8), .A3(G286), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1102), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1108), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(G8), .ZN(new_n1113));
  NAND2_X1  g688(.A1(G303), .A2(G8), .ZN(new_n1114));
  XNOR2_X1  g689(.A(new_n1114), .B(KEYINPUT55), .ZN(new_n1115));
  INV_X1    g690(.A(G2090), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1069), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(KEYINPUT45), .B1(new_n509), .B2(new_n994), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n980), .B1(new_n1014), .B2(new_n977), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n746), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  AOI211_X1 g695(.A(new_n1113), .B(new_n1115), .C1(new_n1117), .C2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT49), .ZN(new_n1122));
  XNOR2_X1  g697(.A(KEYINPUT117), .B(G1981), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n587), .A2(new_n588), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(G1981), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n548), .A2(G86), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1125), .B1(new_n587), .B2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1122), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT118), .ZN(new_n1129));
  OR3_X1    g704(.A1(new_n1124), .A2(new_n1127), .A3(new_n1122), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT118), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1131), .B(new_n1122), .C1(new_n1124), .C2(new_n1127), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1113), .B1(new_n1032), .B2(new_n980), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1129), .A2(new_n1130), .A3(new_n1132), .A4(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT116), .ZN(new_n1135));
  XNOR2_X1  g710(.A(KEYINPUT115), .B(G1976), .ZN(new_n1136));
  NAND2_X1  g711(.A1(G288), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT52), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1135), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1136), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1140), .B1(new_n575), .B2(new_n578), .ZN(new_n1141));
  NOR3_X1   g716(.A1(new_n1141), .A2(KEYINPUT116), .A3(KEYINPUT52), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1139), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n742), .A2(G1976), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1060), .A2(G8), .A3(new_n1144), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(KEYINPUT52), .B1(new_n1133), .B2(new_n1144), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1134), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT120), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1134), .B(KEYINPUT120), .C1(new_n1146), .C2(new_n1147), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1121), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1000), .A2(new_n1009), .A3(new_n1116), .A4(new_n980), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(G1971), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1155));
  OAI21_X1  g730(.A(G8), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT119), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1156), .A2(new_n1157), .A3(new_n1115), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1113), .B1(new_n1120), .B2(new_n1153), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1115), .ZN(new_n1160));
  OAI21_X1  g735(.A(KEYINPUT119), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1158), .A2(new_n1161), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1100), .A2(new_n1112), .A3(new_n1152), .A4(new_n1162), .ZN(new_n1163));
  NOR3_X1   g738(.A1(new_n1067), .A2(new_n1095), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1117), .A2(new_n1120), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1166), .A2(G8), .A3(new_n1160), .ZN(new_n1167));
  AND3_X1   g742(.A1(new_n1109), .A2(G8), .A3(G168), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1165), .A2(new_n1162), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT63), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NOR3_X1   g746(.A1(new_n1121), .A2(new_n1170), .A3(new_n1148), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1166), .A2(G8), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(new_n1115), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1172), .A2(new_n1168), .A3(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1171), .A2(new_n1175), .ZN(new_n1176));
  AND3_X1   g751(.A1(new_n1165), .A2(new_n1162), .A3(new_n1167), .ZN(new_n1177));
  AND2_X1   g752(.A1(new_n1093), .A2(G171), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1111), .A2(new_n1110), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1106), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1180));
  OAI21_X1  g755(.A(KEYINPUT62), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT62), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1108), .A2(new_n1182), .A3(new_n1110), .A4(new_n1111), .ZN(new_n1183));
  NAND4_X1  g758(.A1(new_n1177), .A2(new_n1178), .A3(new_n1181), .A4(new_n1183), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1167), .A2(new_n1148), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1124), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1134), .ZN(new_n1187));
  OR2_X1    g762(.A1(G288), .A2(G1976), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1186), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1185), .B1(new_n1133), .B2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1176), .A2(new_n1184), .A3(new_n1190), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n992), .B1(new_n1164), .B2(new_n1191), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n989), .A2(new_n982), .ZN(new_n1193));
  XNOR2_X1  g768(.A(new_n1193), .B(KEYINPUT48), .ZN(new_n1194));
  INV_X1    g769(.A(new_n781), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n983), .B1(new_n972), .B2(new_n1195), .ZN(new_n1196));
  XOR2_X1   g771(.A(new_n984), .B(KEYINPUT46), .Z(new_n1197));
  NAND2_X1  g772(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  AND2_X1   g773(.A1(new_n1198), .A2(KEYINPUT47), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n1198), .A2(KEYINPUT47), .ZN(new_n1200));
  OAI22_X1  g775(.A1(new_n988), .A2(new_n1194), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n985), .A2(new_n722), .A3(new_n719), .ZN(new_n1202));
  OR2_X1    g777(.A1(new_n806), .A2(G2067), .ZN(new_n1203));
  AOI21_X1  g778(.A(new_n986), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  NOR2_X1   g779(.A1(new_n1201), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1192), .A2(new_n1205), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g781(.A1(new_n673), .A2(new_n462), .ZN(new_n1208));
  NOR2_X1   g782(.A1(G401), .A2(new_n1208), .ZN(new_n1209));
  AND4_X1   g783(.A1(new_n705), .A2(new_n904), .A3(new_n965), .A4(new_n1209), .ZN(G308));
  NAND4_X1  g784(.A1(new_n705), .A2(new_n904), .A3(new_n965), .A4(new_n1209), .ZN(G225));
endmodule


