//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 0 0 1 1 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 0 1 1 1 0 1 0 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:17 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n559, new_n561, new_n562, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n619, new_n621, new_n622, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1195, new_n1196;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT65), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(KEYINPUT67), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  XNOR2_X1  g046(.A(KEYINPUT3), .B(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(KEYINPUT67), .A3(G125), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n470), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(KEYINPUT66), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT66), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n474), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n479), .A2(new_n472), .A3(G137), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n464), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G101), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n481), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G160));
  NOR2_X1   g063(.A1(new_n468), .A2(new_n479), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n468), .A2(G2105), .ZN(new_n490));
  AOI22_X1  g065(.A1(G124), .A2(new_n489), .B1(new_n490), .B2(G136), .ZN(new_n491));
  OAI221_X1 g066(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n479), .C2(G112), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g068(.A(new_n493), .B(KEYINPUT68), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G162));
  NAND3_X1  g070(.A1(new_n479), .A2(new_n472), .A3(G138), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n465), .A2(new_n467), .A3(G126), .ZN(new_n499));
  NAND2_X1  g074(.A1(G114), .A2(G2104), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G2105), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n483), .A2(G102), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n479), .A2(new_n472), .A3(KEYINPUT4), .A4(G138), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n498), .A2(new_n502), .A3(new_n503), .A4(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  OAI21_X1  g082(.A(KEYINPUT69), .B1(new_n507), .B2(KEYINPUT6), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT69), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n509), .A2(new_n510), .A3(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n507), .A2(KEYINPUT6), .ZN(new_n513));
  AND2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n514), .A2(G50), .B1(G75), .B2(G651), .ZN(new_n515));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n512), .A2(new_n513), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n516), .A2(KEYINPUT5), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT5), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G88), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT5), .B(G543), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n525), .A2(G62), .A3(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n517), .A2(new_n527), .ZN(G166));
  NOR2_X1   g103(.A1(new_n518), .A2(new_n516), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G51), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n523), .A2(G89), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n525), .A2(G63), .A3(G651), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n530), .A2(new_n531), .A3(new_n532), .A4(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  NAND2_X1  g111(.A1(G77), .A2(G543), .ZN(new_n537));
  INV_X1    g112(.A(G64), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n537), .B1(new_n522), .B2(new_n538), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n529), .A2(G52), .B1(G651), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n523), .A2(G90), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  INV_X1    g118(.A(G56), .ZN(new_n544));
  INV_X1    g119(.A(G68), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n522), .A2(new_n544), .B1(new_n545), .B2(new_n516), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(KEYINPUT70), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT70), .ZN(new_n548));
  OAI221_X1 g123(.A(new_n548), .B1(new_n545), .B2(new_n516), .C1(new_n522), .C2(new_n544), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n547), .A2(G651), .A3(new_n549), .ZN(new_n550));
  NAND4_X1  g125(.A1(new_n512), .A2(G43), .A3(G543), .A4(new_n513), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n512), .A2(G81), .A3(new_n513), .A4(new_n525), .ZN(new_n552));
  AND2_X1   g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AND3_X1   g128(.A1(new_n550), .A2(KEYINPUT71), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g129(.A(KEYINPUT71), .B1(new_n550), .B2(new_n553), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  AND3_X1   g133(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G36), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n559), .A2(new_n562), .ZN(G188));
  AND2_X1   g138(.A1(G53), .A2(G543), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n509), .B1(new_n510), .B2(G651), .ZN(new_n565));
  NOR3_X1   g140(.A1(new_n507), .A2(KEYINPUT69), .A3(KEYINPUT6), .ZN(new_n566));
  OAI211_X1 g141(.A(new_n513), .B(new_n564), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT72), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n512), .A2(KEYINPUT72), .A3(new_n513), .A4(new_n564), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n569), .A2(KEYINPUT9), .A3(new_n570), .ZN(new_n571));
  OR2_X1    g146(.A1(new_n567), .A2(KEYINPUT9), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n571), .A2(KEYINPUT73), .A3(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT73), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n569), .A2(new_n574), .A3(KEYINPUT9), .A4(new_n570), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT74), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n525), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n577), .B2(new_n507), .ZN(new_n578));
  NAND2_X1  g153(.A1(G78), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G65), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n522), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n581), .A2(KEYINPUT74), .A3(G651), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n578), .A2(new_n582), .B1(new_n523), .B2(G91), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n573), .A2(new_n575), .A3(new_n583), .ZN(G299));
  OR2_X1    g159(.A1(new_n517), .A2(new_n527), .ZN(G303));
  NAND2_X1  g160(.A1(new_n529), .A2(G49), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n523), .A2(G87), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n525), .B2(G74), .ZN(new_n588));
  AND3_X1   g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G288));
  NAND2_X1  g165(.A1(new_n529), .A2(G48), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n523), .A2(G86), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n525), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n593), .A2(new_n507), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n591), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  XOR2_X1   g170(.A(new_n595), .B(KEYINPUT75), .Z(G305));
  NAND2_X1  g171(.A1(new_n523), .A2(G85), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n529), .A2(G47), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n525), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  OR2_X1    g174(.A1(new_n599), .A2(new_n507), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n597), .A2(new_n598), .A3(new_n600), .ZN(G290));
  NAND2_X1  g176(.A1(G301), .A2(G868), .ZN(new_n602));
  NAND2_X1  g177(.A1(G79), .A2(G543), .ZN(new_n603));
  INV_X1    g178(.A(G66), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n522), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n529), .A2(G54), .B1(G651), .B2(new_n605), .ZN(new_n606));
  NAND4_X1  g181(.A1(new_n512), .A2(G92), .A3(new_n513), .A4(new_n525), .ZN(new_n607));
  XNOR2_X1  g182(.A(KEYINPUT76), .B(KEYINPUT10), .ZN(new_n608));
  OR2_X1    g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n607), .A2(new_n608), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n606), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n602), .B1(new_n612), .B2(G868), .ZN(G284));
  OAI21_X1  g188(.A(new_n602), .B1(new_n612), .B2(G868), .ZN(G321));
  NAND2_X1  g189(.A1(G286), .A2(G868), .ZN(new_n615));
  XNOR2_X1  g190(.A(G299), .B(KEYINPUT77), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G868), .ZN(G297));
  OAI21_X1  g192(.A(new_n615), .B1(new_n616), .B2(G868), .ZN(G280));
  XNOR2_X1  g193(.A(KEYINPUT78), .B(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n612), .B1(G860), .B2(new_n619), .ZN(G148));
  NAND2_X1  g195(.A1(new_n612), .A2(new_n619), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G868), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G868), .B2(new_n557), .ZN(G323));
  XNOR2_X1  g198(.A(KEYINPUT79), .B(KEYINPUT11), .ZN(new_n624));
  XNOR2_X1  g199(.A(G323), .B(new_n624), .ZN(G282));
  NAND2_X1  g200(.A1(new_n472), .A2(new_n483), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2100), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n490), .A2(G135), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT80), .Z(new_n631));
  NAND2_X1  g206(.A1(new_n489), .A2(G123), .ZN(new_n632));
  OAI221_X1 g207(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n479), .C2(G111), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n634), .A2(G2096), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(G2096), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n629), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT81), .Z(G156));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2430), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2435), .ZN(new_n640));
  XOR2_X1   g215(.A(G2427), .B(G2438), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(KEYINPUT14), .ZN(new_n643));
  XOR2_X1   g218(.A(G2451), .B(G2454), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n643), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G1341), .B(G1348), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2443), .B(G2446), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n650), .A2(G14), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT82), .ZN(G401));
  XOR2_X1   g227(.A(G2072), .B(G2078), .Z(new_n653));
  XOR2_X1   g228(.A(G2067), .B(G2678), .Z(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n653), .B1(new_n657), .B2(KEYINPUT18), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2096), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2100), .ZN(new_n660));
  AND2_X1   g235(.A1(new_n657), .A2(KEYINPUT17), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n655), .A2(new_n656), .ZN(new_n662));
  AOI21_X1  g237(.A(KEYINPUT18), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n660), .B(new_n663), .Z(G227));
  XNOR2_X1  g239(.A(G1956), .B(G2474), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT83), .ZN(new_n666));
  XOR2_X1   g241(.A(G1961), .B(G1966), .Z(new_n667));
  AND2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G1971), .B(G1976), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT19), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(KEYINPUT20), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n666), .A2(new_n667), .ZN(new_n673));
  AOI22_X1  g248(.A1(new_n671), .A2(new_n672), .B1(new_n670), .B2(new_n673), .ZN(new_n674));
  OR3_X1    g249(.A1(new_n668), .A2(new_n673), .A3(new_n670), .ZN(new_n675));
  OAI211_X1 g250(.A(new_n674), .B(new_n675), .C1(new_n672), .C2(new_n671), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT84), .B(G1981), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n676), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1991), .B(G1996), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(G1986), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n680), .B(new_n682), .ZN(G229));
  INV_X1    g258(.A(G16), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(G21), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n685), .B1(G168), .B2(new_n684), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT94), .B(G1966), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(G29), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G35), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(G162), .B2(new_n689), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n691), .A2(new_n693), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(G2090), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(G299), .A2(G16), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n684), .A2(KEYINPUT23), .A3(G20), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT23), .ZN(new_n701));
  INV_X1    g276(.A(G20), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n701), .B1(new_n702), .B2(G16), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n699), .A2(new_n700), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(G1956), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(KEYINPUT92), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G29), .B2(G32), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n489), .A2(G129), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n490), .A2(G141), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n483), .A2(G105), .ZN(new_n711));
  NAND3_X1  g286(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT26), .Z(new_n713));
  NAND4_X1  g288(.A1(new_n709), .A2(new_n710), .A3(new_n711), .A4(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n714), .A2(new_n689), .ZN(new_n715));
  MUX2_X1   g290(.A(new_n708), .B(new_n707), .S(new_n715), .Z(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT27), .B(G1996), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT93), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n716), .B(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(KEYINPUT24), .A2(G34), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(KEYINPUT24), .A2(G34), .ZN(new_n722));
  NOR3_X1   g297(.A1(new_n721), .A2(new_n722), .A3(G29), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n487), .B2(G29), .ZN(new_n724));
  INV_X1    g299(.A(G2084), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AND2_X1   g301(.A1(new_n689), .A2(G33), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n479), .A2(G103), .A3(G2104), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT25), .Z(new_n729));
  NAND2_X1  g304(.A1(G115), .A2(G2104), .ZN(new_n730));
  INV_X1    g305(.A(G127), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(new_n468), .B2(new_n731), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n732), .A2(new_n480), .B1(new_n490), .B2(G139), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT91), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n729), .A2(KEYINPUT91), .A3(new_n733), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n727), .B1(new_n738), .B2(G29), .ZN(new_n739));
  INV_X1    g314(.A(G2072), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n724), .A2(new_n725), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n719), .A2(new_n726), .A3(new_n741), .A4(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n684), .A2(G5), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G171), .B2(new_n684), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT95), .B(G1961), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n739), .A2(new_n740), .ZN(new_n748));
  NOR3_X1   g323(.A1(new_n743), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n684), .A2(G19), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(new_n557), .B2(new_n684), .ZN(new_n751));
  INV_X1    g326(.A(G11), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n751), .A2(G1341), .B1(KEYINPUT31), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n751), .A2(G1341), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n689), .A2(G26), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  AOI22_X1  g332(.A1(G128), .A2(new_n489), .B1(new_n490), .B2(G140), .ZN(new_n758));
  OAI21_X1  g333(.A(G2104), .B1(new_n479), .B2(G116), .ZN(new_n759));
  NOR2_X1   g334(.A1(G104), .A2(G2105), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n760), .A2(KEYINPUT89), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(KEYINPUT89), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n758), .B1(new_n759), .B2(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n757), .B1(new_n764), .B2(G29), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G2067), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT30), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n767), .A2(G28), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(G28), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n768), .A2(new_n769), .A3(new_n689), .ZN(new_n770));
  INV_X1    g345(.A(G2078), .ZN(new_n771));
  NAND2_X1  g346(.A1(G164), .A2(G29), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G27), .B2(G29), .ZN(new_n773));
  OAI211_X1 g348(.A(new_n766), .B(new_n770), .C1(new_n771), .C2(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n754), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n773), .A2(new_n771), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n634), .A2(new_n689), .ZN(new_n777));
  AND4_X1   g352(.A1(new_n753), .A2(new_n775), .A3(new_n776), .A4(new_n777), .ZN(new_n778));
  NAND4_X1  g353(.A1(new_n698), .A2(new_n706), .A3(new_n749), .A4(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n684), .A2(G6), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n595), .B(KEYINPUT75), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n781), .B1(new_n782), .B2(new_n684), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT32), .B(G1981), .Z(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n684), .A2(G22), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G166), .B2(new_n684), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G1971), .ZN(new_n788));
  NOR2_X1   g363(.A1(G16), .A2(G23), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n589), .B2(G16), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT33), .B(G1976), .Z(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n788), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n785), .A2(new_n793), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT34), .Z(new_n795));
  INV_X1    g370(.A(KEYINPUT36), .ZN(new_n796));
  INV_X1    g371(.A(G24), .ZN(new_n797));
  OAI21_X1  g372(.A(KEYINPUT86), .B1(new_n797), .B2(G16), .ZN(new_n798));
  OR3_X1    g373(.A1(new_n797), .A2(KEYINPUT86), .A3(G16), .ZN(new_n799));
  INV_X1    g374(.A(G290), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n798), .B(new_n799), .C1(new_n800), .C2(new_n684), .ZN(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT87), .B(G1986), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n689), .A2(G25), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT85), .ZN(new_n805));
  INV_X1    g380(.A(new_n489), .ZN(new_n806));
  INV_X1    g381(.A(G119), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n490), .A2(G131), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n489), .A2(KEYINPUT85), .A3(G119), .ZN(new_n810));
  OAI221_X1 g385(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n479), .C2(G107), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n808), .A2(new_n809), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n804), .B1(new_n813), .B2(new_n689), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT35), .B(G1991), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AND2_X1   g391(.A1(new_n814), .A2(new_n815), .ZN(new_n817));
  NOR3_X1   g392(.A1(new_n803), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  AND3_X1   g393(.A1(new_n795), .A2(new_n796), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n796), .B1(new_n795), .B2(new_n818), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n688), .B(new_n780), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n612), .A2(G16), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(G4), .B2(G16), .ZN(new_n823));
  XOR2_X1   g398(.A(KEYINPUT88), .B(G1348), .Z(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n752), .A2(KEYINPUT31), .ZN(new_n826));
  NOR3_X1   g401(.A1(new_n821), .A2(new_n825), .A3(new_n826), .ZN(G311));
  INV_X1    g402(.A(new_n820), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n795), .A2(new_n796), .A3(new_n818), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n779), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n825), .ZN(new_n831));
  INV_X1    g406(.A(new_n826), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n830), .A2(new_n831), .A3(new_n832), .A4(new_n688), .ZN(G150));
  NAND2_X1  g408(.A1(new_n523), .A2(G93), .ZN(new_n834));
  AOI22_X1  g409(.A1(new_n525), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n835), .A2(new_n507), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n514), .A2(G55), .A3(G543), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n834), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(G860), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(KEYINPUT37), .Z(new_n840));
  OAI211_X1 g415(.A(KEYINPUT98), .B(new_n838), .C1(new_n554), .C2(new_n555), .ZN(new_n841));
  AND3_X1   g416(.A1(new_n834), .A2(new_n836), .A3(new_n837), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n550), .A2(new_n553), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT71), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n550), .A2(KEYINPUT71), .A3(new_n553), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n842), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT98), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(new_n842), .B2(new_n843), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n841), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n612), .A2(G559), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT39), .Z(new_n854));
  XNOR2_X1  g429(.A(new_n852), .B(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n840), .B1(new_n855), .B2(G860), .ZN(G145));
  INV_X1    g431(.A(KEYINPUT99), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n736), .A2(new_n857), .A3(new_n737), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n764), .B(new_n505), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n858), .A2(new_n859), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n714), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n862), .ZN(new_n864));
  INV_X1    g439(.A(new_n714), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n864), .A2(new_n865), .A3(new_n860), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT100), .ZN(new_n868));
  INV_X1    g443(.A(G130), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n868), .B1(new_n806), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n490), .A2(G142), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n489), .A2(KEYINPUT100), .A3(G130), .ZN(new_n872));
  OAI221_X1 g447(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n479), .C2(G118), .ZN(new_n873));
  NAND4_X1  g448(.A1(new_n870), .A2(new_n871), .A3(new_n872), .A4(new_n873), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n874), .B(new_n627), .Z(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(new_n812), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n867), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n863), .A2(new_n866), .A3(new_n876), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n878), .A2(new_n879), .A3(KEYINPUT101), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n634), .B(new_n487), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(new_n494), .ZN(new_n882));
  OAI211_X1 g457(.A(new_n880), .B(new_n882), .C1(KEYINPUT101), .C2(new_n878), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n878), .A2(new_n879), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n884), .A2(new_n882), .ZN(new_n885));
  INV_X1    g460(.A(G37), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n883), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(KEYINPUT102), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT102), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n883), .A2(new_n885), .A3(new_n889), .A4(new_n886), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT40), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n888), .A2(KEYINPUT40), .A3(new_n890), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(G395));
  NAND2_X1  g470(.A1(new_n611), .A2(KEYINPUT103), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT103), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n606), .A2(new_n897), .A3(new_n609), .A4(new_n610), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n896), .A2(G299), .A3(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  NOR3_X1   g475(.A1(G299), .A2(KEYINPUT103), .A3(new_n611), .ZN(new_n901));
  OAI21_X1  g476(.A(KEYINPUT41), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OR3_X1    g477(.A1(G299), .A2(KEYINPUT103), .A3(new_n611), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT41), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n903), .A2(new_n904), .A3(new_n899), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT105), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n902), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n903), .A2(new_n899), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n908), .A2(KEYINPUT105), .A3(KEYINPUT41), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT104), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n911), .B1(new_n900), .B2(new_n901), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n903), .A2(KEYINPUT104), .A3(new_n899), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  XOR2_X1   g489(.A(new_n850), .B(new_n621), .Z(new_n915));
  MUX2_X1   g490(.A(new_n910), .B(new_n914), .S(new_n915), .Z(new_n916));
  NAND2_X1  g491(.A1(G303), .A2(new_n589), .ZN(new_n917));
  NAND2_X1  g492(.A1(G288), .A2(G166), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(new_n782), .ZN(new_n920));
  NAND3_X1  g495(.A1(G305), .A2(new_n918), .A3(new_n917), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n920), .A2(new_n921), .A3(new_n800), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n800), .B1(new_n920), .B2(new_n921), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n924), .B(KEYINPUT42), .ZN(new_n925));
  OR2_X1    g500(.A1(new_n916), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n916), .A2(new_n925), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n926), .A2(new_n927), .A3(G868), .ZN(new_n928));
  OAI21_X1  g503(.A(KEYINPUT106), .B1(new_n842), .B2(G868), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT106), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n930), .B1(new_n931), .B2(new_n928), .ZN(G295));
  OAI21_X1  g507(.A(new_n930), .B1(new_n931), .B2(new_n928), .ZN(G331));
  NAND2_X1  g508(.A1(new_n920), .A2(new_n921), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(G290), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n920), .A2(new_n921), .A3(new_n800), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(G286), .B(G301), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n938), .B(new_n841), .C1(new_n847), .C2(new_n849), .ZN(new_n939));
  XOR2_X1   g514(.A(G286), .B(G301), .Z(new_n940));
  NAND2_X1  g515(.A1(new_n850), .A2(new_n940), .ZN(new_n941));
  AOI22_X1  g516(.A1(new_n907), .A2(new_n909), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n939), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n943), .B1(new_n903), .B2(new_n899), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n937), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n945), .A2(new_n886), .ZN(new_n946));
  AND2_X1   g521(.A1(new_n941), .A2(new_n939), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT109), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n947), .A2(new_n948), .A3(new_n913), .A4(new_n912), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n902), .A2(new_n905), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n943), .ZN(new_n951));
  OAI21_X1  g526(.A(KEYINPUT109), .B1(new_n914), .B2(new_n943), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n949), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(new_n924), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n946), .A2(KEYINPUT43), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n910), .A2(new_n943), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT107), .ZN(new_n957));
  NOR3_X1   g532(.A1(new_n922), .A2(new_n923), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n947), .A2(new_n908), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n956), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n935), .A2(KEYINPUT107), .A3(new_n936), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n961), .B1(new_n942), .B2(new_n944), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n960), .A2(new_n962), .A3(new_n886), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT43), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT44), .B1(new_n955), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT108), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT108), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n963), .A2(new_n969), .A3(KEYINPUT43), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n954), .A2(new_n964), .A3(new_n886), .A4(new_n945), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT110), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n946), .A2(KEYINPUT110), .A3(new_n964), .A4(new_n954), .ZN(new_n974));
  AOI22_X1  g549(.A1(new_n968), .A2(new_n970), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n966), .B1(new_n975), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g551(.A(KEYINPUT54), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT111), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT50), .ZN(new_n979));
  INV_X1    g554(.A(G1384), .ZN(new_n980));
  AND3_X1   g555(.A1(new_n505), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n979), .B1(new_n505), .B2(new_n980), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n978), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G40), .ZN(new_n984));
  AOI211_X1 g559(.A(new_n984), .B(new_n485), .C1(new_n474), .C2(new_n480), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n505), .A2(new_n979), .A3(new_n980), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(KEYINPUT111), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n983), .A2(new_n985), .A3(new_n987), .ZN(new_n988));
  XNOR2_X1  g563(.A(KEYINPUT124), .B(G1961), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT53), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n498), .A2(new_n504), .ZN(new_n991));
  AOI22_X1  g566(.A1(new_n472), .A2(G126), .B1(G114), .B2(G2104), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n503), .B1(new_n992), .B2(new_n475), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n980), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT45), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n505), .A2(KEYINPUT45), .A3(new_n980), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n996), .A2(new_n771), .A3(new_n985), .A4(new_n997), .ZN(new_n998));
  AOI22_X1  g573(.A1(new_n988), .A2(new_n989), .B1(new_n990), .B2(new_n998), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n505), .A2(KEYINPUT45), .A3(new_n980), .ZN(new_n1000));
  AOI21_X1  g575(.A(KEYINPUT45), .B1(new_n505), .B2(new_n980), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n485), .A2(KEYINPUT125), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  NOR3_X1   g578(.A1(new_n1000), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT126), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n984), .B1(new_n474), .B2(new_n480), .ZN(new_n1006));
  OAI211_X1 g581(.A(KEYINPUT53), .B(new_n771), .C1(new_n485), .C2(KEYINPUT125), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .A4(new_n1008), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n996), .A2(new_n1006), .A3(new_n997), .A4(new_n1002), .ZN(new_n1010));
  OAI21_X1  g585(.A(KEYINPUT126), .B1(new_n1010), .B2(new_n1007), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  AND3_X1   g587(.A1(new_n999), .A2(G301), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1006), .A2(new_n486), .ZN(new_n1014));
  NOR3_X1   g589(.A1(new_n1000), .A2(new_n1001), .A3(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1015), .A2(KEYINPUT53), .A3(new_n771), .ZN(new_n1016));
  AOI21_X1  g591(.A(G301), .B1(new_n999), .B2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n977), .B1(new_n1013), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT61), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT119), .ZN(new_n1020));
  NAND2_X1  g595(.A1(G299), .A2(KEYINPUT118), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT118), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n573), .A2(new_n1022), .A3(new_n575), .A4(new_n583), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT57), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1021), .A2(KEYINPUT57), .A3(new_n1023), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g603(.A(KEYINPUT56), .B(G2072), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n994), .A2(KEYINPUT50), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1030), .A2(new_n985), .A3(new_n986), .ZN(new_n1031));
  INV_X1    g606(.A(G1956), .ZN(new_n1032));
  AOI22_X1  g607(.A1(new_n1015), .A2(new_n1029), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1020), .B1(new_n1028), .B2(new_n1033), .ZN(new_n1034));
  AND3_X1   g609(.A1(new_n1021), .A2(KEYINPUT57), .A3(new_n1023), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT57), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n1020), .B(new_n1033), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1019), .B1(new_n1034), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1018), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT127), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n999), .A2(new_n1012), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n977), .B1(new_n1042), .B2(G171), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n999), .A2(G301), .A3(new_n1016), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1041), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n983), .A2(new_n725), .A3(new_n985), .A4(new_n987), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n996), .A2(new_n985), .A3(new_n997), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(new_n687), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(G8), .ZN(new_n1050));
  INV_X1    g625(.A(G8), .ZN(new_n1051));
  NOR2_X1   g626(.A1(G168), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1050), .A2(KEYINPUT123), .A3(KEYINPUT51), .A4(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1049), .A2(G8), .A3(G286), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT51), .B1(new_n1052), .B2(KEYINPUT123), .ZN(new_n1056));
  OAI211_X1 g631(.A(G8), .B(new_n1056), .C1(new_n1049), .C2(G286), .ZN(new_n1057));
  AND3_X1   g632(.A1(new_n1054), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1058));
  NOR3_X1   g633(.A1(new_n1040), .A2(new_n1045), .A3(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G1996), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n996), .A2(new_n1060), .A3(new_n985), .A4(new_n997), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT120), .ZN(new_n1062));
  XOR2_X1   g637(.A(KEYINPUT58), .B(G1341), .Z(new_n1063));
  OAI21_X1  g638(.A(new_n1063), .B1(new_n1014), .B2(new_n994), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1061), .A2(new_n1062), .A3(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1062), .B1(new_n1061), .B2(new_n1064), .ZN(new_n1066));
  NOR3_X1   g641(.A1(new_n1065), .A2(new_n1066), .A3(new_n556), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT59), .ZN(new_n1068));
  OAI21_X1  g643(.A(KEYINPUT121), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT122), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1061), .A2(new_n1064), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT120), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1061), .A2(new_n1062), .A3(new_n1064), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1072), .A2(new_n557), .A3(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1070), .B1(new_n1074), .B2(KEYINPUT59), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1076), .A2(KEYINPUT122), .A3(new_n1068), .A4(new_n557), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT121), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1074), .A2(new_n1078), .A3(KEYINPUT59), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1069), .A2(new_n1075), .A3(new_n1077), .A4(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1033), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n996), .A2(new_n985), .A3(new_n997), .A4(new_n1029), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1026), .A2(new_n1084), .A3(new_n1027), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1081), .A2(new_n1085), .A3(KEYINPUT61), .ZN(new_n1086));
  INV_X1    g661(.A(G1348), .ZN(new_n1087));
  INV_X1    g662(.A(G2067), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1014), .A2(new_n994), .ZN(new_n1089));
  AOI22_X1  g664(.A1(new_n988), .A2(new_n1087), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT60), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1090), .A2(new_n1091), .A3(new_n612), .ZN(new_n1092));
  AND2_X1   g667(.A1(new_n1086), .A2(new_n1092), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n1090), .A2(new_n611), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1090), .A2(new_n611), .ZN(new_n1095));
  OAI21_X1  g670(.A(KEYINPUT60), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1080), .A2(new_n1093), .A3(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1034), .A2(new_n1038), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1085), .B1(new_n611), .B2(new_n1090), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(G303), .A2(G8), .ZN(new_n1102));
  XOR2_X1   g677(.A(new_n1102), .B(KEYINPUT55), .Z(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  OR2_X1    g679(.A1(new_n1015), .A2(G1971), .ZN(new_n1105));
  AND2_X1   g680(.A1(new_n1031), .A2(KEYINPUT116), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n697), .B1(new_n1031), .B2(KEYINPUT116), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1105), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  AND2_X1   g683(.A1(new_n1108), .A2(KEYINPUT117), .ZN(new_n1109));
  OAI21_X1  g684(.A(G8), .B1(new_n1108), .B2(KEYINPUT117), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1104), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  OR3_X1    g686(.A1(new_n988), .A2(KEYINPUT112), .A3(G2090), .ZN(new_n1112));
  OAI21_X1  g687(.A(KEYINPUT112), .B1(new_n988), .B2(G2090), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1112), .A2(new_n1105), .A3(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1114), .A2(G8), .A3(new_n1103), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n595), .A2(G1981), .ZN(new_n1116));
  INV_X1    g691(.A(G1981), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n591), .A2(new_n592), .A3(new_n1117), .A4(new_n594), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1118), .A2(KEYINPUT114), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1118), .A2(KEYINPUT114), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1116), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT49), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1089), .A2(new_n1051), .ZN(new_n1124));
  OAI211_X1 g699(.A(KEYINPUT49), .B(new_n1116), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1123), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(G1976), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1124), .B1(new_n1127), .B2(G288), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT52), .ZN(new_n1129));
  XNOR2_X1  g704(.A(KEYINPUT113), .B(G1976), .ZN(new_n1130));
  AOI21_X1  g705(.A(KEYINPUT52), .B1(G288), .B2(new_n1130), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1131), .B(new_n1124), .C1(new_n1127), .C2(G288), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1126), .A2(new_n1129), .A3(new_n1132), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1111), .A2(new_n1115), .A3(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1043), .A2(new_n1041), .A3(new_n1044), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1059), .A2(new_n1101), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1054), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1137));
  OR2_X1    g712(.A1(new_n1137), .A2(KEYINPUT62), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(KEYINPUT62), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1134), .A2(new_n1138), .A3(new_n1139), .A4(new_n1017), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1050), .A2(G286), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1111), .A2(new_n1115), .A3(new_n1133), .A4(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT63), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1114), .A2(G8), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1143), .B1(new_n1145), .B2(new_n1104), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1146), .A2(new_n1115), .A3(new_n1133), .A4(new_n1141), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1144), .A2(new_n1147), .ZN(new_n1148));
  AND3_X1   g723(.A1(new_n1126), .A2(new_n1127), .A3(new_n589), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1124), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1133), .A2(G8), .A3(new_n1103), .A4(new_n1114), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT115), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1153), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1136), .A2(new_n1140), .A3(new_n1148), .A4(new_n1156), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n996), .A2(new_n1014), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n764), .B(new_n1088), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n714), .B(G1996), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n812), .A2(new_n815), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n812), .A2(new_n815), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1162), .A2(new_n1163), .A3(new_n1165), .ZN(new_n1166));
  AND2_X1   g741(.A1(G290), .A2(G1986), .ZN(new_n1167));
  OR2_X1    g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g743(.A1(G290), .A2(G1986), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1158), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1157), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1158), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1173));
  OR2_X1    g748(.A1(new_n764), .A2(G2067), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1172), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1158), .B1(new_n1160), .B2(new_n714), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT46), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1177), .B1(new_n1172), .B2(G1996), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1158), .A2(KEYINPUT46), .A3(new_n1060), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1176), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  XOR2_X1   g755(.A(new_n1180), .B(KEYINPUT47), .Z(new_n1181));
  NAND2_X1  g756(.A1(new_n1166), .A2(new_n1158), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1158), .A2(new_n1169), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1183), .B(KEYINPUT48), .ZN(new_n1184));
  AOI211_X1 g759(.A(new_n1175), .B(new_n1181), .C1(new_n1182), .C2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1171), .A2(new_n1185), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g761(.A1(G229), .A2(new_n461), .ZN(new_n1188));
  INV_X1    g762(.A(new_n1188), .ZN(new_n1189));
  AOI21_X1  g763(.A(G227), .B1(new_n650), .B2(G14), .ZN(new_n1190));
  NAND2_X1  g764(.A1(new_n887), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g765(.A1(new_n968), .A2(new_n970), .ZN(new_n1192));
  NAND2_X1  g766(.A1(new_n973), .A2(new_n974), .ZN(new_n1193));
  AOI211_X1 g767(.A(new_n1189), .B(new_n1191), .C1(new_n1192), .C2(new_n1193), .ZN(G308));
  NAND2_X1  g768(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1195));
  INV_X1    g769(.A(new_n1191), .ZN(new_n1196));
  NAND3_X1  g770(.A1(new_n1195), .A2(new_n1188), .A3(new_n1196), .ZN(G225));
endmodule


