

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X2 U546 ( .A(n733), .ZN(n700) );
  NOR2_X2 U547 ( .A1(G2105), .A2(n521), .ZN(n894) );
  NOR2_X1 U548 ( .A1(G543), .A2(G651), .ZN(n640) );
  XNOR2_X2 U549 ( .A(n741), .B(KEYINPUT32), .ZN(n765) );
  NOR2_X1 U550 ( .A1(G164), .A2(G1384), .ZN(n781) );
  BUF_X2 U551 ( .A(n895), .Z(n512) );
  XOR2_X1 U552 ( .A(KEYINPUT17), .B(n518), .Z(n895) );
  INV_X1 U553 ( .A(KEYINPUT108), .ZN(n731) );
  XNOR2_X1 U554 ( .A(n732), .B(n731), .ZN(n742) );
  NOR2_X1 U555 ( .A1(n655), .A2(G651), .ZN(n648) );
  INV_X1 U556 ( .A(G2104), .ZN(n521) );
  INV_X1 U557 ( .A(G2105), .ZN(n513) );
  NOR2_X2 U558 ( .A1(n521), .A2(n513), .ZN(n890) );
  NAND2_X1 U559 ( .A1(G114), .A2(n890), .ZN(n515) );
  NOR2_X2 U560 ( .A1(G2104), .A2(n513), .ZN(n891) );
  NAND2_X1 U561 ( .A1(G126), .A2(n891), .ZN(n514) );
  NAND2_X1 U562 ( .A1(n515), .A2(n514), .ZN(n517) );
  INV_X1 U563 ( .A(KEYINPUT88), .ZN(n516) );
  XNOR2_X1 U564 ( .A(n517), .B(n516), .ZN(n520) );
  NOR2_X1 U565 ( .A1(G2104), .A2(G2105), .ZN(n518) );
  NAND2_X1 U566 ( .A1(n512), .A2(G138), .ZN(n519) );
  NAND2_X1 U567 ( .A1(n520), .A2(n519), .ZN(n524) );
  NAND2_X1 U568 ( .A1(G102), .A2(n894), .ZN(n522) );
  XNOR2_X1 U569 ( .A(KEYINPUT89), .B(n522), .ZN(n523) );
  NOR2_X2 U570 ( .A1(n524), .A2(n523), .ZN(G164) );
  NAND2_X1 U571 ( .A1(n890), .A2(G113), .ZN(n527) );
  NAND2_X1 U572 ( .A1(G101), .A2(n894), .ZN(n525) );
  XOR2_X1 U573 ( .A(KEYINPUT23), .B(n525), .Z(n526) );
  NAND2_X1 U574 ( .A1(n527), .A2(n526), .ZN(n531) );
  NAND2_X1 U575 ( .A1(G125), .A2(n891), .ZN(n529) );
  NAND2_X1 U576 ( .A1(G137), .A2(n512), .ZN(n528) );
  NAND2_X1 U577 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X2 U578 ( .A1(n531), .A2(n530), .ZN(G160) );
  XOR2_X1 U579 ( .A(G2443), .B(G2446), .Z(n533) );
  XNOR2_X1 U580 ( .A(G2427), .B(G2451), .ZN(n532) );
  XNOR2_X1 U581 ( .A(n533), .B(n532), .ZN(n539) );
  XOR2_X1 U582 ( .A(G2430), .B(G2454), .Z(n535) );
  XNOR2_X1 U583 ( .A(G1348), .B(G1341), .ZN(n534) );
  XNOR2_X1 U584 ( .A(n535), .B(n534), .ZN(n537) );
  XOR2_X1 U585 ( .A(G2435), .B(G2438), .Z(n536) );
  XNOR2_X1 U586 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U587 ( .A(n539), .B(n538), .Z(n540) );
  AND2_X1 U588 ( .A1(G14), .A2(n540), .ZN(G401) );
  AND2_X1 U589 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U590 ( .A1(G111), .A2(n890), .ZN(n542) );
  NAND2_X1 U591 ( .A1(G99), .A2(n894), .ZN(n541) );
  NAND2_X1 U592 ( .A1(n542), .A2(n541), .ZN(n548) );
  NAND2_X1 U593 ( .A1(G135), .A2(n512), .ZN(n543) );
  XNOR2_X1 U594 ( .A(n543), .B(KEYINPUT78), .ZN(n546) );
  NAND2_X1 U595 ( .A1(G123), .A2(n891), .ZN(n544) );
  XNOR2_X1 U596 ( .A(n544), .B(KEYINPUT18), .ZN(n545) );
  NAND2_X1 U597 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U598 ( .A1(n548), .A2(n547), .ZN(n967) );
  XNOR2_X1 U599 ( .A(n967), .B(G2096), .ZN(n549) );
  XNOR2_X1 U600 ( .A(n549), .B(KEYINPUT79), .ZN(n550) );
  OR2_X1 U601 ( .A1(G2100), .A2(n550), .ZN(G156) );
  INV_X1 U602 ( .A(G57), .ZN(G237) );
  INV_X1 U603 ( .A(G651), .ZN(n555) );
  NOR2_X1 U604 ( .A1(G543), .A2(n555), .ZN(n551) );
  XOR2_X1 U605 ( .A(KEYINPUT1), .B(n551), .Z(n651) );
  NAND2_X1 U606 ( .A1(G63), .A2(n651), .ZN(n553) );
  XOR2_X1 U607 ( .A(KEYINPUT0), .B(G543), .Z(n655) );
  NAND2_X1 U608 ( .A1(G51), .A2(n648), .ZN(n552) );
  NAND2_X1 U609 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U610 ( .A(KEYINPUT6), .B(n554), .Z(n563) );
  NOR2_X1 U611 ( .A1(n655), .A2(n555), .ZN(n638) );
  NAND2_X1 U612 ( .A1(G76), .A2(n638), .ZN(n559) );
  XOR2_X1 U613 ( .A(KEYINPUT4), .B(KEYINPUT73), .Z(n557) );
  NAND2_X1 U614 ( .A1(G89), .A2(n640), .ZN(n556) );
  XNOR2_X1 U615 ( .A(n557), .B(n556), .ZN(n558) );
  NAND2_X1 U616 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U617 ( .A(n560), .B(KEYINPUT74), .ZN(n561) );
  XNOR2_X1 U618 ( .A(KEYINPUT5), .B(n561), .ZN(n562) );
  NAND2_X1 U619 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U620 ( .A(KEYINPUT7), .B(n564), .ZN(G168) );
  XOR2_X1 U621 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U622 ( .A1(G7), .A2(G661), .ZN(n565) );
  XNOR2_X1 U623 ( .A(n565), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U624 ( .A(G223), .ZN(n831) );
  NAND2_X1 U625 ( .A1(n831), .A2(G567), .ZN(n566) );
  XNOR2_X1 U626 ( .A(n566), .B(KEYINPUT69), .ZN(n567) );
  XNOR2_X1 U627 ( .A(KEYINPUT11), .B(n567), .ZN(G234) );
  XOR2_X1 U628 ( .A(G860), .B(KEYINPUT72), .Z(n605) );
  NAND2_X1 U629 ( .A1(G56), .A2(n651), .ZN(n568) );
  XNOR2_X1 U630 ( .A(n568), .B(KEYINPUT14), .ZN(n571) );
  NAND2_X1 U631 ( .A1(G43), .A2(n648), .ZN(n569) );
  XOR2_X1 U632 ( .A(KEYINPUT71), .B(n569), .Z(n570) );
  NAND2_X1 U633 ( .A1(n571), .A2(n570), .ZN(n578) );
  NAND2_X1 U634 ( .A1(G81), .A2(n640), .ZN(n572) );
  XNOR2_X1 U635 ( .A(n572), .B(KEYINPUT70), .ZN(n573) );
  XNOR2_X1 U636 ( .A(n573), .B(KEYINPUT12), .ZN(n575) );
  NAND2_X1 U637 ( .A1(G68), .A2(n638), .ZN(n574) );
  NAND2_X1 U638 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U639 ( .A(KEYINPUT13), .B(n576), .Z(n577) );
  NOR2_X1 U640 ( .A1(n578), .A2(n577), .ZN(n988) );
  INV_X1 U641 ( .A(n988), .ZN(n611) );
  OR2_X1 U642 ( .A1(n605), .A2(n611), .ZN(G153) );
  NAND2_X1 U643 ( .A1(n638), .A2(G77), .ZN(n579) );
  XOR2_X1 U644 ( .A(KEYINPUT67), .B(n579), .Z(n581) );
  NAND2_X1 U645 ( .A1(n640), .A2(G90), .ZN(n580) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(KEYINPUT9), .B(n582), .ZN(n586) );
  NAND2_X1 U648 ( .A1(G64), .A2(n651), .ZN(n584) );
  NAND2_X1 U649 ( .A1(G52), .A2(n648), .ZN(n583) );
  AND2_X1 U650 ( .A1(n584), .A2(n583), .ZN(n585) );
  NAND2_X1 U651 ( .A1(n586), .A2(n585), .ZN(G301) );
  NAND2_X1 U652 ( .A1(G868), .A2(G301), .ZN(n595) );
  NAND2_X1 U653 ( .A1(G79), .A2(n638), .ZN(n588) );
  NAND2_X1 U654 ( .A1(G92), .A2(n640), .ZN(n587) );
  NAND2_X1 U655 ( .A1(n588), .A2(n587), .ZN(n592) );
  NAND2_X1 U656 ( .A1(G66), .A2(n651), .ZN(n590) );
  NAND2_X1 U657 ( .A1(G54), .A2(n648), .ZN(n589) );
  NAND2_X1 U658 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U659 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U660 ( .A(n593), .B(KEYINPUT15), .ZN(n987) );
  INV_X1 U661 ( .A(G868), .ZN(n667) );
  NAND2_X1 U662 ( .A1(n987), .A2(n667), .ZN(n594) );
  NAND2_X1 U663 ( .A1(n595), .A2(n594), .ZN(G284) );
  NAND2_X1 U664 ( .A1(G65), .A2(n651), .ZN(n597) );
  NAND2_X1 U665 ( .A1(G53), .A2(n648), .ZN(n596) );
  NAND2_X1 U666 ( .A1(n597), .A2(n596), .ZN(n601) );
  NAND2_X1 U667 ( .A1(G78), .A2(n638), .ZN(n599) );
  NAND2_X1 U668 ( .A1(G91), .A2(n640), .ZN(n598) );
  NAND2_X1 U669 ( .A1(n599), .A2(n598), .ZN(n600) );
  NOR2_X1 U670 ( .A1(n601), .A2(n600), .ZN(n984) );
  XOR2_X1 U671 ( .A(n984), .B(KEYINPUT68), .Z(G299) );
  NOR2_X1 U672 ( .A1(G868), .A2(G299), .ZN(n602) );
  XOR2_X1 U673 ( .A(KEYINPUT75), .B(n602), .Z(n604) );
  NOR2_X1 U674 ( .A1(G286), .A2(n667), .ZN(n603) );
  NOR2_X1 U675 ( .A1(n604), .A2(n603), .ZN(G297) );
  NAND2_X1 U676 ( .A1(G559), .A2(n605), .ZN(n606) );
  XNOR2_X1 U677 ( .A(KEYINPUT76), .B(n606), .ZN(n607) );
  INV_X1 U678 ( .A(n987), .ZN(n838) );
  NAND2_X1 U679 ( .A1(n607), .A2(n838), .ZN(n608) );
  XNOR2_X1 U680 ( .A(KEYINPUT16), .B(n608), .ZN(G148) );
  NOR2_X1 U681 ( .A1(n987), .A2(n667), .ZN(n609) );
  XNOR2_X1 U682 ( .A(n609), .B(KEYINPUT77), .ZN(n610) );
  NOR2_X1 U683 ( .A1(G559), .A2(n610), .ZN(n613) );
  NOR2_X1 U684 ( .A1(G868), .A2(n611), .ZN(n612) );
  NOR2_X1 U685 ( .A1(n613), .A2(n612), .ZN(G282) );
  NAND2_X1 U686 ( .A1(G559), .A2(n838), .ZN(n614) );
  XOR2_X1 U687 ( .A(n988), .B(n614), .Z(n664) );
  NOR2_X1 U688 ( .A1(n664), .A2(G860), .ZN(n623) );
  NAND2_X1 U689 ( .A1(G93), .A2(n640), .ZN(n616) );
  NAND2_X1 U690 ( .A1(G67), .A2(n651), .ZN(n615) );
  NAND2_X1 U691 ( .A1(n616), .A2(n615), .ZN(n619) );
  NAND2_X1 U692 ( .A1(G55), .A2(n648), .ZN(n617) );
  XNOR2_X1 U693 ( .A(KEYINPUT81), .B(n617), .ZN(n618) );
  NOR2_X1 U694 ( .A1(n619), .A2(n618), .ZN(n621) );
  NAND2_X1 U695 ( .A1(n638), .A2(G80), .ZN(n620) );
  NAND2_X1 U696 ( .A1(n621), .A2(n620), .ZN(n666) );
  XOR2_X1 U697 ( .A(n666), .B(KEYINPUT80), .Z(n622) );
  XNOR2_X1 U698 ( .A(n623), .B(n622), .ZN(G145) );
  NAND2_X1 U699 ( .A1(G75), .A2(n638), .ZN(n625) );
  NAND2_X1 U700 ( .A1(G88), .A2(n640), .ZN(n624) );
  NAND2_X1 U701 ( .A1(n625), .A2(n624), .ZN(n629) );
  NAND2_X1 U702 ( .A1(G62), .A2(n651), .ZN(n627) );
  NAND2_X1 U703 ( .A1(G50), .A2(n648), .ZN(n626) );
  NAND2_X1 U704 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U705 ( .A1(n629), .A2(n628), .ZN(G166) );
  XOR2_X1 U706 ( .A(KEYINPUT84), .B(KEYINPUT2), .Z(n631) );
  NAND2_X1 U707 ( .A1(G73), .A2(n638), .ZN(n630) );
  XNOR2_X1 U708 ( .A(n631), .B(n630), .ZN(n635) );
  NAND2_X1 U709 ( .A1(G61), .A2(n651), .ZN(n633) );
  NAND2_X1 U710 ( .A1(G48), .A2(n648), .ZN(n632) );
  NAND2_X1 U711 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U712 ( .A1(n635), .A2(n634), .ZN(n637) );
  NAND2_X1 U713 ( .A1(n640), .A2(G86), .ZN(n636) );
  NAND2_X1 U714 ( .A1(n637), .A2(n636), .ZN(G305) );
  NAND2_X1 U715 ( .A1(n638), .A2(G72), .ZN(n639) );
  XOR2_X1 U716 ( .A(KEYINPUT65), .B(n639), .Z(n642) );
  NAND2_X1 U717 ( .A1(n640), .A2(G85), .ZN(n641) );
  NAND2_X1 U718 ( .A1(n642), .A2(n641), .ZN(n643) );
  XOR2_X1 U719 ( .A(KEYINPUT66), .B(n643), .Z(n647) );
  NAND2_X1 U720 ( .A1(G60), .A2(n651), .ZN(n645) );
  NAND2_X1 U721 ( .A1(G47), .A2(n648), .ZN(n644) );
  AND2_X1 U722 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U723 ( .A1(n647), .A2(n646), .ZN(G290) );
  NAND2_X1 U724 ( .A1(n648), .A2(G49), .ZN(n649) );
  XOR2_X1 U725 ( .A(KEYINPUT82), .B(n649), .Z(n650) );
  NOR2_X1 U726 ( .A1(n651), .A2(n650), .ZN(n653) );
  NAND2_X1 U727 ( .A1(G651), .A2(G74), .ZN(n652) );
  NAND2_X1 U728 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U729 ( .A(n654), .B(KEYINPUT83), .ZN(n657) );
  NAND2_X1 U730 ( .A1(G87), .A2(n655), .ZN(n656) );
  NAND2_X1 U731 ( .A1(n657), .A2(n656), .ZN(G288) );
  XOR2_X1 U732 ( .A(G299), .B(KEYINPUT19), .Z(n659) );
  XNOR2_X1 U733 ( .A(G166), .B(KEYINPUT85), .ZN(n658) );
  XNOR2_X1 U734 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U735 ( .A(n660), .B(G305), .ZN(n661) );
  XNOR2_X1 U736 ( .A(n661), .B(n666), .ZN(n662) );
  XNOR2_X1 U737 ( .A(n662), .B(G290), .ZN(n663) );
  XNOR2_X1 U738 ( .A(n663), .B(G288), .ZN(n837) );
  XNOR2_X1 U739 ( .A(n664), .B(n837), .ZN(n665) );
  NAND2_X1 U740 ( .A1(n665), .A2(G868), .ZN(n669) );
  NAND2_X1 U741 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U742 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U743 ( .A(KEYINPUT86), .B(n670), .ZN(G295) );
  NAND2_X1 U744 ( .A1(G2078), .A2(G2084), .ZN(n671) );
  XOR2_X1 U745 ( .A(KEYINPUT20), .B(n671), .Z(n672) );
  NAND2_X1 U746 ( .A1(G2090), .A2(n672), .ZN(n673) );
  XNOR2_X1 U747 ( .A(KEYINPUT21), .B(n673), .ZN(n674) );
  NAND2_X1 U748 ( .A1(n674), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U749 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U750 ( .A(KEYINPUT87), .B(KEYINPUT22), .Z(n676) );
  NAND2_X1 U751 ( .A1(G132), .A2(G82), .ZN(n675) );
  XNOR2_X1 U752 ( .A(n676), .B(n675), .ZN(n677) );
  NOR2_X1 U753 ( .A1(n677), .A2(G218), .ZN(n678) );
  NAND2_X1 U754 ( .A1(G96), .A2(n678), .ZN(n835) );
  NAND2_X1 U755 ( .A1(n835), .A2(G2106), .ZN(n682) );
  NAND2_X1 U756 ( .A1(G69), .A2(G120), .ZN(n679) );
  NOR2_X1 U757 ( .A1(G237), .A2(n679), .ZN(n680) );
  NAND2_X1 U758 ( .A1(G108), .A2(n680), .ZN(n836) );
  NAND2_X1 U759 ( .A1(n836), .A2(G567), .ZN(n681) );
  NAND2_X1 U760 ( .A1(n682), .A2(n681), .ZN(n914) );
  NAND2_X1 U761 ( .A1(G483), .A2(G661), .ZN(n683) );
  NOR2_X1 U762 ( .A1(n914), .A2(n683), .ZN(n834) );
  NAND2_X1 U763 ( .A1(n834), .A2(G36), .ZN(G176) );
  INV_X1 U764 ( .A(G166), .ZN(G303) );
  INV_X1 U765 ( .A(G301), .ZN(G171) );
  NAND2_X1 U766 ( .A1(G160), .A2(G40), .ZN(n780) );
  INV_X1 U767 ( .A(n780), .ZN(n685) );
  NAND2_X2 U768 ( .A1(n781), .A2(n685), .ZN(n733) );
  XNOR2_X1 U769 ( .A(G1961), .B(KEYINPUT97), .ZN(n915) );
  NAND2_X1 U770 ( .A1(n733), .A2(n915), .ZN(n687) );
  XNOR2_X1 U771 ( .A(KEYINPUT25), .B(G2078), .ZN(n951) );
  NAND2_X1 U772 ( .A1(n700), .A2(n951), .ZN(n686) );
  NAND2_X1 U773 ( .A1(n687), .A2(n686), .ZN(n724) );
  NOR2_X1 U774 ( .A1(G171), .A2(n724), .ZN(n693) );
  NAND2_X1 U775 ( .A1(G8), .A2(n733), .ZN(n773) );
  NOR2_X1 U776 ( .A1(G1966), .A2(n773), .ZN(n743) );
  NOR2_X1 U777 ( .A1(G2084), .A2(n733), .ZN(n745) );
  NOR2_X1 U778 ( .A1(n743), .A2(n745), .ZN(n688) );
  XOR2_X1 U779 ( .A(KEYINPUT107), .B(n688), .Z(n689) );
  NAND2_X1 U780 ( .A1(G8), .A2(n689), .ZN(n690) );
  XNOR2_X1 U781 ( .A(KEYINPUT30), .B(n690), .ZN(n691) );
  NOR2_X1 U782 ( .A1(G168), .A2(n691), .ZN(n692) );
  NOR2_X1 U783 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U784 ( .A(KEYINPUT31), .B(n694), .ZN(n730) );
  INV_X1 U785 ( .A(KEYINPUT103), .ZN(n696) );
  NAND2_X1 U786 ( .A1(G2067), .A2(n700), .ZN(n695) );
  XNOR2_X1 U787 ( .A(n696), .B(n695), .ZN(n698) );
  NAND2_X1 U788 ( .A1(G1348), .A2(n733), .ZN(n697) );
  NAND2_X1 U789 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U790 ( .A1(n987), .A2(n699), .ZN(n711) );
  NAND2_X1 U791 ( .A1(n699), .A2(n987), .ZN(n705) );
  XOR2_X1 U792 ( .A(KEYINPUT26), .B(KEYINPUT101), .Z(n702) );
  XNOR2_X1 U793 ( .A(G1996), .B(KEYINPUT100), .ZN(n946) );
  NAND2_X1 U794 ( .A1(n700), .A2(n946), .ZN(n701) );
  XNOR2_X1 U795 ( .A(n702), .B(n701), .ZN(n703) );
  XNOR2_X1 U796 ( .A(n703), .B(KEYINPUT64), .ZN(n704) );
  NAND2_X1 U797 ( .A1(n705), .A2(n704), .ZN(n709) );
  NAND2_X1 U798 ( .A1(n733), .A2(G1341), .ZN(n706) );
  XNOR2_X1 U799 ( .A(n706), .B(KEYINPUT102), .ZN(n707) );
  NAND2_X1 U800 ( .A1(n988), .A2(n707), .ZN(n708) );
  NOR2_X1 U801 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U802 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U803 ( .A(n712), .B(KEYINPUT104), .ZN(n717) );
  NAND2_X1 U804 ( .A1(n700), .A2(G2072), .ZN(n713) );
  XNOR2_X1 U805 ( .A(n713), .B(KEYINPUT27), .ZN(n715) );
  XNOR2_X1 U806 ( .A(G1956), .B(KEYINPUT99), .ZN(n916) );
  NOR2_X1 U807 ( .A1(n916), .A2(n700), .ZN(n714) );
  NOR2_X1 U808 ( .A1(n715), .A2(n714), .ZN(n718) );
  NAND2_X1 U809 ( .A1(n718), .A2(n984), .ZN(n716) );
  NAND2_X1 U810 ( .A1(n717), .A2(n716), .ZN(n721) );
  NOR2_X1 U811 ( .A1(n718), .A2(n984), .ZN(n719) );
  XOR2_X1 U812 ( .A(n719), .B(KEYINPUT28), .Z(n720) );
  NAND2_X1 U813 ( .A1(n721), .A2(n720), .ZN(n723) );
  XOR2_X1 U814 ( .A(KEYINPUT29), .B(KEYINPUT105), .Z(n722) );
  XNOR2_X1 U815 ( .A(n723), .B(n722), .ZN(n727) );
  AND2_X1 U816 ( .A1(n724), .A2(G171), .ZN(n725) );
  XNOR2_X1 U817 ( .A(n725), .B(KEYINPUT98), .ZN(n726) );
  NOR2_X1 U818 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U819 ( .A(KEYINPUT106), .B(n728), .ZN(n729) );
  NOR2_X1 U820 ( .A1(n730), .A2(n729), .ZN(n732) );
  NAND2_X1 U821 ( .A1(n742), .A2(G286), .ZN(n740) );
  INV_X1 U822 ( .A(G8), .ZN(n738) );
  NOR2_X1 U823 ( .A1(G1971), .A2(n773), .ZN(n735) );
  NOR2_X1 U824 ( .A1(G2090), .A2(n733), .ZN(n734) );
  NOR2_X1 U825 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U826 ( .A1(n736), .A2(G303), .ZN(n737) );
  OR2_X1 U827 ( .A1(n738), .A2(n737), .ZN(n739) );
  AND2_X1 U828 ( .A1(n740), .A2(n739), .ZN(n741) );
  INV_X1 U829 ( .A(n742), .ZN(n744) );
  NOR2_X1 U830 ( .A1(n744), .A2(n743), .ZN(n747) );
  NAND2_X1 U831 ( .A1(G8), .A2(n745), .ZN(n746) );
  NAND2_X1 U832 ( .A1(n747), .A2(n746), .ZN(n766) );
  NAND2_X1 U833 ( .A1(G1976), .A2(G288), .ZN(n993) );
  INV_X1 U834 ( .A(n773), .ZN(n748) );
  NAND2_X1 U835 ( .A1(n993), .A2(n748), .ZN(n757) );
  INV_X1 U836 ( .A(n757), .ZN(n752) );
  NOR2_X1 U837 ( .A1(G1976), .A2(G288), .ZN(n756) );
  NAND2_X1 U838 ( .A1(KEYINPUT33), .A2(n756), .ZN(n749) );
  NOR2_X1 U839 ( .A1(n773), .A2(n749), .ZN(n750) );
  XOR2_X1 U840 ( .A(KEYINPUT109), .B(n750), .Z(n760) );
  INV_X1 U841 ( .A(n760), .ZN(n751) );
  AND2_X1 U842 ( .A1(n752), .A2(n751), .ZN(n753) );
  AND2_X1 U843 ( .A1(n766), .A2(n753), .ZN(n754) );
  NAND2_X1 U844 ( .A1(n765), .A2(n754), .ZN(n762) );
  NOR2_X1 U845 ( .A1(G1971), .A2(G303), .ZN(n755) );
  NOR2_X1 U846 ( .A1(n756), .A2(n755), .ZN(n1004) );
  NOR2_X1 U847 ( .A1(n757), .A2(n1004), .ZN(n758) );
  NOR2_X1 U848 ( .A1(n758), .A2(KEYINPUT33), .ZN(n759) );
  OR2_X1 U849 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U850 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U851 ( .A(n763), .B(KEYINPUT110), .ZN(n764) );
  XOR2_X1 U852 ( .A(G1981), .B(G305), .Z(n995) );
  AND2_X1 U853 ( .A1(n764), .A2(n995), .ZN(n779) );
  NAND2_X1 U854 ( .A1(n766), .A2(n765), .ZN(n769) );
  NOR2_X1 U855 ( .A1(G2090), .A2(G303), .ZN(n767) );
  NAND2_X1 U856 ( .A1(G8), .A2(n767), .ZN(n768) );
  NAND2_X1 U857 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U858 ( .A1(n773), .A2(n770), .ZN(n777) );
  NOR2_X1 U859 ( .A1(G1981), .A2(G305), .ZN(n771) );
  XNOR2_X1 U860 ( .A(n771), .B(KEYINPUT24), .ZN(n772) );
  XNOR2_X1 U861 ( .A(n772), .B(KEYINPUT95), .ZN(n774) );
  NOR2_X1 U862 ( .A1(n774), .A2(n773), .ZN(n775) );
  XOR2_X1 U863 ( .A(n775), .B(KEYINPUT96), .Z(n776) );
  NAND2_X1 U864 ( .A1(n777), .A2(n776), .ZN(n778) );
  NOR2_X1 U865 ( .A1(n779), .A2(n778), .ZN(n812) );
  NOR2_X1 U866 ( .A1(n781), .A2(n780), .ZN(n826) );
  XNOR2_X1 U867 ( .A(KEYINPUT91), .B(KEYINPUT35), .ZN(n785) );
  NAND2_X1 U868 ( .A1(G116), .A2(n890), .ZN(n783) );
  NAND2_X1 U869 ( .A1(G128), .A2(n891), .ZN(n782) );
  NAND2_X1 U870 ( .A1(n783), .A2(n782), .ZN(n784) );
  XNOR2_X1 U871 ( .A(n785), .B(n784), .ZN(n791) );
  NAND2_X1 U872 ( .A1(n894), .A2(G104), .ZN(n786) );
  XNOR2_X1 U873 ( .A(n786), .B(KEYINPUT90), .ZN(n788) );
  NAND2_X1 U874 ( .A1(G140), .A2(n512), .ZN(n787) );
  NAND2_X1 U875 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U876 ( .A(KEYINPUT34), .B(n789), .ZN(n790) );
  NOR2_X1 U877 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U878 ( .A(KEYINPUT36), .B(n792), .ZN(n887) );
  XNOR2_X1 U879 ( .A(G2067), .B(KEYINPUT37), .ZN(n824) );
  NOR2_X1 U880 ( .A1(n887), .A2(n824), .ZN(n979) );
  NAND2_X1 U881 ( .A1(n826), .A2(n979), .ZN(n822) );
  NAND2_X1 U882 ( .A1(G95), .A2(n894), .ZN(n794) );
  NAND2_X1 U883 ( .A1(G131), .A2(n512), .ZN(n793) );
  NAND2_X1 U884 ( .A1(n794), .A2(n793), .ZN(n797) );
  NAND2_X1 U885 ( .A1(n890), .A2(G107), .ZN(n795) );
  XOR2_X1 U886 ( .A(KEYINPUT92), .B(n795), .Z(n796) );
  NOR2_X1 U887 ( .A1(n797), .A2(n796), .ZN(n799) );
  NAND2_X1 U888 ( .A1(n891), .A2(G119), .ZN(n798) );
  NAND2_X1 U889 ( .A1(n799), .A2(n798), .ZN(n873) );
  NAND2_X1 U890 ( .A1(n873), .A2(G1991), .ZN(n810) );
  NAND2_X1 U891 ( .A1(G117), .A2(n890), .ZN(n801) );
  NAND2_X1 U892 ( .A1(G141), .A2(n512), .ZN(n800) );
  NAND2_X1 U893 ( .A1(n801), .A2(n800), .ZN(n806) );
  XOR2_X1 U894 ( .A(KEYINPUT38), .B(KEYINPUT94), .Z(n803) );
  NAND2_X1 U895 ( .A1(G105), .A2(n894), .ZN(n802) );
  XNOR2_X1 U896 ( .A(n803), .B(n802), .ZN(n804) );
  XOR2_X1 U897 ( .A(KEYINPUT93), .B(n804), .Z(n805) );
  NOR2_X1 U898 ( .A1(n806), .A2(n805), .ZN(n808) );
  NAND2_X1 U899 ( .A1(n891), .A2(G129), .ZN(n807) );
  NAND2_X1 U900 ( .A1(n808), .A2(n807), .ZN(n901) );
  NAND2_X1 U901 ( .A1(G1996), .A2(n901), .ZN(n809) );
  NAND2_X1 U902 ( .A1(n810), .A2(n809), .ZN(n971) );
  NAND2_X1 U903 ( .A1(n971), .A2(n826), .ZN(n815) );
  NAND2_X1 U904 ( .A1(n822), .A2(n815), .ZN(n811) );
  NOR2_X1 U905 ( .A1(n812), .A2(n811), .ZN(n814) );
  XNOR2_X1 U906 ( .A(G1986), .B(G290), .ZN(n999) );
  NAND2_X1 U907 ( .A1(n999), .A2(n826), .ZN(n813) );
  NAND2_X1 U908 ( .A1(n814), .A2(n813), .ZN(n829) );
  NOR2_X1 U909 ( .A1(G1996), .A2(n901), .ZN(n965) );
  INV_X1 U910 ( .A(n815), .ZN(n818) );
  NOR2_X1 U911 ( .A1(G1986), .A2(G290), .ZN(n816) );
  NOR2_X1 U912 ( .A1(G1991), .A2(n873), .ZN(n968) );
  NOR2_X1 U913 ( .A1(n816), .A2(n968), .ZN(n817) );
  NOR2_X1 U914 ( .A1(n818), .A2(n817), .ZN(n819) );
  XOR2_X1 U915 ( .A(KEYINPUT111), .B(n819), .Z(n820) );
  NOR2_X1 U916 ( .A1(n965), .A2(n820), .ZN(n821) );
  XNOR2_X1 U917 ( .A(n821), .B(KEYINPUT39), .ZN(n823) );
  NAND2_X1 U918 ( .A1(n823), .A2(n822), .ZN(n825) );
  NAND2_X1 U919 ( .A1(n887), .A2(n824), .ZN(n980) );
  NAND2_X1 U920 ( .A1(n825), .A2(n980), .ZN(n827) );
  NAND2_X1 U921 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U922 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U923 ( .A(KEYINPUT40), .B(n830), .ZN(G329) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n831), .ZN(G217) );
  AND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n832) );
  NAND2_X1 U926 ( .A1(G661), .A2(n832), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n833) );
  NAND2_X1 U928 ( .A1(n834), .A2(n833), .ZN(G188) );
  XOR2_X1 U929 ( .A(G96), .B(KEYINPUT112), .Z(G221) );
  INV_X1 U931 ( .A(G132), .ZN(G219) );
  INV_X1 U932 ( .A(G120), .ZN(G236) );
  INV_X1 U933 ( .A(G82), .ZN(G220) );
  INV_X1 U934 ( .A(G69), .ZN(G235) );
  NOR2_X1 U935 ( .A1(n836), .A2(n835), .ZN(G325) );
  INV_X1 U936 ( .A(G325), .ZN(G261) );
  XOR2_X1 U937 ( .A(KEYINPUT121), .B(n837), .Z(n840) );
  XNOR2_X1 U938 ( .A(n838), .B(n988), .ZN(n839) );
  XNOR2_X1 U939 ( .A(n840), .B(n839), .ZN(n842) );
  XNOR2_X1 U940 ( .A(G286), .B(G171), .ZN(n841) );
  XNOR2_X1 U941 ( .A(n842), .B(n841), .ZN(n843) );
  NOR2_X1 U942 ( .A1(G37), .A2(n843), .ZN(G397) );
  XNOR2_X1 U943 ( .A(G1991), .B(G2474), .ZN(n853) );
  XOR2_X1 U944 ( .A(G1956), .B(G1961), .Z(n845) );
  XNOR2_X1 U945 ( .A(G1996), .B(G1976), .ZN(n844) );
  XNOR2_X1 U946 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U947 ( .A(G1966), .B(G1971), .Z(n847) );
  XNOR2_X1 U948 ( .A(G1986), .B(G1981), .ZN(n846) );
  XNOR2_X1 U949 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U950 ( .A(n849), .B(n848), .Z(n851) );
  XNOR2_X1 U951 ( .A(KEYINPUT116), .B(KEYINPUT41), .ZN(n850) );
  XNOR2_X1 U952 ( .A(n851), .B(n850), .ZN(n852) );
  XNOR2_X1 U953 ( .A(n853), .B(n852), .ZN(G229) );
  XNOR2_X1 U954 ( .A(G2067), .B(G2078), .ZN(n854) );
  XNOR2_X1 U955 ( .A(n854), .B(KEYINPUT42), .ZN(n864) );
  XOR2_X1 U956 ( .A(KEYINPUT114), .B(KEYINPUT113), .Z(n856) );
  XNOR2_X1 U957 ( .A(KEYINPUT115), .B(G2096), .ZN(n855) );
  XNOR2_X1 U958 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U959 ( .A(G2100), .B(G2090), .Z(n858) );
  XNOR2_X1 U960 ( .A(G2084), .B(G2072), .ZN(n857) );
  XNOR2_X1 U961 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U962 ( .A(n860), .B(n859), .Z(n862) );
  XNOR2_X1 U963 ( .A(G2678), .B(KEYINPUT43), .ZN(n861) );
  XNOR2_X1 U964 ( .A(n862), .B(n861), .ZN(n863) );
  XNOR2_X1 U965 ( .A(n864), .B(n863), .ZN(G227) );
  NAND2_X1 U966 ( .A1(G124), .A2(n891), .ZN(n865) );
  XOR2_X1 U967 ( .A(KEYINPUT117), .B(n865), .Z(n866) );
  XNOR2_X1 U968 ( .A(n866), .B(KEYINPUT44), .ZN(n868) );
  NAND2_X1 U969 ( .A1(G112), .A2(n890), .ZN(n867) );
  NAND2_X1 U970 ( .A1(n868), .A2(n867), .ZN(n872) );
  NAND2_X1 U971 ( .A1(G100), .A2(n894), .ZN(n870) );
  NAND2_X1 U972 ( .A1(G136), .A2(n512), .ZN(n869) );
  NAND2_X1 U973 ( .A1(n870), .A2(n869), .ZN(n871) );
  NOR2_X1 U974 ( .A1(n872), .A2(n871), .ZN(G162) );
  XNOR2_X1 U975 ( .A(KEYINPUT46), .B(KEYINPUT119), .ZN(n875) );
  XNOR2_X1 U976 ( .A(n873), .B(KEYINPUT48), .ZN(n874) );
  XNOR2_X1 U977 ( .A(n875), .B(n874), .ZN(n886) );
  NAND2_X1 U978 ( .A1(G103), .A2(n894), .ZN(n877) );
  NAND2_X1 U979 ( .A1(G139), .A2(n512), .ZN(n876) );
  NAND2_X1 U980 ( .A1(n877), .A2(n876), .ZN(n882) );
  NAND2_X1 U981 ( .A1(G115), .A2(n890), .ZN(n879) );
  NAND2_X1 U982 ( .A1(G127), .A2(n891), .ZN(n878) );
  NAND2_X1 U983 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U984 ( .A(KEYINPUT47), .B(n880), .Z(n881) );
  NOR2_X1 U985 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U986 ( .A(KEYINPUT118), .B(n883), .Z(n960) );
  XNOR2_X1 U987 ( .A(G160), .B(n960), .ZN(n884) );
  XNOR2_X1 U988 ( .A(n884), .B(G162), .ZN(n885) );
  XNOR2_X1 U989 ( .A(n886), .B(n885), .ZN(n889) );
  XNOR2_X1 U990 ( .A(n887), .B(n967), .ZN(n888) );
  XNOR2_X1 U991 ( .A(n889), .B(n888), .ZN(n905) );
  NAND2_X1 U992 ( .A1(G118), .A2(n890), .ZN(n893) );
  NAND2_X1 U993 ( .A1(G130), .A2(n891), .ZN(n892) );
  NAND2_X1 U994 ( .A1(n893), .A2(n892), .ZN(n900) );
  NAND2_X1 U995 ( .A1(G106), .A2(n894), .ZN(n897) );
  NAND2_X1 U996 ( .A1(G142), .A2(n512), .ZN(n896) );
  NAND2_X1 U997 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U998 ( .A(n898), .B(KEYINPUT45), .Z(n899) );
  NOR2_X1 U999 ( .A1(n900), .A2(n899), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(n902), .B(n901), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(G164), .B(n903), .ZN(n904) );
  XNOR2_X1 U1002 ( .A(n905), .B(n904), .ZN(n906) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n906), .ZN(n907) );
  XNOR2_X1 U1004 ( .A(KEYINPUT120), .B(n907), .ZN(G395) );
  NOR2_X1 U1005 ( .A1(G229), .A2(G227), .ZN(n908) );
  XNOR2_X1 U1006 ( .A(KEYINPUT49), .B(n908), .ZN(n909) );
  NOR2_X1 U1007 ( .A1(G397), .A2(n909), .ZN(n913) );
  NOR2_X1 U1008 ( .A1(n914), .A2(G401), .ZN(n910) );
  XOR2_X1 U1009 ( .A(KEYINPUT122), .B(n910), .Z(n911) );
  NOR2_X1 U1010 ( .A1(G395), .A2(n911), .ZN(n912) );
  NAND2_X1 U1011 ( .A1(n913), .A2(n912), .ZN(G225) );
  INV_X1 U1012 ( .A(G225), .ZN(G308) );
  INV_X1 U1013 ( .A(n914), .ZN(G319) );
  INV_X1 U1014 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1015 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n1016) );
  XNOR2_X1 U1016 ( .A(G5), .B(n915), .ZN(n928) );
  XNOR2_X1 U1017 ( .A(G20), .B(n916), .ZN(n920) );
  XNOR2_X1 U1018 ( .A(G1981), .B(G6), .ZN(n918) );
  XNOR2_X1 U1019 ( .A(G1341), .B(G19), .ZN(n917) );
  NOR2_X1 U1020 ( .A1(n918), .A2(n917), .ZN(n919) );
  NAND2_X1 U1021 ( .A1(n920), .A2(n919), .ZN(n923) );
  XOR2_X1 U1022 ( .A(KEYINPUT59), .B(G1348), .Z(n921) );
  XNOR2_X1 U1023 ( .A(G4), .B(n921), .ZN(n922) );
  NOR2_X1 U1024 ( .A1(n923), .A2(n922), .ZN(n924) );
  XOR2_X1 U1025 ( .A(KEYINPUT60), .B(n924), .Z(n926) );
  XNOR2_X1 U1026 ( .A(G1966), .B(G21), .ZN(n925) );
  NOR2_X1 U1027 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1028 ( .A1(n928), .A2(n927), .ZN(n936) );
  XNOR2_X1 U1029 ( .A(G1986), .B(G24), .ZN(n930) );
  XNOR2_X1 U1030 ( .A(G23), .B(G1976), .ZN(n929) );
  NOR2_X1 U1031 ( .A1(n930), .A2(n929), .ZN(n933) );
  XOR2_X1 U1032 ( .A(G1971), .B(KEYINPUT124), .Z(n931) );
  XNOR2_X1 U1033 ( .A(G22), .B(n931), .ZN(n932) );
  NAND2_X1 U1034 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1035 ( .A(KEYINPUT58), .B(n934), .ZN(n935) );
  NOR2_X1 U1036 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1037 ( .A(KEYINPUT61), .B(n937), .Z(n938) );
  NOR2_X1 U1038 ( .A1(G16), .A2(n938), .ZN(n939) );
  XOR2_X1 U1039 ( .A(KEYINPUT125), .B(n939), .Z(n1014) );
  XOR2_X1 U1040 ( .A(G2090), .B(G35), .Z(n942) );
  XOR2_X1 U1041 ( .A(KEYINPUT54), .B(G34), .Z(n940) );
  XNOR2_X1 U1042 ( .A(G2084), .B(n940), .ZN(n941) );
  NAND2_X1 U1043 ( .A1(n942), .A2(n941), .ZN(n956) );
  XNOR2_X1 U1044 ( .A(G1991), .B(G25), .ZN(n944) );
  XNOR2_X1 U1045 ( .A(G33), .B(G2072), .ZN(n943) );
  NOR2_X1 U1046 ( .A1(n944), .A2(n943), .ZN(n950) );
  XOR2_X1 U1047 ( .A(G2067), .B(G26), .Z(n945) );
  NAND2_X1 U1048 ( .A1(n945), .A2(G28), .ZN(n948) );
  XNOR2_X1 U1049 ( .A(G32), .B(n946), .ZN(n947) );
  NOR2_X1 U1050 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1051 ( .A1(n950), .A2(n949), .ZN(n953) );
  XOR2_X1 U1052 ( .A(G27), .B(n951), .Z(n952) );
  NOR2_X1 U1053 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1054 ( .A(n954), .B(KEYINPUT53), .ZN(n955) );
  NOR2_X1 U1055 ( .A1(n956), .A2(n955), .ZN(n957) );
  XOR2_X1 U1056 ( .A(KEYINPUT123), .B(n957), .Z(n958) );
  NOR2_X1 U1057 ( .A1(G29), .A2(n958), .ZN(n959) );
  XOR2_X1 U1058 ( .A(KEYINPUT55), .B(n959), .Z(n1011) );
  XOR2_X1 U1059 ( .A(G164), .B(G2078), .Z(n962) );
  XNOR2_X1 U1060 ( .A(G2072), .B(n960), .ZN(n961) );
  NOR2_X1 U1061 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1062 ( .A(KEYINPUT50), .B(n963), .ZN(n977) );
  XOR2_X1 U1063 ( .A(G2090), .B(G162), .Z(n964) );
  NOR2_X1 U1064 ( .A1(n965), .A2(n964), .ZN(n966) );
  XOR2_X1 U1065 ( .A(KEYINPUT51), .B(n966), .Z(n970) );
  NOR2_X1 U1066 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1067 ( .A1(n970), .A2(n969), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(G160), .B(G2084), .ZN(n973) );
  INV_X1 U1069 ( .A(n971), .ZN(n972) );
  NAND2_X1 U1070 ( .A1(n973), .A2(n972), .ZN(n974) );
  NOR2_X1 U1071 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n978) );
  NOR2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n981) );
  NAND2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1075 ( .A(n982), .B(KEYINPUT52), .ZN(n983) );
  NAND2_X1 U1076 ( .A1(n983), .A2(G29), .ZN(n1009) );
  XNOR2_X1 U1077 ( .A(KEYINPUT56), .B(G16), .ZN(n1007) );
  XNOR2_X1 U1078 ( .A(G1956), .B(n984), .ZN(n986) );
  NAND2_X1 U1079 ( .A1(G1971), .A2(G303), .ZN(n985) );
  NAND2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n992) );
  XOR2_X1 U1081 ( .A(n987), .B(G1348), .Z(n990) );
  XNOR2_X1 U1082 ( .A(n988), .B(G1341), .ZN(n989) );
  NAND2_X1 U1083 ( .A1(n990), .A2(n989), .ZN(n991) );
  NOR2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n994) );
  NAND2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n1003) );
  XNOR2_X1 U1086 ( .A(G1966), .B(G168), .ZN(n996) );
  NAND2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1088 ( .A(n997), .B(KEYINPUT57), .ZN(n1001) );
  XNOR2_X1 U1089 ( .A(G1961), .B(G301), .ZN(n998) );
  NOR2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NOR2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1005) );
  NAND2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1094 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1095 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NOR2_X1 U1096 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1097 ( .A1(n1012), .A2(G11), .ZN(n1013) );
  NOR2_X1 U1098 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1099 ( .A(n1016), .B(n1015), .ZN(G311) );
  XNOR2_X1 U1100 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
endmodule

