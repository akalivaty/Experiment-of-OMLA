//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 1 1 0 1 1 0 1 1 1 0 1 0 1 0 0 0 1 0 1 1 1 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:12 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n569, new_n570, new_n571, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n626, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT65), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  XNOR2_X1  g030(.A(G325), .B(KEYINPUT66), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT67), .Z(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT68), .Z(G319));
  INV_X1    g034(.A(KEYINPUT69), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  OAI21_X1  g036(.A(new_n460), .B1(new_n461), .B2(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n464), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n462), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G137), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n464), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(new_n463), .ZN(new_n471));
  INV_X1    g046(.A(G125), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2104), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT70), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n476), .B(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G101), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n468), .A2(new_n474), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  NAND4_X1  g056(.A1(new_n462), .A2(new_n465), .A3(G2105), .A4(new_n463), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  AND2_X1   g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(G112), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n485), .B1(new_n486), .B2(G2105), .ZN(new_n487));
  OR3_X1    g062(.A1(new_n466), .A2(KEYINPUT71), .A3(G2105), .ZN(new_n488));
  OAI21_X1  g063(.A(KEYINPUT71), .B1(new_n466), .B2(G2105), .ZN(new_n489));
  AND2_X1   g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AOI211_X1 g065(.A(new_n484), .B(new_n487), .C1(new_n490), .C2(G136), .ZN(G162));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n462), .A2(new_n465), .A3(new_n493), .A4(new_n463), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n470), .A2(new_n463), .ZN(new_n495));
  NOR3_X1   g070(.A1(new_n492), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n496));
  AOI22_X1  g071(.A1(new_n494), .A2(KEYINPUT4), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OR2_X1    g072(.A1(G102), .A2(G2105), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n498), .B(G2104), .C1(G114), .C2(new_n475), .ZN(new_n499));
  INV_X1    g074(.A(G126), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n499), .B1(new_n482), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n497), .A2(new_n501), .ZN(G164));
  INV_X1    g077(.A(KEYINPUT72), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT6), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n503), .B1(new_n504), .B2(G651), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(KEYINPUT72), .A3(KEYINPUT6), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT73), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n509), .B1(new_n506), .B2(KEYINPUT6), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n504), .A2(KEYINPUT73), .A3(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OR2_X1    g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n508), .A2(new_n512), .A3(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT74), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g093(.A1(new_n508), .A2(new_n512), .A3(KEYINPUT74), .A4(new_n515), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G88), .ZN(new_n521));
  AND3_X1   g096(.A1(new_n508), .A2(new_n512), .A3(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(G75), .A2(G543), .ZN(new_n523));
  XOR2_X1   g098(.A(KEYINPUT5), .B(G543), .Z(new_n524));
  INV_X1    g099(.A(G62), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n522), .A2(G50), .B1(new_n526), .B2(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n521), .A2(new_n527), .ZN(G303));
  INV_X1    g103(.A(G303), .ZN(G166));
  NAND3_X1  g104(.A1(new_n518), .A2(G89), .A3(new_n519), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT75), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n530), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  AND2_X1   g109(.A1(G63), .A2(G651), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n522), .A2(G51), .B1(new_n515), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n531), .B1(new_n530), .B2(new_n533), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n537), .A2(new_n538), .ZN(G168));
  NAND2_X1  g114(.A1(new_n518), .A2(new_n519), .ZN(new_n540));
  INV_X1    g115(.A(G90), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT76), .ZN(new_n543));
  NAND2_X1  g118(.A1(G77), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G64), .ZN(new_n545));
  OAI211_X1 g120(.A(new_n543), .B(new_n544), .C1(new_n524), .C2(new_n545), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n545), .B1(new_n513), .B2(new_n514), .ZN(new_n547));
  INV_X1    g122(.A(new_n544), .ZN(new_n548));
  OAI21_X1  g123(.A(KEYINPUT76), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n546), .A2(new_n549), .A3(G651), .ZN(new_n550));
  INV_X1    g125(.A(new_n522), .ZN(new_n551));
  INV_X1    g126(.A(G52), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n542), .A2(new_n553), .ZN(G171));
  NAND2_X1  g129(.A1(G68), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G56), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n524), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n557), .A2(KEYINPUT77), .A3(G651), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT77), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n560), .B2(new_n506), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n522), .A2(G43), .ZN(new_n563));
  INV_X1    g138(.A(G81), .ZN(new_n564));
  OAI211_X1 g139(.A(new_n562), .B(new_n563), .C1(new_n564), .C2(new_n540), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g143(.A(KEYINPUT78), .B(KEYINPUT8), .Z(new_n569));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n569), .B(new_n570), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(G188));
  NAND4_X1  g147(.A1(new_n508), .A2(new_n512), .A3(G53), .A4(G543), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT79), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(KEYINPUT9), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n573), .B(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(G78), .A2(G543), .ZN(new_n578));
  XNOR2_X1  g153(.A(KEYINPUT80), .B(G65), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n524), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(G651), .ZN(new_n581));
  INV_X1    g156(.A(G91), .ZN(new_n582));
  OAI211_X1 g157(.A(new_n577), .B(new_n581), .C1(new_n582), .C2(new_n540), .ZN(G299));
  OAI221_X1 g158(.A(new_n550), .B1(new_n551), .B2(new_n552), .C1(new_n540), .C2(new_n541), .ZN(G301));
  INV_X1    g159(.A(G168), .ZN(G286));
  NAND2_X1  g160(.A1(new_n520), .A2(G87), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n515), .A2(G74), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n522), .A2(G49), .B1(new_n587), .B2(G651), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n586), .A2(new_n588), .ZN(G288));
  NAND2_X1  g164(.A1(new_n520), .A2(G86), .ZN(new_n590));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G61), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n524), .B2(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n522), .A2(G48), .B1(new_n593), .B2(G651), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n590), .A2(new_n594), .ZN(G305));
  NAND2_X1  g170(.A1(new_n520), .A2(G85), .ZN(new_n596));
  NAND2_X1  g171(.A1(G72), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G60), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n524), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n522), .A2(G47), .B1(new_n599), .B2(G651), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n596), .A2(new_n600), .ZN(G290));
  NAND2_X1  g176(.A1(G301), .A2(G868), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n518), .A2(G92), .A3(new_n519), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(KEYINPUT81), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT81), .ZN(new_n605));
  NAND4_X1  g180(.A1(new_n518), .A2(new_n605), .A3(G92), .A4(new_n519), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT10), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n604), .A2(KEYINPUT10), .A3(new_n606), .ZN(new_n610));
  NAND2_X1  g185(.A1(G79), .A2(G543), .ZN(new_n611));
  INV_X1    g186(.A(G66), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n524), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(G651), .ZN(new_n614));
  INV_X1    g189(.A(G54), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n551), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(KEYINPUT82), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT82), .ZN(new_n618));
  OAI211_X1 g193(.A(new_n618), .B(new_n614), .C1(new_n551), .C2(new_n615), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  AND3_X1   g195(.A1(new_n609), .A2(new_n610), .A3(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n602), .B1(new_n621), .B2(G868), .ZN(G284));
  OAI21_X1  g197(.A(new_n602), .B1(new_n621), .B2(G868), .ZN(G321));
  MUX2_X1   g198(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g199(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g200(.A(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n621), .B1(new_n626), .B2(G860), .ZN(G148));
  NAND2_X1  g202(.A1(new_n621), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G868), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(G868), .B2(new_n566), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g206(.A1(new_n478), .A2(new_n495), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT12), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT13), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2100), .ZN(new_n635));
  INV_X1    g210(.A(G123), .ZN(new_n636));
  OAI21_X1  g211(.A(KEYINPUT83), .B1(new_n475), .B2(G111), .ZN(new_n637));
  OR2_X1    g212(.A1(G99), .A2(G2105), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n637), .A2(G2104), .A3(new_n638), .ZN(new_n639));
  NOR3_X1   g214(.A1(new_n475), .A2(KEYINPUT83), .A3(G111), .ZN(new_n640));
  OAI22_X1  g215(.A1(new_n482), .A2(new_n636), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(new_n490), .ZN(new_n643));
  INV_X1    g218(.A(G135), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n642), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n645), .A2(G2096), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(G2096), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n635), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT84), .Z(G156));
  XNOR2_X1  g224(.A(G2427), .B(G2438), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2430), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT15), .B(G2435), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n652), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(KEYINPUT14), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G1341), .B(G1348), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2451), .B(G2454), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT16), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT85), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n659), .A2(new_n663), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n664), .A2(G14), .A3(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(G401));
  INV_X1    g242(.A(KEYINPUT18), .ZN(new_n668));
  XOR2_X1   g243(.A(G2084), .B(G2090), .Z(new_n669));
  XNOR2_X1  g244(.A(G2067), .B(G2678), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(KEYINPUT17), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n669), .A2(new_n670), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n668), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(G2100), .ZN(new_n675));
  XOR2_X1   g250(.A(G2072), .B(G2078), .Z(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(new_n671), .B2(KEYINPUT18), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G2096), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n675), .B(new_n678), .ZN(G227));
  XNOR2_X1  g254(.A(G1961), .B(G1966), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT86), .ZN(new_n681));
  XOR2_X1   g256(.A(G1956), .B(G2474), .Z(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1971), .B(G1976), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT19), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n686), .B(KEYINPUT20), .Z(new_n687));
  OR2_X1    g262(.A1(new_n681), .A2(new_n682), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(new_n683), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n689), .A2(KEYINPUT87), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(KEYINPUT87), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(new_n685), .ZN(new_n692));
  OAI221_X1 g267(.A(new_n687), .B1(new_n688), .B2(new_n685), .C1(new_n690), .C2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT88), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1991), .B(G1996), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n698));
  XOR2_X1   g273(.A(new_n697), .B(new_n698), .Z(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n694), .A2(new_n700), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n693), .A2(KEYINPUT88), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n693), .A2(KEYINPUT88), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n702), .A2(new_n703), .A3(new_n699), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n701), .A2(new_n704), .ZN(G229));
  INV_X1    g280(.A(G16), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G22), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G166), .B2(new_n706), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(G1971), .Z(new_n709));
  NOR2_X1   g284(.A1(G16), .A2(G23), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT90), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G288), .B2(new_n706), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT33), .B(G1976), .Z(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(G6), .A2(G16), .ZN(new_n715));
  INV_X1    g290(.A(G305), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n715), .B1(new_n716), .B2(G16), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT32), .B(G1981), .Z(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n709), .A2(new_n714), .A3(new_n719), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n720), .A2(KEYINPUT34), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(KEYINPUT34), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n706), .A2(G24), .ZN(new_n723));
  INV_X1    g298(.A(G290), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(new_n724), .B2(new_n706), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G1986), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n726), .A2(KEYINPUT89), .ZN(new_n727));
  INV_X1    g302(.A(G29), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G25), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n490), .A2(G131), .ZN(new_n730));
  OAI21_X1  g305(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n731));
  INV_X1    g306(.A(G107), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n731), .B1(new_n732), .B2(G2105), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n483), .B2(G119), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n730), .A2(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n729), .B1(new_n736), .B2(new_n728), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT35), .B(G1991), .Z(new_n738));
  XOR2_X1   g313(.A(new_n737), .B(new_n738), .Z(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(KEYINPUT89), .B2(new_n726), .ZN(new_n740));
  NAND4_X1  g315(.A1(new_n721), .A2(new_n722), .A3(new_n727), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT36), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n728), .A2(G32), .ZN(new_n743));
  NAND3_X1  g318(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT26), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n478), .A2(G105), .ZN(new_n746));
  AOI211_X1 g321(.A(new_n745), .B(new_n746), .C1(G129), .C2(new_n483), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n490), .A2(G141), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n743), .B1(new_n750), .B2(new_n728), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT93), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT27), .B(G1996), .ZN(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n706), .A2(G20), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT23), .Z(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G299), .B2(G16), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G1956), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n755), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n752), .A2(new_n754), .ZN(new_n761));
  NOR2_X1   g336(.A1(G4), .A2(G16), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n621), .B2(G16), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT91), .B(G1348), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n763), .A2(new_n765), .ZN(new_n767));
  NOR4_X1   g342(.A1(new_n760), .A2(new_n761), .A3(new_n766), .A4(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n728), .A2(G35), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G162), .B2(new_n728), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT29), .Z(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G2090), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n728), .A2(G27), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G164), .B2(new_n728), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G2078), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n706), .A2(G19), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n566), .B2(new_n706), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G1341), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n728), .A2(G26), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT28), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n490), .A2(G140), .ZN(new_n781));
  OAI21_X1  g356(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n782));
  INV_X1    g357(.A(G116), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(G2105), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n483), .B2(G128), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n780), .B1(new_n787), .B2(new_n728), .ZN(new_n788));
  AOI211_X1 g363(.A(new_n775), .B(new_n778), .C1(G2067), .C2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n706), .A2(G5), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G171), .B2(new_n706), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G1961), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n788), .A2(G2067), .ZN(new_n793));
  INV_X1    g368(.A(G34), .ZN(new_n794));
  AOI21_X1  g369(.A(G29), .B1(new_n794), .B2(KEYINPUT24), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(KEYINPUT24), .B2(new_n794), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n480), .B2(new_n728), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G2084), .ZN(new_n798));
  INV_X1    g373(.A(G28), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n799), .A2(KEYINPUT30), .ZN(new_n800));
  AOI21_X1  g375(.A(G29), .B1(new_n799), .B2(KEYINPUT30), .ZN(new_n801));
  OR2_X1    g376(.A1(KEYINPUT31), .A2(G11), .ZN(new_n802));
  NAND2_X1  g377(.A1(KEYINPUT31), .A2(G11), .ZN(new_n803));
  AOI22_X1  g378(.A1(new_n800), .A2(new_n801), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  OAI211_X1 g379(.A(new_n798), .B(new_n804), .C1(new_n728), .C2(new_n645), .ZN(new_n805));
  NOR3_X1   g380(.A1(new_n792), .A2(new_n793), .A3(new_n805), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n772), .A2(new_n789), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n706), .A2(G21), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G168), .B2(new_n706), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT94), .Z(new_n810));
  NOR2_X1   g385(.A1(new_n810), .A2(G1966), .ZN(new_n811));
  AND2_X1   g386(.A1(new_n810), .A2(G1966), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n490), .A2(G139), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT92), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(G115), .A2(G2104), .ZN(new_n816));
  INV_X1    g391(.A(G127), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n471), .B2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT25), .ZN(new_n819));
  NAND2_X1  g394(.A1(G103), .A2(G2104), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n819), .B1(new_n820), .B2(G2105), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n475), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n822));
  AOI22_X1  g397(.A1(new_n818), .A2(G2105), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n815), .A2(new_n823), .ZN(new_n824));
  MUX2_X1   g399(.A(G33), .B(new_n824), .S(G29), .Z(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G2072), .ZN(new_n826));
  NOR4_X1   g401(.A1(new_n807), .A2(new_n811), .A3(new_n812), .A4(new_n826), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n742), .A2(new_n768), .A3(new_n827), .ZN(G150));
  INV_X1    g403(.A(G150), .ZN(G311));
  NAND3_X1  g404(.A1(new_n518), .A2(G93), .A3(new_n519), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n508), .A2(new_n512), .A3(G55), .A4(G543), .ZN(new_n831));
  INV_X1    g406(.A(G67), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n832), .B1(new_n513), .B2(new_n514), .ZN(new_n833));
  AND2_X1   g408(.A1(G80), .A2(G543), .ZN(new_n834));
  OAI21_X1  g409(.A(G651), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AND2_X1   g410(.A1(new_n831), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n830), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(KEYINPUT95), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT95), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n830), .A2(new_n839), .A3(new_n836), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(G860), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT37), .Z(new_n843));
  NAND2_X1  g418(.A1(new_n621), .A2(G559), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT38), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT96), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n838), .A2(new_n565), .A3(new_n846), .A4(new_n840), .ZN(new_n847));
  AND3_X1   g422(.A1(new_n838), .A2(new_n565), .A3(new_n840), .ZN(new_n848));
  INV_X1    g423(.A(new_n837), .ZN(new_n849));
  OAI21_X1  g424(.A(KEYINPUT96), .B1(new_n565), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n847), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n845), .B(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT39), .ZN(new_n853));
  AOI21_X1  g428(.A(G860), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n854), .B1(new_n853), .B2(new_n852), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n855), .A2(KEYINPUT97), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n855), .A2(KEYINPUT97), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n843), .B1(new_n856), .B2(new_n857), .ZN(G145));
  NAND2_X1  g433(.A1(new_n490), .A2(G142), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT98), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  OR2_X1    g436(.A1(G106), .A2(G2105), .ZN(new_n862));
  OAI211_X1 g437(.A(new_n862), .B(G2104), .C1(G118), .C2(new_n475), .ZN(new_n863));
  INV_X1    g438(.A(G130), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n863), .B1(new_n482), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n861), .A2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(G164), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n786), .B(new_n867), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n866), .A2(new_n868), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n824), .A2(new_n749), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n815), .A2(new_n750), .A3(new_n823), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n735), .B(new_n633), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n872), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n875), .B1(new_n872), .B2(new_n873), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n871), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n872), .A2(new_n873), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(new_n874), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n881), .A2(new_n876), .A3(new_n869), .A4(new_n870), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n645), .B(G160), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(G162), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n879), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(G37), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n884), .B1(new_n879), .B2(new_n882), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  XOR2_X1   g464(.A(new_n889), .B(KEYINPUT40), .Z(G395));
  XOR2_X1   g465(.A(G303), .B(G288), .Z(new_n891));
  XOR2_X1   g466(.A(G305), .B(G290), .Z(new_n892));
  XOR2_X1   g467(.A(new_n891), .B(new_n892), .Z(new_n893));
  XOR2_X1   g468(.A(new_n893), .B(KEYINPUT42), .Z(new_n894));
  XOR2_X1   g469(.A(new_n628), .B(new_n851), .Z(new_n895));
  NAND4_X1  g470(.A1(new_n609), .A2(G299), .A3(new_n610), .A4(new_n620), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(KEYINPUT99), .ZN(new_n897));
  AOI22_X1  g472(.A1(new_n607), .A2(new_n608), .B1(new_n617), .B2(new_n619), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT99), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n898), .A2(new_n899), .A3(G299), .A4(new_n610), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT100), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n902), .B1(new_n621), .B2(G299), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n898), .A2(new_n610), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n520), .A2(G91), .ZN(new_n905));
  AND2_X1   g480(.A1(new_n577), .A2(new_n581), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n904), .A2(KEYINPUT100), .A3(new_n905), .A4(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n901), .A2(new_n903), .A3(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  OR2_X1    g484(.A1(new_n895), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT101), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n910), .B(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n908), .A2(KEYINPUT41), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT41), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n901), .A2(new_n903), .A3(new_n914), .A4(new_n907), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n895), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n894), .B1(new_n912), .B2(new_n916), .ZN(new_n917));
  OR2_X1    g492(.A1(new_n910), .A2(KEYINPUT101), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n910), .A2(KEYINPUT101), .ZN(new_n919));
  AND4_X1   g494(.A1(new_n916), .A2(new_n918), .A3(new_n919), .A4(new_n894), .ZN(new_n920));
  OAI21_X1  g495(.A(G868), .B1(new_n917), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n841), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n921), .B1(G868), .B2(new_n922), .ZN(G295));
  OAI21_X1  g498(.A(new_n921), .B1(G868), .B2(new_n922), .ZN(G331));
  XOR2_X1   g499(.A(KEYINPUT102), .B(KEYINPUT43), .Z(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(G301), .B1(new_n537), .B2(new_n538), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n530), .A2(new_n533), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(KEYINPUT75), .ZN(new_n929));
  NAND4_X1  g504(.A1(G171), .A2(new_n929), .A3(new_n534), .A4(new_n536), .ZN(new_n930));
  AND2_X1   g505(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n851), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n838), .A2(new_n565), .A3(new_n840), .ZN(new_n933));
  OAI211_X1 g508(.A(new_n933), .B(KEYINPUT96), .C1(new_n565), .C2(new_n849), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n927), .A2(new_n930), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n934), .A2(new_n935), .A3(new_n847), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n932), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n913), .A2(new_n915), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n908), .A2(new_n937), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT103), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n893), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n908), .A2(new_n937), .A3(KEYINPUT103), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n939), .A2(new_n942), .A3(new_n943), .A4(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n886), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n908), .A2(KEYINPUT103), .A3(new_n937), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT103), .B1(new_n908), .B2(new_n937), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n943), .B1(new_n949), .B2(new_n939), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n926), .B1(new_n946), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n943), .B1(new_n939), .B2(new_n940), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n954), .A2(new_n886), .A3(new_n945), .A4(new_n925), .ZN(new_n955));
  AND3_X1   g530(.A1(new_n951), .A2(new_n952), .A3(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n939), .A2(new_n942), .A3(new_n944), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(new_n893), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n958), .A2(new_n886), .A3(new_n945), .A4(new_n925), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT104), .ZN(new_n960));
  INV_X1    g535(.A(new_n946), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT104), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n961), .A2(new_n962), .A3(new_n958), .A4(new_n925), .ZN(new_n963));
  OAI21_X1  g538(.A(KEYINPUT43), .B1(new_n946), .B2(new_n953), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n960), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n956), .B1(new_n965), .B2(KEYINPUT44), .ZN(G397));
  NAND4_X1  g541(.A1(new_n468), .A2(new_n474), .A3(G40), .A4(new_n479), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(G1384), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n969), .B1(new_n497), .B2(new_n501), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT45), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OAI211_X1 g547(.A(KEYINPUT45), .B(new_n969), .C1(new_n497), .C2(new_n501), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n968), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT107), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n968), .A2(new_n972), .A3(KEYINPUT107), .A4(new_n973), .ZN(new_n977));
  XNOR2_X1  g552(.A(KEYINPUT108), .B(G1971), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT110), .ZN(new_n980));
  INV_X1    g555(.A(new_n970), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT50), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n980), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n970), .A2(KEYINPUT110), .A3(KEYINPUT50), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT109), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n986), .B1(new_n970), .B2(KEYINPUT50), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n987), .A2(new_n968), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n981), .A2(KEYINPUT109), .A3(new_n982), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n985), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n979), .B1(new_n990), .B2(G2090), .ZN(new_n991));
  NOR2_X1   g566(.A1(KEYINPUT111), .A2(KEYINPUT55), .ZN(new_n992));
  AND2_X1   g567(.A1(KEYINPUT111), .A2(KEYINPUT55), .ZN(new_n993));
  OAI211_X1 g568(.A(G303), .B(G8), .C1(new_n992), .C2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G8), .ZN(new_n995));
  NOR2_X1   g570(.A1(G166), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n994), .B1(new_n996), .B2(new_n993), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n991), .A2(G8), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT112), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n991), .A2(new_n997), .A3(KEYINPUT112), .A4(G8), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1981), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n716), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1003), .B1(new_n590), .B2(new_n594), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1004), .A2(KEYINPUT49), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT49), .ZN(new_n1008));
  NOR2_X1   g583(.A1(G305), .A2(G1981), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1008), .B1(new_n1009), .B2(new_n1005), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n995), .B1(new_n968), .B2(new_n981), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1007), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT114), .ZN(new_n1013));
  INV_X1    g588(.A(G1976), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n1011), .B(new_n1013), .C1(new_n1014), .C2(G288), .ZN(new_n1015));
  XOR2_X1   g590(.A(KEYINPUT113), .B(G1976), .Z(new_n1016));
  AOI21_X1  g591(.A(new_n1016), .B1(new_n586), .B2(new_n588), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT52), .B1(new_n1017), .B2(new_n1011), .ZN(new_n1018));
  AND2_X1   g593(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1012), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n967), .B1(KEYINPUT50), .B2(new_n970), .ZN(new_n1022));
  OR2_X1    g597(.A1(new_n1022), .A2(KEYINPUT116), .ZN(new_n1023));
  AOI22_X1  g598(.A1(new_n1022), .A2(KEYINPUT116), .B1(new_n982), .B2(new_n981), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n979), .B1(new_n1025), .B2(G2090), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n997), .B1(new_n1026), .B2(G8), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1021), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1002), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G1966), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n974), .A2(new_n1030), .ZN(new_n1031));
  OAI211_X1 g606(.A(G168), .B(new_n1031), .C1(new_n990), .C2(G2084), .ZN(new_n1032));
  OAI21_X1  g607(.A(G8), .B1(KEYINPUT123), .B2(KEYINPUT51), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(KEYINPUT123), .A2(KEYINPUT51), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1032), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1031), .B1(new_n990), .B2(G2084), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1037), .A2(G8), .A3(G286), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1035), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1029), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n1043));
  AOI21_X1  g618(.A(G2078), .B1(new_n976), .B2(new_n977), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT124), .ZN(new_n1045));
  OR3_X1    g620(.A1(new_n1044), .A2(new_n1045), .A3(KEYINPUT53), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1045), .B1(new_n1044), .B2(KEYINPUT53), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n1049));
  NOR3_X1   g624(.A1(new_n974), .A2(new_n1049), .A3(G2078), .ZN(new_n1050));
  INV_X1    g625(.A(G1961), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1050), .B1(new_n990), .B2(new_n1051), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n1048), .A2(G301), .A3(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(G301), .B1(new_n1048), .B2(new_n1052), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1043), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1048), .A2(new_n1052), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(G171), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1048), .A2(G301), .A3(new_n1052), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1057), .A2(KEYINPUT54), .A3(new_n1058), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n1042), .A2(new_n1055), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n968), .A2(new_n981), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1061), .A2(G2067), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1062), .B1(new_n990), .B2(new_n764), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  OR2_X1    g639(.A1(new_n904), .A2(KEYINPUT60), .ZN(new_n1065));
  XOR2_X1   g640(.A(KEYINPUT58), .B(G1341), .Z(new_n1066));
  NAND2_X1  g641(.A1(new_n1061), .A2(new_n1066), .ZN(new_n1067));
  XNOR2_X1  g642(.A(KEYINPUT121), .B(G1996), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1067), .B1(new_n974), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n1069), .A2(new_n566), .A3(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1070), .B1(new_n1069), .B2(new_n566), .ZN(new_n1072));
  OAI22_X1  g647(.A1(new_n1064), .A2(new_n1065), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  XNOR2_X1  g648(.A(new_n1063), .B(new_n904), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1073), .B1(new_n1074), .B2(KEYINPUT60), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT61), .ZN(new_n1076));
  AOI21_X1  g651(.A(G1956), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1077));
  XOR2_X1   g652(.A(KEYINPUT56), .B(G2072), .Z(new_n1078));
  NOR2_X1   g653(.A1(new_n974), .A2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT118), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT57), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n905), .A2(new_n1083), .A3(new_n581), .A4(new_n577), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n1081), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1082), .B1(new_n1081), .B2(new_n1084), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(KEYINPUT119), .B1(new_n1080), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT119), .ZN(new_n1089));
  OAI221_X1 g664(.A(new_n1089), .B1(new_n1085), .B2(new_n1086), .C1(new_n1077), .C2(new_n1079), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1081), .A2(new_n1084), .ZN(new_n1092));
  NOR3_X1   g667(.A1(new_n1077), .A2(new_n1092), .A3(new_n1079), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1076), .B1(new_n1091), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1080), .B1(new_n1081), .B2(new_n1084), .ZN(new_n1096));
  NOR3_X1   g671(.A1(new_n1096), .A2(new_n1093), .A3(KEYINPUT61), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1075), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT120), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT117), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1100), .B1(new_n1063), .B2(new_n904), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n989), .A2(new_n968), .A3(new_n987), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n765), .B1(new_n1102), .B2(new_n985), .ZN(new_n1103));
  OAI211_X1 g678(.A(KEYINPUT117), .B(new_n621), .C1(new_n1103), .C2(new_n1062), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1105), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1099), .B1(new_n1106), .B2(new_n1093), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1091), .A2(new_n1101), .A3(new_n1104), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1108), .A2(KEYINPUT120), .A3(new_n1094), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1098), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1060), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT125), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT62), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1113), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1040), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1115), .A2(KEYINPUT62), .A3(new_n1038), .A4(new_n1036), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1054), .A2(new_n1002), .A3(new_n1028), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1112), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1118), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1120), .A2(KEYINPUT125), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1123));
  AND4_X1   g698(.A1(new_n1014), .A2(new_n1012), .A3(new_n586), .A4(new_n588), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n1009), .B(KEYINPUT115), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1011), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1126), .B1(new_n1002), .B2(new_n1021), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT63), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1037), .A2(G8), .A3(G168), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1128), .B1(new_n1029), .B2(new_n1129), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n1021), .A2(new_n1129), .A3(new_n1128), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n991), .A2(G8), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n1131), .B(new_n1002), .C1(new_n1132), .C2(new_n997), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1127), .B1(new_n1130), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1111), .A2(new_n1123), .A3(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n972), .A2(new_n967), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n735), .B(new_n738), .ZN(new_n1137));
  XOR2_X1   g712(.A(new_n1137), .B(KEYINPUT106), .Z(new_n1138));
  XNOR2_X1  g713(.A(new_n749), .B(G1996), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n786), .B(G2067), .ZN(new_n1140));
  OR2_X1    g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1138), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(G1986), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n724), .A2(new_n1144), .ZN(new_n1145));
  XOR2_X1   g720(.A(new_n1145), .B(KEYINPUT105), .Z(new_n1146));
  INV_X1    g721(.A(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1147), .B1(new_n1144), .B2(new_n724), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1136), .B1(new_n1143), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1135), .A2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1136), .B1(new_n1140), .B2(new_n749), .ZN(new_n1151));
  NOR3_X1   g726(.A1(new_n972), .A2(G1996), .A3(new_n967), .ZN(new_n1152));
  XOR2_X1   g727(.A(new_n1152), .B(KEYINPUT46), .Z(new_n1153));
  NAND2_X1  g728(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  XOR2_X1   g729(.A(new_n1154), .B(KEYINPUT47), .Z(new_n1155));
  NAND2_X1  g730(.A1(new_n736), .A2(new_n738), .ZN(new_n1156));
  OAI22_X1  g731(.A1(new_n1141), .A2(new_n1156), .B1(G2067), .B2(new_n786), .ZN(new_n1157));
  AND2_X1   g732(.A1(new_n1157), .A2(new_n1136), .ZN(new_n1158));
  AOI21_X1  g733(.A(KEYINPUT126), .B1(new_n1143), .B2(new_n1136), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1146), .A2(new_n1136), .ZN(new_n1160));
  XOR2_X1   g735(.A(new_n1160), .B(KEYINPUT48), .Z(new_n1161));
  NOR2_X1   g736(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1143), .A2(KEYINPUT126), .A3(new_n1136), .ZN(new_n1163));
  AOI211_X1 g738(.A(new_n1155), .B(new_n1158), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1150), .A2(new_n1164), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g740(.A(KEYINPUT127), .ZN(new_n1167));
  NAND2_X1  g741(.A1(new_n951), .A2(new_n955), .ZN(new_n1168));
  NOR2_X1   g742(.A1(new_n458), .A2(G227), .ZN(new_n1169));
  NAND2_X1  g743(.A1(new_n666), .A2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g744(.A1(G229), .A2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g745(.A(new_n1171), .B1(new_n887), .B2(new_n888), .ZN(new_n1172));
  INV_X1    g746(.A(new_n1172), .ZN(new_n1173));
  AOI21_X1  g747(.A(new_n1167), .B1(new_n1168), .B2(new_n1173), .ZN(new_n1174));
  AOI211_X1 g748(.A(KEYINPUT127), .B(new_n1172), .C1(new_n951), .C2(new_n955), .ZN(new_n1175));
  NOR2_X1   g749(.A1(new_n1174), .A2(new_n1175), .ZN(G308));
  NAND2_X1  g750(.A1(new_n1168), .A2(new_n1173), .ZN(G225));
endmodule


