

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592;

  NOR2_X1 U325 ( .A1(n587), .A2(n504), .ZN(n505) );
  XOR2_X1 U326 ( .A(n347), .B(G64GAT), .Z(n429) );
  XNOR2_X1 U327 ( .A(n490), .B(n489), .ZN(n491) );
  INV_X1 U328 ( .A(n429), .ZN(n348) );
  XNOR2_X1 U329 ( .A(n376), .B(n341), .ZN(n345) );
  XNOR2_X1 U330 ( .A(KEYINPUT55), .B(n441), .ZN(n579) );
  XNOR2_X1 U331 ( .A(n389), .B(n388), .ZN(n587) );
  XNOR2_X1 U332 ( .A(n508), .B(n507), .ZN(n519) );
  XOR2_X1 U333 ( .A(n432), .B(KEYINPUT94), .Z(n293) );
  INV_X1 U334 ( .A(KEYINPUT78), .ZN(n377) );
  XNOR2_X1 U335 ( .A(KEYINPUT54), .B(KEYINPUT120), .ZN(n438) );
  XNOR2_X1 U336 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U337 ( .A(n340), .B(KEYINPUT31), .ZN(n341) );
  INV_X1 U338 ( .A(KEYINPUT96), .ZN(n489) );
  XNOR2_X1 U339 ( .A(n380), .B(n379), .ZN(n383) );
  XNOR2_X1 U340 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U341 ( .A(n351), .B(n350), .ZN(n415) );
  XNOR2_X1 U342 ( .A(n466), .B(KEYINPUT123), .ZN(n590) );
  XOR2_X1 U343 ( .A(n372), .B(n371), .Z(n582) );
  NOR2_X1 U344 ( .A1(n519), .A2(n516), .ZN(n517) );
  XOR2_X1 U345 ( .A(n436), .B(n435), .Z(n536) );
  XNOR2_X1 U346 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U347 ( .A(n470), .B(n469), .ZN(G1353GAT) );
  XOR2_X1 U348 ( .A(G204GAT), .B(KEYINPUT22), .Z(n295) );
  XNOR2_X1 U349 ( .A(KEYINPUT23), .B(G78GAT), .ZN(n294) );
  XNOR2_X1 U350 ( .A(n295), .B(n294), .ZN(n310) );
  XOR2_X1 U351 ( .A(KEYINPUT85), .B(KEYINPUT84), .Z(n297) );
  XOR2_X1 U352 ( .A(G106GAT), .B(G148GAT), .Z(n346) );
  XOR2_X1 U353 ( .A(G22GAT), .B(G155GAT), .Z(n375) );
  XNOR2_X1 U354 ( .A(n346), .B(n375), .ZN(n296) );
  XNOR2_X1 U355 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U356 ( .A(G50GAT), .B(G162GAT), .Z(n398) );
  XOR2_X1 U357 ( .A(n298), .B(n398), .Z(n308) );
  XNOR2_X1 U358 ( .A(G211GAT), .B(KEYINPUT86), .ZN(n299) );
  XNOR2_X1 U359 ( .A(n299), .B(KEYINPUT21), .ZN(n300) );
  XOR2_X1 U360 ( .A(n300), .B(KEYINPUT87), .Z(n302) );
  XNOR2_X1 U361 ( .A(G197GAT), .B(G218GAT), .ZN(n301) );
  XNOR2_X1 U362 ( .A(n302), .B(n301), .ZN(n427) );
  XNOR2_X1 U363 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n303) );
  XNOR2_X1 U364 ( .A(n303), .B(KEYINPUT2), .ZN(n331) );
  XOR2_X1 U365 ( .A(n331), .B(KEYINPUT24), .Z(n305) );
  NAND2_X1 U366 ( .A1(G228GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U367 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U368 ( .A(n427), .B(n306), .ZN(n307) );
  XNOR2_X1 U369 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U370 ( .A(n310), .B(n309), .Z(n485) );
  XOR2_X1 U371 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n312) );
  XNOR2_X1 U372 ( .A(G1GAT), .B(KEYINPUT88), .ZN(n311) );
  XNOR2_X1 U373 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U374 ( .A(G57GAT), .B(KEYINPUT5), .Z(n314) );
  XNOR2_X1 U375 ( .A(KEYINPUT92), .B(KEYINPUT4), .ZN(n313) );
  XNOR2_X1 U376 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U377 ( .A(n316), .B(n315), .Z(n321) );
  XOR2_X1 U378 ( .A(KEYINPUT89), .B(KEYINPUT90), .Z(n318) );
  NAND2_X1 U379 ( .A1(G225GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U380 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U381 ( .A(KEYINPUT91), .B(n319), .ZN(n320) );
  XNOR2_X1 U382 ( .A(n321), .B(n320), .ZN(n328) );
  XOR2_X1 U383 ( .A(G155GAT), .B(G148GAT), .Z(n323) );
  XNOR2_X1 U384 ( .A(G120GAT), .B(G127GAT), .ZN(n322) );
  XNOR2_X1 U385 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U386 ( .A(G29GAT), .B(G85GAT), .Z(n401) );
  XOR2_X1 U387 ( .A(n324), .B(n401), .Z(n326) );
  XNOR2_X1 U388 ( .A(G134GAT), .B(G162GAT), .ZN(n325) );
  XNOR2_X1 U389 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U390 ( .A(n328), .B(n327), .Z(n333) );
  XOR2_X1 U391 ( .A(KEYINPUT80), .B(KEYINPUT0), .Z(n330) );
  XNOR2_X1 U392 ( .A(G113GAT), .B(KEYINPUT79), .ZN(n329) );
  XNOR2_X1 U393 ( .A(n330), .B(n329), .ZN(n442) );
  XNOR2_X1 U394 ( .A(n442), .B(n331), .ZN(n332) );
  XOR2_X1 U395 ( .A(n333), .B(n332), .Z(n509) );
  INV_X1 U396 ( .A(n509), .ZN(n534) );
  INV_X1 U397 ( .A(KEYINPUT41), .ZN(n352) );
  XNOR2_X1 U398 ( .A(G71GAT), .B(G78GAT), .ZN(n339) );
  INV_X1 U399 ( .A(KEYINPUT13), .ZN(n334) );
  NAND2_X1 U400 ( .A1(n334), .A2(G57GAT), .ZN(n337) );
  INV_X1 U401 ( .A(G57GAT), .ZN(n335) );
  NAND2_X1 U402 ( .A1(n335), .A2(KEYINPUT13), .ZN(n336) );
  NAND2_X1 U403 ( .A1(n337), .A2(n336), .ZN(n338) );
  XNOR2_X1 U404 ( .A(n339), .B(n338), .ZN(n376) );
  AND2_X1 U405 ( .A1(G230GAT), .A2(G233GAT), .ZN(n340) );
  XOR2_X1 U406 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n343) );
  XNOR2_X1 U407 ( .A(G176GAT), .B(G85GAT), .ZN(n342) );
  XNOR2_X1 U408 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U409 ( .A(n345), .B(n344), .ZN(n351) );
  XOR2_X1 U410 ( .A(G99GAT), .B(G120GAT), .Z(n446) );
  XOR2_X1 U411 ( .A(n446), .B(n346), .Z(n349) );
  XNOR2_X1 U412 ( .A(G204GAT), .B(G92GAT), .ZN(n347) );
  XNOR2_X1 U413 ( .A(n352), .B(n415), .ZN(n567) );
  XOR2_X1 U414 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n354) );
  XNOR2_X1 U415 ( .A(G8GAT), .B(KEYINPUT70), .ZN(n353) );
  XNOR2_X1 U416 ( .A(n354), .B(n353), .ZN(n359) );
  XNOR2_X1 U417 ( .A(G1GAT), .B(KEYINPUT73), .ZN(n355) );
  XNOR2_X1 U418 ( .A(n355), .B(KEYINPUT74), .ZN(n381) );
  XOR2_X1 U419 ( .A(n381), .B(G29GAT), .Z(n357) );
  XOR2_X1 U420 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n409) );
  XNOR2_X1 U421 ( .A(G36GAT), .B(n409), .ZN(n356) );
  XNOR2_X1 U422 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U423 ( .A(n359), .B(n358), .ZN(n372) );
  XOR2_X1 U424 ( .A(G22GAT), .B(G141GAT), .Z(n361) );
  XNOR2_X1 U425 ( .A(G50GAT), .B(G43GAT), .ZN(n360) );
  XNOR2_X1 U426 ( .A(n361), .B(n360), .ZN(n365) );
  XOR2_X1 U427 ( .A(G113GAT), .B(G15GAT), .Z(n363) );
  XNOR2_X1 U428 ( .A(G169GAT), .B(G197GAT), .ZN(n362) );
  XNOR2_X1 U429 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U430 ( .A(n365), .B(n364), .Z(n370) );
  XOR2_X1 U431 ( .A(KEYINPUT75), .B(KEYINPUT72), .Z(n367) );
  NAND2_X1 U432 ( .A1(G229GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U433 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U434 ( .A(KEYINPUT71), .B(n368), .ZN(n369) );
  XNOR2_X1 U435 ( .A(n370), .B(n369), .ZN(n371) );
  NAND2_X1 U436 ( .A1(n567), .A2(n582), .ZN(n373) );
  XNOR2_X1 U437 ( .A(n373), .B(KEYINPUT109), .ZN(n374) );
  XNOR2_X1 U438 ( .A(n374), .B(KEYINPUT46), .ZN(n390) );
  XOR2_X1 U439 ( .A(n376), .B(n375), .Z(n380) );
  NAND2_X1 U440 ( .A1(G231GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U441 ( .A(n381), .B(KEYINPUT12), .ZN(n382) );
  XNOR2_X1 U442 ( .A(n383), .B(n382), .ZN(n387) );
  XOR2_X1 U443 ( .A(G64GAT), .B(KEYINPUT14), .Z(n385) );
  XNOR2_X1 U444 ( .A(G211GAT), .B(KEYINPUT15), .ZN(n384) );
  XNOR2_X1 U445 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U446 ( .A(n387), .B(n386), .Z(n389) );
  XOR2_X1 U447 ( .A(G15GAT), .B(G127GAT), .Z(n445) );
  XOR2_X1 U448 ( .A(G8GAT), .B(G183GAT), .Z(n433) );
  XNOR2_X1 U449 ( .A(n445), .B(n433), .ZN(n388) );
  XNOR2_X1 U450 ( .A(KEYINPUT108), .B(n587), .ZN(n574) );
  NOR2_X1 U451 ( .A1(n390), .A2(n574), .ZN(n391) );
  XNOR2_X1 U452 ( .A(n391), .B(KEYINPUT110), .ZN(n412) );
  XOR2_X1 U453 ( .A(KEYINPUT77), .B(KEYINPUT67), .Z(n393) );
  XNOR2_X1 U454 ( .A(G218GAT), .B(KEYINPUT69), .ZN(n392) );
  XNOR2_X1 U455 ( .A(n393), .B(n392), .ZN(n397) );
  XOR2_X1 U456 ( .A(G92GAT), .B(KEYINPUT10), .Z(n395) );
  XNOR2_X1 U457 ( .A(G99GAT), .B(G106GAT), .ZN(n394) );
  XNOR2_X1 U458 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U459 ( .A(n397), .B(n396), .Z(n400) );
  XOR2_X1 U460 ( .A(G43GAT), .B(G134GAT), .Z(n449) );
  XNOR2_X1 U461 ( .A(n449), .B(n398), .ZN(n399) );
  XNOR2_X1 U462 ( .A(n400), .B(n399), .ZN(n405) );
  XOR2_X1 U463 ( .A(G36GAT), .B(G190GAT), .Z(n428) );
  XOR2_X1 U464 ( .A(n428), .B(n401), .Z(n403) );
  NAND2_X1 U465 ( .A1(G232GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U466 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U467 ( .A(n405), .B(n404), .Z(n411) );
  XOR2_X1 U468 ( .A(KEYINPUT65), .B(KEYINPUT9), .Z(n407) );
  XNOR2_X1 U469 ( .A(KEYINPUT76), .B(KEYINPUT11), .ZN(n406) );
  XNOR2_X1 U470 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U471 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U472 ( .A(n411), .B(n410), .Z(n577) );
  INV_X1 U473 ( .A(n577), .ZN(n475) );
  NAND2_X1 U474 ( .A1(n412), .A2(n475), .ZN(n413) );
  XNOR2_X1 U475 ( .A(n413), .B(KEYINPUT111), .ZN(n414) );
  XNOR2_X1 U476 ( .A(n414), .B(KEYINPUT47), .ZN(n421) );
  XOR2_X1 U477 ( .A(KEYINPUT36), .B(n475), .Z(n589) );
  NAND2_X1 U478 ( .A1(n589), .A2(n587), .ZN(n416) );
  XNOR2_X1 U479 ( .A(n416), .B(KEYINPUT45), .ZN(n417) );
  XNOR2_X1 U480 ( .A(n417), .B(KEYINPUT68), .ZN(n418) );
  NOR2_X1 U481 ( .A1(n415), .A2(n418), .ZN(n419) );
  INV_X1 U482 ( .A(n582), .ZN(n521) );
  NAND2_X1 U483 ( .A1(n419), .A2(n521), .ZN(n420) );
  NAND2_X1 U484 ( .A1(n421), .A2(n420), .ZN(n423) );
  XNOR2_X1 U485 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n422) );
  XNOR2_X1 U486 ( .A(n423), .B(n422), .ZN(n545) );
  XOR2_X1 U487 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n425) );
  XNOR2_X1 U488 ( .A(KEYINPUT18), .B(G176GAT), .ZN(n424) );
  XNOR2_X1 U489 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U490 ( .A(G169GAT), .B(n426), .Z(n454) );
  XNOR2_X1 U491 ( .A(n454), .B(n427), .ZN(n436) );
  XNOR2_X1 U492 ( .A(n429), .B(n428), .ZN(n431) );
  NAND2_X1 U493 ( .A1(G226GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U494 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U495 ( .A(n433), .B(KEYINPUT93), .ZN(n434) );
  XNOR2_X1 U496 ( .A(n293), .B(n434), .ZN(n435) );
  XOR2_X1 U497 ( .A(KEYINPUT119), .B(n536), .Z(n437) );
  NAND2_X1 U498 ( .A1(n545), .A2(n437), .ZN(n439) );
  XNOR2_X1 U499 ( .A(n439), .B(n438), .ZN(n440) );
  NOR2_X1 U500 ( .A1(n534), .A2(n440), .ZN(n464) );
  NAND2_X1 U501 ( .A1(n485), .A2(n464), .ZN(n441) );
  XOR2_X1 U502 ( .A(G71GAT), .B(n442), .Z(n444) );
  NAND2_X1 U503 ( .A1(G227GAT), .A2(G233GAT), .ZN(n443) );
  XNOR2_X1 U504 ( .A(n444), .B(n443), .ZN(n458) );
  XOR2_X1 U505 ( .A(G183GAT), .B(G190GAT), .Z(n448) );
  XNOR2_X1 U506 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U507 ( .A(n448), .B(n447), .ZN(n450) );
  XOR2_X1 U508 ( .A(n450), .B(n449), .Z(n456) );
  XOR2_X1 U509 ( .A(KEYINPUT81), .B(KEYINPUT20), .Z(n452) );
  XNOR2_X1 U510 ( .A(KEYINPUT82), .B(KEYINPUT66), .ZN(n451) );
  XNOR2_X1 U511 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U512 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U513 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U514 ( .A(n458), .B(n457), .ZN(n516) );
  INV_X1 U515 ( .A(n516), .ZN(n576) );
  AND2_X1 U516 ( .A1(n576), .A2(n582), .ZN(n459) );
  AND2_X1 U517 ( .A1(n579), .A2(n459), .ZN(n461) );
  XNOR2_X1 U518 ( .A(KEYINPUT121), .B(G169GAT), .ZN(n460) );
  XNOR2_X1 U519 ( .A(n461), .B(n460), .ZN(G1348GAT) );
  NOR2_X1 U520 ( .A1(n576), .A2(n485), .ZN(n462) );
  XOR2_X1 U521 ( .A(KEYINPUT97), .B(n462), .Z(n463) );
  XOR2_X1 U522 ( .A(KEYINPUT26), .B(n463), .Z(n561) );
  INV_X1 U523 ( .A(n561), .ZN(n465) );
  NAND2_X1 U524 ( .A1(n465), .A2(n464), .ZN(n466) );
  NAND2_X1 U525 ( .A1(n590), .A2(n415), .ZN(n470) );
  XOR2_X1 U526 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n468) );
  XOR2_X1 U527 ( .A(G204GAT), .B(KEYINPUT125), .Z(n467) );
  AND2_X1 U528 ( .A1(n579), .A2(n576), .ZN(n573) );
  AND2_X1 U529 ( .A1(n567), .A2(n573), .ZN(n474) );
  XOR2_X1 U530 ( .A(KEYINPUT122), .B(KEYINPUT57), .Z(n472) );
  XNOR2_X1 U531 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n471) );
  XOR2_X1 U532 ( .A(n472), .B(n471), .Z(n473) );
  XNOR2_X1 U533 ( .A(n474), .B(n473), .ZN(G1349GAT) );
  XOR2_X1 U534 ( .A(KEYINPUT34), .B(KEYINPUT100), .Z(n495) );
  OR2_X1 U535 ( .A1(n415), .A2(n521), .ZN(n506) );
  NAND2_X1 U536 ( .A1(n475), .A2(n587), .ZN(n476) );
  XOR2_X1 U537 ( .A(KEYINPUT16), .B(n476), .Z(n493) );
  NAND2_X1 U538 ( .A1(n576), .A2(n536), .ZN(n477) );
  NAND2_X1 U539 ( .A1(n485), .A2(n477), .ZN(n478) );
  XNOR2_X1 U540 ( .A(n478), .B(KEYINPUT25), .ZN(n480) );
  XOR2_X1 U541 ( .A(n536), .B(KEYINPUT27), .Z(n484) );
  NOR2_X1 U542 ( .A1(n484), .A2(n561), .ZN(n479) );
  NOR2_X1 U543 ( .A1(n480), .A2(n479), .ZN(n481) );
  XNOR2_X1 U544 ( .A(n481), .B(KEYINPUT98), .ZN(n482) );
  NOR2_X1 U545 ( .A1(n534), .A2(n482), .ZN(n483) );
  XNOR2_X1 U546 ( .A(KEYINPUT99), .B(n483), .ZN(n492) );
  NOR2_X1 U547 ( .A1(n509), .A2(n484), .ZN(n544) );
  XOR2_X1 U548 ( .A(n485), .B(KEYINPUT28), .Z(n539) );
  INV_X1 U549 ( .A(n539), .ZN(n547) );
  NAND2_X1 U550 ( .A1(n544), .A2(n547), .ZN(n486) );
  XOR2_X1 U551 ( .A(KEYINPUT95), .B(n486), .Z(n488) );
  XNOR2_X1 U552 ( .A(n516), .B(KEYINPUT83), .ZN(n487) );
  NOR2_X1 U553 ( .A1(n488), .A2(n487), .ZN(n490) );
  NAND2_X1 U554 ( .A1(n492), .A2(n491), .ZN(n503) );
  NAND2_X1 U555 ( .A1(n493), .A2(n503), .ZN(n522) );
  NOR2_X1 U556 ( .A1(n506), .A2(n522), .ZN(n501) );
  NAND2_X1 U557 ( .A1(n501), .A2(n534), .ZN(n494) );
  XNOR2_X1 U558 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U559 ( .A(G1GAT), .B(n496), .Z(G1324GAT) );
  XOR2_X1 U560 ( .A(G8GAT), .B(KEYINPUT101), .Z(n498) );
  NAND2_X1 U561 ( .A1(n501), .A2(n536), .ZN(n497) );
  XNOR2_X1 U562 ( .A(n498), .B(n497), .ZN(G1325GAT) );
  XOR2_X1 U563 ( .A(G15GAT), .B(KEYINPUT35), .Z(n500) );
  NAND2_X1 U564 ( .A1(n501), .A2(n576), .ZN(n499) );
  XNOR2_X1 U565 ( .A(n500), .B(n499), .ZN(G1326GAT) );
  NAND2_X1 U566 ( .A1(n501), .A2(n539), .ZN(n502) );
  XNOR2_X1 U567 ( .A(n502), .B(G22GAT), .ZN(G1327GAT) );
  XNOR2_X1 U568 ( .A(KEYINPUT102), .B(KEYINPUT39), .ZN(n513) );
  NAND2_X1 U569 ( .A1(n589), .A2(n503), .ZN(n504) );
  XNOR2_X1 U570 ( .A(KEYINPUT37), .B(n505), .ZN(n533) );
  NOR2_X1 U571 ( .A1(n533), .A2(n506), .ZN(n508) );
  XNOR2_X1 U572 ( .A(KEYINPUT103), .B(KEYINPUT38), .ZN(n507) );
  NOR2_X1 U573 ( .A1(n519), .A2(n509), .ZN(n511) );
  XNOR2_X1 U574 ( .A(G29GAT), .B(KEYINPUT104), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U576 ( .A(n513), .B(n512), .ZN(G1328GAT) );
  INV_X1 U577 ( .A(n536), .ZN(n514) );
  NOR2_X1 U578 ( .A1(n514), .A2(n519), .ZN(n515) );
  XOR2_X1 U579 ( .A(G36GAT), .B(n515), .Z(G1329GAT) );
  XOR2_X1 U580 ( .A(n517), .B(KEYINPUT40), .Z(n518) );
  XNOR2_X1 U581 ( .A(G43GAT), .B(n518), .ZN(G1330GAT) );
  NOR2_X1 U582 ( .A1(n519), .A2(n547), .ZN(n520) );
  XOR2_X1 U583 ( .A(G50GAT), .B(n520), .Z(G1331GAT) );
  XNOR2_X1 U584 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n524) );
  NAND2_X1 U585 ( .A1(n521), .A2(n567), .ZN(n532) );
  NOR2_X1 U586 ( .A1(n532), .A2(n522), .ZN(n528) );
  NAND2_X1 U587 ( .A1(n534), .A2(n528), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n524), .B(n523), .ZN(G1332GAT) );
  XOR2_X1 U589 ( .A(G64GAT), .B(KEYINPUT105), .Z(n526) );
  NAND2_X1 U590 ( .A1(n528), .A2(n536), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n526), .B(n525), .ZN(G1333GAT) );
  NAND2_X1 U592 ( .A1(n528), .A2(n576), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n527), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT106), .B(KEYINPUT43), .Z(n530) );
  NAND2_X1 U595 ( .A1(n528), .A2(n539), .ZN(n529) );
  XNOR2_X1 U596 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U597 ( .A(G78GAT), .B(n531), .ZN(G1335GAT) );
  NOR2_X1 U598 ( .A1(n533), .A2(n532), .ZN(n540) );
  NAND2_X1 U599 ( .A1(n534), .A2(n540), .ZN(n535) );
  XNOR2_X1 U600 ( .A(G85GAT), .B(n535), .ZN(G1336GAT) );
  NAND2_X1 U601 ( .A1(n536), .A2(n540), .ZN(n537) );
  XNOR2_X1 U602 ( .A(n537), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U603 ( .A1(n540), .A2(n576), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n538), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT44), .B(KEYINPUT107), .Z(n542) );
  NAND2_X1 U606 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U608 ( .A(G106GAT), .B(n543), .ZN(G1339GAT) );
  XOR2_X1 U609 ( .A(G113GAT), .B(KEYINPUT113), .Z(n550) );
  NAND2_X1 U610 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U611 ( .A(n546), .B(KEYINPUT112), .ZN(n560) );
  NAND2_X1 U612 ( .A1(n576), .A2(n547), .ZN(n548) );
  NOR2_X1 U613 ( .A1(n560), .A2(n548), .ZN(n556) );
  NAND2_X1 U614 ( .A1(n556), .A2(n582), .ZN(n549) );
  XNOR2_X1 U615 ( .A(n550), .B(n549), .ZN(G1340GAT) );
  XOR2_X1 U616 ( .A(G120GAT), .B(KEYINPUT49), .Z(n552) );
  NAND2_X1 U617 ( .A1(n556), .A2(n567), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(G1341GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n554) );
  NAND2_X1 U620 ( .A1(n556), .A2(n574), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(n555) );
  XOR2_X1 U622 ( .A(G127GAT), .B(n555), .Z(G1342GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT51), .B(KEYINPUT115), .Z(n558) );
  NAND2_X1 U624 ( .A1(n556), .A2(n577), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(n559) );
  XOR2_X1 U626 ( .A(G134GAT), .B(n559), .Z(G1343GAT) );
  XNOR2_X1 U627 ( .A(G141GAT), .B(KEYINPUT116), .ZN(n563) );
  NOR2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n571) );
  NAND2_X1 U629 ( .A1(n571), .A2(n582), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(G1344GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n565) );
  XNOR2_X1 U632 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n564) );
  XNOR2_X1 U633 ( .A(n565), .B(n564), .ZN(n566) );
  XOR2_X1 U634 ( .A(KEYINPUT53), .B(n566), .Z(n569) );
  NAND2_X1 U635 ( .A1(n571), .A2(n567), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(G1345GAT) );
  NAND2_X1 U637 ( .A1(n571), .A2(n587), .ZN(n570) );
  XNOR2_X1 U638 ( .A(n570), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U639 ( .A1(n577), .A2(n571), .ZN(n572) );
  XNOR2_X1 U640 ( .A(n572), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U641 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n575), .B(G183GAT), .ZN(G1350GAT) );
  AND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n580), .B(KEYINPUT58), .ZN(n581) );
  XNOR2_X1 U646 ( .A(G190GAT), .B(n581), .ZN(G1351GAT) );
  NAND2_X1 U647 ( .A1(n582), .A2(n590), .ZN(n586) );
  XOR2_X1 U648 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n584) );
  XNOR2_X1 U649 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(G1352GAT) );
  NAND2_X1 U652 ( .A1(n590), .A2(n587), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n588), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U655 ( .A(n591), .B(KEYINPUT62), .ZN(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

