//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 1 1 0 1 1 1 0 1 1 0 0 0 1 0 1 0 1 0 1 0 0 1 1 0 0 0 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 0 1 1 1 1 0 0 1 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n740, new_n742, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n991, new_n992, new_n993;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT11), .ZN(new_n204));
  INV_X1    g003(.A(G169gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(KEYINPUT12), .ZN(new_n207));
  XNOR2_X1  g006(.A(G15gat), .B(G22gat), .ZN(new_n208));
  INV_X1    g007(.A(G1gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT16), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(G1gat), .B2(new_n208), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G8gat), .ZN(new_n213));
  INV_X1    g012(.A(G8gat), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n211), .B(new_n214), .C1(G1gat), .C2(new_n208), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G43gat), .B(G50gat), .ZN(new_n217));
  OR2_X1    g016(.A1(new_n217), .A2(KEYINPUT15), .ZN(new_n218));
  NAND2_X1  g017(.A1(G29gat), .A2(G36gat), .ZN(new_n219));
  XOR2_X1   g018(.A(new_n219), .B(KEYINPUT81), .Z(new_n220));
  NOR2_X1   g019(.A1(G29gat), .A2(G36gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT14), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n221), .B(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n217), .A2(KEYINPUT15), .ZN(new_n224));
  NAND4_X1  g023(.A1(new_n218), .A2(new_n220), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n221), .B(KEYINPUT14), .ZN(new_n226));
  INV_X1    g025(.A(new_n219), .ZN(new_n227));
  OAI211_X1 g026(.A(KEYINPUT15), .B(new_n217), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n216), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT83), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT83), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n216), .A2(new_n229), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n216), .A2(new_n229), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(G229gat), .A2(G233gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n238), .B(KEYINPUT13), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n237), .A2(KEYINPUT85), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT85), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n235), .B1(new_n231), .B2(new_n233), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n242), .B1(new_n243), .B2(new_n239), .ZN(new_n244));
  INV_X1    g043(.A(new_n216), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT82), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT17), .B1(new_n229), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT17), .ZN(new_n248));
  AOI211_X1 g047(.A(KEYINPUT82), .B(new_n248), .C1(new_n225), .C2(new_n228), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n245), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n234), .A2(new_n250), .A3(KEYINPUT18), .A4(new_n238), .ZN(new_n251));
  AND3_X1   g050(.A1(new_n241), .A2(new_n244), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n207), .B1(new_n252), .B2(KEYINPUT84), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n234), .A2(new_n250), .A3(new_n238), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT18), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n252), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n252), .B(new_n256), .C1(KEYINPUT84), .C2(new_n207), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(G230gat), .ZN(new_n262));
  INV_X1    g061(.A(G233gat), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT10), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT93), .ZN(new_n266));
  OR2_X1    g065(.A1(G99gat), .A2(G106gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(G99gat), .A2(G106gat), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n267), .A2(new_n266), .A3(new_n268), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n270), .A2(KEYINPUT96), .A3(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G57gat), .B(G64gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(G71gat), .A2(G78gat), .ZN(new_n274));
  NOR2_X1   g073(.A1(G71gat), .A2(G78gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(KEYINPUT9), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n273), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(G64gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(G57gat), .ZN(new_n280));
  INV_X1    g079(.A(G57gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(G64gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT9), .ZN(new_n284));
  INV_X1    g083(.A(new_n274), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n285), .A2(new_n275), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT86), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT9), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n288), .B1(new_n280), .B2(new_n282), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT86), .ZN(new_n290));
  XNOR2_X1  g089(.A(G71gat), .B(G78gat), .ZN(new_n291));
  NOR3_X1   g090(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n272), .B(new_n278), .C1(new_n287), .C2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(KEYINPUT92), .A2(KEYINPUT7), .ZN(new_n294));
  INV_X1    g093(.A(G85gat), .ZN(new_n295));
  INV_X1    g094(.A(G92gat), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND4_X1  g096(.A1(KEYINPUT92), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AOI22_X1  g098(.A1(KEYINPUT8), .A2(new_n268), .B1(new_n295), .B2(new_n296), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n270), .A2(new_n299), .A3(new_n271), .A4(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n300), .A2(new_n297), .A3(new_n298), .ZN(new_n302));
  INV_X1    g101(.A(new_n271), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n302), .B1(new_n303), .B2(new_n269), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n293), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n290), .B1(new_n289), .B2(new_n291), .ZN(new_n307));
  OAI211_X1 g106(.A(new_n286), .B(KEYINPUT86), .C1(new_n273), .C2(new_n288), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n277), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  AOI22_X1  g108(.A1(new_n309), .A2(new_n272), .B1(new_n301), .B2(new_n304), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n265), .B1(new_n306), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n305), .A2(KEYINPUT10), .A3(new_n309), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n264), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n264), .ZN(new_n314));
  NOR3_X1   g113(.A1(new_n306), .A2(new_n310), .A3(new_n314), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G120gat), .B(G148gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n317), .B(KEYINPUT97), .ZN(new_n318));
  INV_X1    g117(.A(G176gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n318), .B(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(G204gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n320), .B(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n316), .B(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n261), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(G155gat), .ZN(new_n326));
  INV_X1    g125(.A(G162gat), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n326), .A2(new_n327), .A3(KEYINPUT71), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT71), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n329), .B1(G155gat), .B2(G162gat), .ZN(new_n330));
  AND2_X1   g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT2), .ZN(new_n332));
  INV_X1    g131(.A(G141gat), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n333), .A2(G148gat), .ZN(new_n334));
  INV_X1    g133(.A(G148gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n335), .A2(G141gat), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n332), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  AND2_X1   g136(.A1(G155gat), .A2(G162gat), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n331), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  NOR2_X1   g139(.A1(G155gat), .A2(G162gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(new_n332), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(new_n339), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n333), .A2(KEYINPUT72), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT72), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(G141gat), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n335), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n343), .B1(new_n347), .B2(new_n334), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n340), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT1), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n350), .B1(G113gat), .B2(G120gat), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(G127gat), .ZN(new_n353));
  INV_X1    g152(.A(G134gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(G127gat), .A2(G134gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(G113gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT68), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT68), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(G113gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(G120gat), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n352), .B(new_n357), .C1(new_n362), .C2(new_n363), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n358), .A2(new_n363), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n355), .B(new_n356), .C1(new_n365), .C2(new_n351), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NOR3_X1   g166(.A1(new_n349), .A2(KEYINPUT4), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(KEYINPUT75), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n335), .A2(G141gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n333), .A2(G148gat), .ZN(new_n371));
  AOI21_X1  g170(.A(KEYINPUT2), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n372), .A2(new_n338), .ZN(new_n373));
  XNOR2_X1  g172(.A(KEYINPUT72), .B(G141gat), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n370), .B1(new_n374), .B2(new_n335), .ZN(new_n375));
  AOI22_X1  g174(.A1(new_n373), .A2(new_n331), .B1(new_n375), .B2(new_n343), .ZN(new_n376));
  AND2_X1   g175(.A1(new_n364), .A2(new_n366), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT4), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT75), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT4), .B1(new_n349), .B2(new_n367), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n369), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT5), .ZN(new_n384));
  NAND2_X1  g183(.A1(G225gat), .A2(G233gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n328), .A2(new_n330), .ZN(new_n386));
  NOR3_X1   g185(.A1(new_n372), .A2(new_n386), .A3(new_n338), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n338), .B1(new_n332), .B2(new_n341), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n345), .A2(G141gat), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n333), .A2(KEYINPUT72), .ZN(new_n390));
  OAI21_X1  g189(.A(G148gat), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n388), .B1(new_n391), .B2(new_n370), .ZN(new_n392));
  OAI21_X1  g191(.A(KEYINPUT3), .B1(new_n387), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT3), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n340), .A2(new_n394), .A3(new_n348), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n393), .A2(new_n367), .A3(new_n395), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n383), .A2(new_n384), .A3(new_n385), .A4(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n397), .B(KEYINPUT76), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT74), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n378), .B1(new_n376), .B2(new_n377), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n396), .B(new_n385), .C1(new_n368), .C2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT73), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n382), .A2(new_n379), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n404), .A2(KEYINPUT73), .A3(new_n385), .A4(new_n396), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n349), .B(new_n367), .ZN(new_n407));
  INV_X1    g206(.A(new_n385), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AND4_X1   g208(.A1(new_n399), .A2(new_n406), .A3(KEYINPUT5), .A4(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n384), .B1(new_n403), .B2(new_n405), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n399), .B1(new_n411), .B2(new_n409), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n398), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(G1gat), .B(G29gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n414), .B(KEYINPUT0), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n415), .B(G57gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n416), .B(G85gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n413), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT6), .ZN(new_n419));
  INV_X1    g218(.A(new_n417), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n420), .B(new_n398), .C1(new_n410), .C2(new_n412), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n418), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n413), .A2(KEYINPUT6), .A3(new_n417), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G8gat), .B(G36gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n425), .B(new_n279), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n426), .B(new_n296), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(G197gat), .B(G204gat), .ZN(new_n429));
  NAND2_X1  g228(.A1(G211gat), .A2(G218gat), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n429), .B1(KEYINPUT22), .B2(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(G211gat), .B(G218gat), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n433), .A2(KEYINPUT69), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  OAI221_X1 g234(.A(new_n429), .B1(new_n431), .B2(KEYINPUT22), .C1(new_n433), .C2(KEYINPUT69), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(G226gat), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n438), .A2(new_n263), .ZN(new_n439));
  INV_X1    g238(.A(G183gat), .ZN(new_n440));
  OAI21_X1  g239(.A(KEYINPUT27), .B1(new_n440), .B2(KEYINPUT65), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT65), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT27), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n442), .A2(new_n443), .A3(G183gat), .ZN(new_n444));
  INV_X1    g243(.A(G190gat), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n441), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT66), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT28), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n441), .A2(new_n444), .A3(KEYINPUT66), .A4(new_n445), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  AND2_X1   g250(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n452));
  NOR2_X1   g251(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n453));
  OAI211_X1 g252(.A(KEYINPUT28), .B(new_n445), .C1(new_n452), .C2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT67), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g255(.A(KEYINPUT27), .B(G183gat), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n457), .A2(KEYINPUT67), .A3(KEYINPUT28), .A4(new_n445), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n451), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g259(.A1(G169gat), .A2(G176gat), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT26), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(G169gat), .A2(G176gat), .ZN(new_n464));
  OAI21_X1  g263(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(G183gat), .A2(G190gat), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n460), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NOR2_X1   g267(.A1(KEYINPUT64), .A2(KEYINPUT25), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n440), .A2(new_n445), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n470), .A2(KEYINPUT24), .A3(new_n467), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT24), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n472), .A2(G183gat), .A3(G190gat), .ZN(new_n473));
  AND3_X1   g272(.A1(new_n471), .A2(new_n464), .A3(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT23), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n461), .B(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n469), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n473), .A2(new_n464), .ZN(new_n478));
  AND4_X1   g277(.A1(new_n476), .A2(new_n478), .A3(new_n471), .A4(new_n469), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT64), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT25), .ZN(new_n481));
  OAI22_X1  g280(.A1(new_n477), .A2(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n468), .A2(new_n482), .A3(KEYINPUT70), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(KEYINPUT70), .B1(new_n468), .B2(new_n482), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n439), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n468), .A2(new_n482), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n439), .A2(KEYINPUT29), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n437), .B1(new_n486), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT70), .ZN(new_n491));
  INV_X1    g290(.A(new_n466), .ZN(new_n492));
  INV_X1    g291(.A(new_n467), .ZN(new_n493));
  AOI211_X1 g292(.A(new_n492), .B(new_n493), .C1(new_n451), .C2(new_n459), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n480), .A2(new_n481), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n476), .A2(new_n478), .A3(new_n471), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n496), .B1(KEYINPUT64), .B2(KEYINPUT25), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n474), .A2(new_n476), .A3(new_n469), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n495), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n491), .B1(new_n494), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n500), .A2(new_n483), .A3(new_n488), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n494), .A2(new_n499), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(new_n439), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n501), .A2(new_n437), .A3(new_n503), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n428), .B1(new_n490), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n437), .ZN(new_n506));
  INV_X1    g305(.A(new_n439), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n507), .B1(new_n500), .B2(new_n483), .ZN(new_n508));
  INV_X1    g307(.A(new_n489), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n506), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n501), .A2(new_n437), .A3(new_n503), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n510), .A2(new_n427), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n505), .A2(KEYINPUT30), .A3(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT30), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n514), .B(new_n428), .C1(new_n490), .C2(new_n504), .ZN(new_n515));
  AND2_X1   g314(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT29), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n395), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(new_n506), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT77), .ZN(new_n521));
  AOI21_X1  g320(.A(KEYINPUT29), .B1(new_n432), .B2(new_n433), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n522), .B1(new_n432), .B2(new_n433), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(new_n394), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(new_n349), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n437), .B1(new_n395), .B2(new_n518), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT77), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n521), .A2(new_n525), .A3(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(G228gat), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n530), .A2(new_n263), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT78), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n532), .B1(new_n520), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n394), .B1(new_n506), .B2(KEYINPUT29), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(new_n349), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n526), .A2(KEYINPUT78), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n535), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n533), .A2(KEYINPUT79), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(G22gat), .ZN(new_n541));
  INV_X1    g340(.A(G22gat), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n533), .A2(KEYINPUT79), .A3(new_n542), .A4(new_n539), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n533), .A2(new_n539), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT79), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  XOR2_X1   g346(.A(G78gat), .B(G106gat), .Z(new_n548));
  XNOR2_X1  g347(.A(KEYINPUT31), .B(G50gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n548), .B(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n544), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n541), .A2(new_n547), .A3(new_n550), .A4(new_n543), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(G227gat), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n555), .A2(new_n263), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n487), .A2(new_n377), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n468), .A2(new_n482), .A3(new_n367), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n557), .A2(new_n556), .A3(new_n558), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT34), .ZN(new_n561));
  AND3_X1   g360(.A1(new_n560), .A2(KEYINPUT32), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n561), .B1(new_n560), .B2(KEYINPUT32), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n559), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n560), .A2(KEYINPUT32), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(KEYINPUT34), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n560), .A2(KEYINPUT32), .A3(new_n561), .ZN(new_n567));
  INV_X1    g366(.A(new_n559), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G15gat), .B(G43gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(G71gat), .ZN(new_n571));
  INV_X1    g370(.A(G99gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT33), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n574), .B1(new_n560), .B2(new_n575), .ZN(new_n576));
  AND3_X1   g375(.A1(new_n564), .A2(new_n569), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n576), .B1(new_n564), .B2(new_n569), .ZN(new_n578));
  NOR3_X1   g377(.A1(new_n554), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  AND4_X1   g378(.A1(KEYINPUT35), .A2(new_n424), .A3(new_n517), .A4(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n516), .B1(new_n422), .B2(new_n423), .ZN(new_n581));
  AOI21_X1  g380(.A(KEYINPUT35), .B1(new_n581), .B2(new_n579), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(KEYINPUT37), .B1(new_n510), .B2(new_n511), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n510), .A2(KEYINPUT37), .A3(new_n511), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n585), .A2(KEYINPUT38), .A3(new_n586), .A4(new_n427), .ZN(new_n587));
  NOR3_X1   g386(.A1(new_n508), .A2(new_n509), .A3(new_n506), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n437), .B1(new_n501), .B2(new_n503), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT37), .ZN(new_n590));
  NOR3_X1   g389(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NOR3_X1   g390(.A1(new_n591), .A2(new_n584), .A3(new_n428), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n587), .B1(new_n592), .B2(KEYINPUT38), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n593), .A2(new_n422), .A3(new_n423), .A4(new_n505), .ZN(new_n594));
  INV_X1    g393(.A(new_n554), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n385), .B1(new_n383), .B2(new_n396), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT39), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n407), .A2(new_n408), .ZN(new_n598));
  OR3_X1    g397(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n417), .B1(new_n596), .B2(new_n597), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n599), .A2(KEYINPUT40), .A3(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT80), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  AND2_X1   g402(.A1(new_n599), .A2(new_n600), .ZN(new_n604));
  OR2_X1    g403(.A1(new_n604), .A2(KEYINPUT40), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n603), .A2(new_n516), .A3(new_n418), .A4(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n594), .A2(new_n595), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n421), .A2(new_n419), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n406), .A2(KEYINPUT5), .A3(new_n409), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(KEYINPUT74), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n411), .A2(new_n399), .A3(new_n409), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n420), .B1(new_n612), .B2(new_n398), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n423), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n517), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(new_n554), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n577), .A2(new_n578), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(KEYINPUT36), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT36), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n620), .B1(new_n577), .B2(new_n578), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n607), .A2(new_n617), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n325), .B1(new_n583), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n309), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT21), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n625), .A2(new_n216), .A3(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n245), .B1(KEYINPUT21), .B2(new_n309), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n625), .A2(new_n626), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  XOR2_X1   g429(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G127gat), .B(G155gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT89), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n632), .B(new_n634), .ZN(new_n635));
  XOR2_X1   g434(.A(G183gat), .B(G211gat), .Z(new_n636));
  XNOR2_X1  g435(.A(KEYINPUT87), .B(KEYINPUT88), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(G231gat), .A2(G233gat), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n638), .B(new_n639), .Z(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n635), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n635), .A2(new_n641), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(G232gat), .A2(G233gat), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT41), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n647), .B1(new_n229), .B2(new_n305), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n648), .B(KEYINPUT95), .Z(new_n649));
  XNOR2_X1  g448(.A(new_n305), .B(KEYINPUT94), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n650), .B1(new_n247), .B2(new_n249), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(KEYINPUT90), .B(KEYINPUT91), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n645), .A2(new_n646), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n652), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(G190gat), .B(G218gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(new_n354), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(G162gat), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n656), .B(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n644), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n624), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n663), .A2(new_n424), .ZN(new_n664));
  XOR2_X1   g463(.A(KEYINPUT98), .B(G1gat), .Z(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(G1324gat));
  NAND3_X1  g465(.A1(new_n624), .A2(new_n662), .A3(new_n516), .ZN(new_n667));
  OR2_X1    g466(.A1(new_n667), .A2(KEYINPUT99), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(KEYINPUT99), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(G8gat), .ZN(new_n671));
  XOR2_X1   g470(.A(KEYINPUT16), .B(G8gat), .Z(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(KEYINPUT42), .ZN(new_n673));
  AND3_X1   g472(.A1(new_n668), .A2(new_n669), .A3(new_n672), .ZN(new_n674));
  OAI221_X1 g473(.A(new_n671), .B1(new_n667), .B2(new_n673), .C1(new_n674), .C2(KEYINPUT42), .ZN(G1325gat));
  INV_X1    g474(.A(G15gat), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n663), .A2(new_n676), .A3(new_n622), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n624), .A2(new_n662), .A3(new_n618), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n677), .B1(new_n676), .B2(new_n678), .ZN(G1326gat));
  NAND3_X1  g478(.A1(new_n624), .A2(new_n662), .A3(new_n554), .ZN(new_n680));
  XNOR2_X1  g479(.A(KEYINPUT43), .B(G22gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(KEYINPUT100), .B(KEYINPUT101), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(G1327gat));
  INV_X1    g483(.A(new_n644), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n325), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n583), .A2(new_n623), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n687), .B1(new_n688), .B2(new_n661), .ZN(new_n689));
  INV_X1    g488(.A(new_n661), .ZN(new_n690));
  AOI211_X1 g489(.A(KEYINPUT44), .B(new_n690), .C1(new_n583), .C2(new_n623), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n686), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(G29gat), .B1(new_n692), .B2(new_n424), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n690), .B1(new_n583), .B2(new_n623), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(new_n686), .ZN(new_n695));
  OR3_X1    g494(.A1(new_n695), .A2(G29gat), .A3(new_n424), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(KEYINPUT102), .ZN(new_n697));
  OR4_X1    g496(.A1(KEYINPUT102), .A2(new_n695), .A3(G29gat), .A4(new_n424), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT45), .ZN(new_n699));
  AND3_X1   g498(.A1(new_n697), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n699), .B1(new_n697), .B2(new_n698), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n693), .B1(new_n700), .B2(new_n701), .ZN(G1328gat));
  NOR3_X1   g501(.A1(new_n695), .A2(G36gat), .A3(new_n517), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT46), .ZN(new_n704));
  OAI21_X1  g503(.A(G36gat), .B1(new_n692), .B2(new_n517), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(G1329gat));
  INV_X1    g505(.A(G43gat), .ZN(new_n707));
  INV_X1    g506(.A(new_n686), .ZN(new_n708));
  INV_X1    g507(.A(new_n689), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n687), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n622), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n707), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT47), .ZN(new_n714));
  INV_X1    g513(.A(new_n618), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n695), .A2(G43gat), .A3(new_n715), .ZN(new_n716));
  OR3_X1    g515(.A1(new_n713), .A2(new_n714), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n714), .B1(new_n713), .B2(new_n716), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(G1330gat));
  OAI21_X1  g518(.A(G50gat), .B1(new_n692), .B2(new_n595), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n695), .A2(G50gat), .A3(new_n595), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT103), .ZN(new_n724));
  AOI21_X1  g523(.A(KEYINPUT48), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n723), .B(new_n725), .ZN(G1331gat));
  AND3_X1   g525(.A1(new_n688), .A2(new_n662), .A3(new_n261), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(new_n323), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n424), .B(KEYINPUT104), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XOR2_X1   g529(.A(KEYINPUT105), .B(G57gat), .Z(new_n731));
  XNOR2_X1  g530(.A(new_n730), .B(new_n731), .ZN(G1332gat));
  NOR2_X1   g531(.A1(new_n728), .A2(new_n517), .ZN(new_n733));
  NOR2_X1   g532(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n734));
  AND2_X1   g533(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n736), .B1(new_n733), .B2(new_n734), .ZN(G1333gat));
  NOR2_X1   g536(.A1(new_n728), .A2(new_n715), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n712), .A2(G71gat), .ZN(new_n739));
  OAI22_X1  g538(.A1(new_n738), .A2(G71gat), .B1(new_n728), .B2(new_n739), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g540(.A1(new_n728), .A2(new_n595), .ZN(new_n742));
  XOR2_X1   g541(.A(new_n742), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g542(.A1(new_n685), .A2(new_n260), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n694), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT51), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n424), .A2(G85gat), .ZN(new_n748));
  AND3_X1   g547(.A1(new_n747), .A2(new_n323), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n744), .A2(new_n323), .ZN(new_n750));
  XOR2_X1   g549(.A(new_n750), .B(KEYINPUT106), .Z(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n752), .B1(new_n709), .B2(new_n710), .ZN(new_n753));
  INV_X1    g552(.A(new_n424), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n295), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(KEYINPUT107), .B1(new_n749), .B2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT107), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n747), .A2(new_n323), .A3(new_n748), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n753), .A2(new_n754), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n757), .B(new_n758), .C1(new_n759), .C2(new_n295), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n756), .A2(new_n760), .ZN(G1336gat));
  NOR2_X1   g560(.A1(new_n517), .A2(G92gat), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n747), .A2(new_n323), .A3(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT52), .ZN(new_n764));
  OAI211_X1 g563(.A(new_n516), .B(new_n751), .C1(new_n689), .C2(new_n691), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(G92gat), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n763), .A2(new_n764), .A3(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT109), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n746), .A2(KEYINPUT108), .ZN(new_n769));
  AND3_X1   g568(.A1(new_n694), .A2(new_n744), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n769), .B1(new_n694), .B2(new_n744), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n323), .B(new_n762), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n766), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n768), .B1(new_n773), .B2(KEYINPUT52), .ZN(new_n774));
  AOI211_X1 g573(.A(KEYINPUT109), .B(new_n764), .C1(new_n766), .C2(new_n772), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n767), .B1(new_n774), .B2(new_n775), .ZN(G1337gat));
  NAND3_X1  g575(.A1(new_n747), .A2(new_n323), .A3(new_n618), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n622), .A2(new_n572), .ZN(new_n778));
  AOI22_X1  g577(.A1(new_n777), .A2(new_n572), .B1(new_n753), .B2(new_n778), .ZN(G1338gat));
  NAND2_X1  g578(.A1(new_n753), .A2(new_n554), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(G106gat), .ZN(new_n781));
  INV_X1    g580(.A(new_n323), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n595), .A2(G106gat), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(KEYINPUT53), .B1(new_n747), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n781), .A2(new_n784), .ZN(new_n785));
  OR2_X1    g584(.A1(new_n770), .A2(new_n771), .ZN(new_n786));
  AOI22_X1  g585(.A1(new_n780), .A2(G106gat), .B1(new_n786), .B2(new_n783), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT53), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n785), .B1(new_n787), .B2(new_n788), .ZN(G1339gat));
  NAND3_X1  g588(.A1(new_n662), .A2(new_n782), .A3(new_n261), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT111), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n311), .A2(new_n264), .A3(new_n312), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n293), .A2(new_n305), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n309), .A2(new_n301), .A3(new_n304), .A4(new_n272), .ZN(new_n794));
  AOI21_X1  g593(.A(KEYINPUT10), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(new_n312), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n314), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n792), .A2(new_n797), .A3(KEYINPUT54), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(KEYINPUT110), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT110), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n792), .A2(new_n797), .A3(new_n800), .A4(KEYINPUT54), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n322), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n803), .B1(new_n797), .B2(KEYINPUT54), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n802), .A2(KEYINPUT55), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n316), .A2(new_n322), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n804), .B1(new_n799), .B2(new_n801), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n809), .A2(KEYINPUT55), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n791), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  OR2_X1    g610(.A1(new_n809), .A2(KEYINPUT55), .ZN(new_n812));
  INV_X1    g611(.A(new_n807), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n813), .B1(new_n809), .B2(KEYINPUT55), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n812), .A2(new_n814), .A3(KEYINPUT111), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n811), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT112), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n238), .B1(new_n234), .B2(new_n250), .ZN(new_n818));
  INV_X1    g617(.A(new_n233), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n232), .B1(new_n216), .B2(new_n229), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n236), .B(new_n239), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n817), .B(new_n206), .C1(new_n818), .C2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  AND4_X1   g623(.A1(new_n244), .A2(new_n256), .A3(new_n241), .A4(new_n251), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n824), .B1(new_n825), .B2(new_n207), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n206), .B1(new_n818), .B2(new_n822), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(KEYINPUT112), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n816), .A2(new_n661), .A3(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n252), .A2(new_n207), .A3(new_n256), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n831), .A2(new_n323), .A3(new_n828), .A4(new_n823), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT113), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n826), .A2(KEYINPUT113), .A3(new_n323), .A4(new_n828), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n836), .B1(new_n816), .B2(new_n260), .ZN(new_n837));
  OAI211_X1 g636(.A(KEYINPUT114), .B(new_n830), .C1(new_n837), .C2(new_n661), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n644), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n261), .B1(new_n811), .B2(new_n815), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n690), .B1(new_n840), .B2(new_n836), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT114), .B1(new_n841), .B2(new_n830), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n790), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n843), .A2(new_n579), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n729), .A2(new_n516), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n846), .A2(new_n362), .A3(new_n260), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT115), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n424), .A2(new_n516), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n843), .A2(new_n579), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n260), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n848), .B1(new_n851), .B2(G113gat), .ZN(new_n852));
  AOI211_X1 g651(.A(KEYINPUT115), .B(new_n358), .C1(new_n850), .C2(new_n260), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n847), .B1(new_n852), .B2(new_n853), .ZN(G1340gat));
  NAND2_X1  g653(.A1(new_n323), .A2(new_n363), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n855), .B(KEYINPUT117), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n846), .A2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT116), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n850), .A2(new_n323), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n858), .B1(new_n859), .B2(G120gat), .ZN(new_n860));
  AOI211_X1 g659(.A(KEYINPUT116), .B(new_n363), .C1(new_n850), .C2(new_n323), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n857), .B1(new_n860), .B2(new_n861), .ZN(G1341gat));
  AOI21_X1  g661(.A(G127gat), .B1(new_n846), .B2(new_n685), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n644), .A2(new_n353), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n863), .B1(new_n850), .B2(new_n864), .ZN(G1342gat));
  XNOR2_X1  g664(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n844), .A2(new_n354), .A3(new_n845), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n866), .B1(new_n867), .B2(new_n690), .ZN(new_n868));
  NAND2_X1  g667(.A1(KEYINPUT119), .A2(KEYINPUT56), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n846), .A2(new_n354), .A3(new_n661), .A4(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n850), .A2(new_n661), .ZN(new_n871));
  AND3_X1   g670(.A1(new_n871), .A2(KEYINPUT118), .A3(G134gat), .ZN(new_n872));
  AOI21_X1  g671(.A(KEYINPUT118), .B1(new_n871), .B2(G134gat), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n868), .B(new_n870), .C1(new_n872), .C2(new_n873), .ZN(G1343gat));
  AND3_X1   g673(.A1(new_n816), .A2(new_n661), .A3(new_n829), .ZN(new_n875));
  XNOR2_X1  g674(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n260), .B(new_n814), .C1(new_n809), .C2(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n661), .B1(new_n877), .B2(new_n832), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n644), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n595), .B1(new_n879), .B2(new_n790), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT57), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n622), .B(new_n849), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n843), .A2(new_n554), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n883), .B1(KEYINPUT57), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n374), .B1(new_n885), .B2(new_n261), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n884), .A2(new_n712), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n887), .A2(new_n333), .A3(new_n260), .A4(new_n845), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT58), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n886), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(new_n374), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT114), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n808), .A2(new_n791), .A3(new_n810), .ZN(new_n893));
  AOI21_X1  g692(.A(KEYINPUT111), .B1(new_n812), .B2(new_n814), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n260), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n836), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n661), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n892), .B1(new_n897), .B2(new_n875), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n644), .A3(new_n838), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n595), .B1(new_n899), .B2(new_n790), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n882), .B1(new_n900), .B2(new_n881), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n891), .B1(new_n901), .B2(new_n260), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n900), .A2(new_n622), .A3(new_n845), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n903), .A2(G141gat), .A3(new_n261), .ZN(new_n904));
  OAI21_X1  g703(.A(KEYINPUT58), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n890), .A2(new_n905), .ZN(G1344gat));
  NAND4_X1  g705(.A1(new_n887), .A2(new_n335), .A3(new_n323), .A4(new_n845), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT59), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n884), .A2(KEYINPUT57), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n595), .A2(KEYINPUT57), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n661), .A2(new_n814), .A3(new_n812), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n911), .B(KEYINPUT122), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n829), .ZN(new_n913));
  INV_X1    g712(.A(new_n878), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n685), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(new_n790), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n910), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n849), .A2(new_n622), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT121), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n909), .A2(new_n323), .A3(new_n917), .A4(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n908), .B1(new_n920), .B2(G148gat), .ZN(new_n921));
  AOI211_X1 g720(.A(KEYINPUT59), .B(new_n335), .C1(new_n901), .C2(new_n323), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n907), .B1(new_n921), .B2(new_n922), .ZN(G1345gat));
  NAND3_X1  g722(.A1(new_n887), .A2(new_n685), .A3(new_n845), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n644), .A2(new_n326), .ZN(new_n925));
  AOI22_X1  g724(.A1(new_n924), .A2(new_n326), .B1(new_n901), .B2(new_n925), .ZN(G1346gat));
  NAND3_X1  g725(.A1(new_n887), .A2(new_n661), .A3(new_n845), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n690), .A2(new_n327), .ZN(new_n928));
  AOI22_X1  g727(.A1(new_n927), .A2(new_n327), .B1(new_n901), .B2(new_n928), .ZN(G1347gat));
  AND2_X1   g728(.A1(new_n729), .A2(new_n516), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n843), .A2(new_n260), .A3(new_n579), .A4(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(G169gat), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n754), .A2(new_n517), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n844), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n260), .A2(new_n205), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n932), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT123), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n936), .B(new_n937), .ZN(G1348gat));
  INV_X1    g737(.A(new_n934), .ZN(new_n939));
  AOI21_X1  g738(.A(G176gat), .B1(new_n939), .B2(new_n323), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n844), .A2(new_n930), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n782), .A2(new_n319), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(G1349gat));
  NAND4_X1  g742(.A1(new_n843), .A2(new_n685), .A3(new_n579), .A4(new_n930), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(G183gat), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n685), .A2(new_n457), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n945), .B1(new_n934), .B2(new_n946), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g747(.A1(new_n939), .A2(new_n445), .A3(new_n661), .ZN(new_n949));
  NAND4_X1  g748(.A1(new_n843), .A2(new_n661), .A3(new_n579), .A4(new_n930), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT124), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n950), .A2(new_n951), .A3(G190gat), .ZN(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n951), .B1(new_n950), .B2(G190gat), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n953), .A2(new_n954), .A3(KEYINPUT61), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT61), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n950), .A2(G190gat), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(KEYINPUT124), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n956), .B1(new_n958), .B2(new_n952), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n949), .B1(new_n955), .B2(new_n959), .ZN(G1351gat));
  OR2_X1    g759(.A1(new_n915), .A2(new_n916), .ZN(new_n961));
  AOI22_X1  g760(.A1(new_n884), .A2(KEYINPUT57), .B1(new_n961), .B2(new_n910), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT125), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n930), .A2(new_n622), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n962), .A2(new_n963), .A3(new_n260), .A4(new_n964), .ZN(new_n965));
  OAI211_X1 g764(.A(new_n917), .B(new_n964), .C1(new_n900), .C2(new_n881), .ZN(new_n966));
  OAI21_X1  g765(.A(KEYINPUT125), .B1(new_n966), .B2(new_n261), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n965), .A2(new_n967), .A3(G197gat), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n887), .A2(new_n933), .ZN(new_n969));
  INV_X1    g768(.A(G197gat), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n969), .A2(new_n970), .A3(new_n260), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n968), .A2(new_n971), .ZN(G1352gat));
  XNOR2_X1  g771(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n973));
  INV_X1    g772(.A(new_n973), .ZN(new_n974));
  NAND4_X1  g773(.A1(new_n969), .A2(new_n321), .A3(new_n323), .A4(new_n974), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n962), .A2(new_n323), .A3(new_n964), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n976), .A2(G204gat), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n887), .A2(new_n321), .A3(new_n933), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n973), .B1(new_n978), .B2(new_n782), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n975), .A2(new_n977), .A3(new_n979), .ZN(G1353gat));
  INV_X1    g779(.A(KEYINPUT127), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n966), .A2(new_n644), .ZN(new_n982));
  INV_X1    g781(.A(G211gat), .ZN(new_n983));
  OAI211_X1 g782(.A(new_n981), .B(KEYINPUT63), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n969), .A2(new_n983), .A3(new_n685), .ZN(new_n985));
  NAND4_X1  g784(.A1(new_n909), .A2(new_n685), .A3(new_n917), .A4(new_n964), .ZN(new_n986));
  OR2_X1    g785(.A1(new_n981), .A2(KEYINPUT63), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n981), .A2(KEYINPUT63), .ZN(new_n988));
  NAND4_X1  g787(.A1(new_n986), .A2(G211gat), .A3(new_n987), .A4(new_n988), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n984), .A2(new_n985), .A3(new_n989), .ZN(G1354gat));
  INV_X1    g789(.A(G218gat), .ZN(new_n991));
  NOR3_X1   g790(.A1(new_n966), .A2(new_n991), .A3(new_n690), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n969), .A2(new_n661), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n992), .B1(new_n993), .B2(new_n991), .ZN(G1355gat));
endmodule


