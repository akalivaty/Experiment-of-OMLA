//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 0 1 1 0 0 1 0 0 1 0 0 0 0 1 1 0 0 0 0 0 1 0 0 0 0 1 1 1 0 0 0 1 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 1 0 1 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:12 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1312, new_n1313, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1375, new_n1376, new_n1377,
    new_n1378, new_n1379, new_n1380, new_n1381, new_n1382, new_n1383;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(new_n202), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G50), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(G1), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n210), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(G13), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT65), .Z(new_n218));
  INV_X1    g0018(.A(KEYINPUT0), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n212), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AOI21_X1  g0020(.A(new_n220), .B1(new_n219), .B2(new_n218), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT66), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  INV_X1    g0023(.A(G77), .ZN(new_n224));
  INV_X1    g0024(.A(G244), .ZN(new_n225));
  INV_X1    g0025(.A(G107), .ZN(new_n226));
  INV_X1    g0026(.A(G264), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n215), .B1(new_n228), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT1), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n222), .A2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  INV_X1    g0035(.A(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G264), .B(G270), .Z(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G358));
  XNOR2_X1  g0043(.A(G68), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT67), .ZN(new_n245));
  XOR2_X1   g0045(.A(G50), .B(G58), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(KEYINPUT3), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n256), .A2(G232), .A3(G1698), .ZN(new_n257));
  NAND2_X1  g0057(.A1(G33), .A2(G97), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G226), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n257), .B(new_n258), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n209), .B1(G33), .B2(G41), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G41), .ZN(new_n265));
  INV_X1    g0065(.A(G45), .ZN(new_n266));
  AOI21_X1  g0066(.A(G1), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G33), .A2(G41), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(G1), .A3(G13), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n267), .A2(new_n269), .A3(G274), .ZN(new_n270));
  INV_X1    g0070(.A(G238), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n213), .B1(G41), .B2(G45), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n270), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n264), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT13), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT75), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n274), .B1(new_n262), .B2(new_n263), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT13), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n277), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n276), .A2(new_n278), .A3(KEYINPUT13), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n282), .A2(G169), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT14), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT14), .ZN(new_n286));
  NAND4_X1  g0086(.A1(new_n282), .A2(new_n286), .A3(G169), .A4(new_n283), .ZN(new_n287));
  INV_X1    g0087(.A(G179), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n288), .B1(new_n279), .B2(new_n280), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n277), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n285), .A2(new_n287), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n209), .ZN(new_n293));
  NOR2_X1   g0093(.A1(G20), .A2(G33), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G50), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n210), .A2(G33), .ZN(new_n298));
  OAI22_X1  g0098(.A1(new_n298), .A2(new_n224), .B1(new_n210), .B2(G68), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n293), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n300), .B(KEYINPUT11), .ZN(new_n301));
  INV_X1    g0101(.A(G68), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n293), .B1(new_n213), .B2(G20), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(KEYINPUT76), .A2(KEYINPUT12), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n213), .A2(G13), .A3(G20), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(G68), .B1(KEYINPUT76), .B2(KEYINPUT12), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n305), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NOR4_X1   g0109(.A1(new_n306), .A2(KEYINPUT76), .A3(KEYINPUT12), .A4(G68), .ZN(new_n310));
  OAI221_X1 g0110(.A(new_n301), .B1(new_n302), .B2(new_n304), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n291), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G190), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n314), .B1(new_n279), .B2(new_n280), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n311), .B1(new_n315), .B2(new_n277), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n282), .A2(G200), .A3(new_n283), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n313), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n263), .A2(new_n267), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(G226), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n270), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT68), .ZN(new_n324));
  XNOR2_X1  g0124(.A(new_n323), .B(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n256), .A2(G222), .A3(new_n259), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n256), .A2(G1698), .ZN(new_n327));
  INV_X1    g0127(.A(G223), .ZN(new_n328));
  OAI221_X1 g0128(.A(new_n326), .B1(new_n224), .B2(new_n256), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n263), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(KEYINPUT69), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT69), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n325), .A2(new_n333), .A3(new_n330), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n288), .ZN(new_n336));
  INV_X1    g0136(.A(G169), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n332), .A2(new_n337), .A3(new_n334), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n303), .A2(G50), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n307), .A2(new_n296), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n294), .ZN(new_n342));
  INV_X1    g0142(.A(G58), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(KEYINPUT70), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT70), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(G58), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(KEYINPUT8), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n348), .B1(KEYINPUT8), .B2(G58), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n342), .B1(new_n298), .B2(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n341), .B1(new_n350), .B2(new_n293), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n336), .A2(new_n338), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n332), .A2(G200), .A3(new_n334), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n351), .A2(KEYINPUT9), .ZN(new_n356));
  AND2_X1   g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT74), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(new_n351), .B2(KEYINPUT9), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT9), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n352), .A2(KEYINPUT74), .A3(new_n360), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n335), .A2(G190), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT10), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n357), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  AND3_X1   g0164(.A1(new_n325), .A2(new_n333), .A3(new_n330), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n333), .B1(new_n325), .B2(new_n330), .ZN(new_n366));
  OAI21_X1  g0166(.A(G190), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n361), .A2(new_n359), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n367), .A2(new_n355), .A3(new_n368), .A4(new_n356), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT10), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n354), .B1(new_n364), .B2(new_n370), .ZN(new_n371));
  XNOR2_X1  g0171(.A(KEYINPUT70), .B(G58), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n206), .B1(new_n372), .B2(new_n302), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n373), .A2(G20), .B1(G159), .B2(new_n294), .ZN(new_n374));
  XNOR2_X1  g0174(.A(KEYINPUT77), .B(G33), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n210), .B(new_n254), .C1(new_n375), .C2(new_n252), .ZN(new_n376));
  OAI21_X1  g0176(.A(G68), .B1(new_n376), .B2(KEYINPUT7), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT7), .ZN(new_n378));
  NOR2_X1   g0178(.A1(KEYINPUT3), .A2(G33), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n253), .A2(KEYINPUT77), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT77), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(G33), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n379), .B1(new_n383), .B2(KEYINPUT3), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n378), .B1(new_n384), .B2(new_n210), .ZN(new_n385));
  OAI211_X1 g0185(.A(KEYINPUT16), .B(new_n374), .C1(new_n377), .C2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT16), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n202), .B1(new_n347), .B2(G68), .ZN(new_n388));
  INV_X1    g0188(.A(G159), .ZN(new_n389));
  OAI22_X1  g0189(.A1(new_n388), .A2(new_n210), .B1(new_n389), .B2(new_n295), .ZN(new_n390));
  AND3_X1   g0190(.A1(new_n255), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(new_n383), .B2(KEYINPUT3), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n255), .A2(new_n210), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n378), .B1(new_n393), .B2(new_n379), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n302), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n387), .B1(new_n390), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n386), .A2(new_n293), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n349), .A2(new_n306), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n398), .B1(new_n303), .B2(new_n349), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT78), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n269), .A2(G232), .A3(new_n272), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n401), .B1(new_n270), .B2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n270), .A2(new_n402), .A3(new_n401), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n328), .A2(new_n259), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n261), .A2(G1698), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n252), .B1(new_n380), .B2(new_n382), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n407), .B(new_n408), .C1(new_n409), .C2(new_n379), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G33), .A2(G87), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n269), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(G169), .B1(new_n406), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n410), .A2(new_n411), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n263), .ZN(new_n415));
  AND3_X1   g0215(.A1(new_n270), .A2(new_n402), .A3(new_n401), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n416), .A2(new_n403), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n415), .A2(new_n417), .A3(G179), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n413), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n400), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(KEYINPUT18), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT18), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n400), .A2(new_n422), .A3(new_n419), .ZN(new_n423));
  INV_X1    g0223(.A(G200), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n424), .B1(new_n406), .B2(new_n412), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n415), .A2(new_n417), .A3(new_n314), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n427), .A2(new_n397), .A3(new_n399), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT17), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n427), .A2(new_n397), .A3(KEYINPUT17), .A4(new_n399), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n421), .A2(new_n423), .A3(new_n430), .A4(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  XOR2_X1   g0233(.A(KEYINPUT8), .B(G58), .Z(new_n434));
  AOI22_X1  g0234(.A1(new_n434), .A2(new_n294), .B1(G20), .B2(G77), .ZN(new_n435));
  XNOR2_X1  g0235(.A(KEYINPUT15), .B(G87), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n435), .B1(new_n436), .B2(new_n298), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n293), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n306), .A2(G77), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n439), .B1(new_n303), .B2(G77), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  OR2_X1    g0241(.A1(new_n441), .A2(KEYINPUT71), .ZN(new_n442));
  INV_X1    g0242(.A(new_n255), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n443), .A2(new_n379), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(G107), .ZN(new_n445));
  OAI221_X1 g0245(.A(new_n445), .B1(new_n260), .B2(new_n236), .C1(new_n271), .C2(new_n327), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n263), .ZN(new_n447));
  INV_X1    g0247(.A(G274), .ZN(new_n448));
  AND2_X1   g0248(.A1(G1), .A2(G13), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n448), .B1(new_n449), .B2(new_n268), .ZN(new_n450));
  AOI22_X1  g0250(.A1(new_n321), .A2(G244), .B1(new_n450), .B2(new_n267), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n447), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(G200), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n441), .A2(KEYINPUT71), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n442), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(KEYINPUT72), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT72), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n442), .A2(new_n457), .A3(new_n453), .A4(new_n454), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n456), .B(new_n458), .C1(new_n314), .C2(new_n452), .ZN(new_n459));
  INV_X1    g0259(.A(new_n441), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n460), .B1(new_n452), .B2(new_n337), .ZN(new_n461));
  OR2_X1    g0261(.A1(new_n461), .A2(KEYINPUT73), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n447), .A2(new_n288), .A3(new_n451), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n461), .A2(KEYINPUT73), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  AND2_X1   g0265(.A1(new_n459), .A2(new_n465), .ZN(new_n466));
  AND4_X1   g0266(.A1(new_n320), .A2(new_n371), .A3(new_n433), .A4(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT22), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n210), .A2(G87), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n468), .B1(new_n444), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n383), .A2(new_n210), .A3(G116), .ZN(new_n471));
  OAI21_X1  g0271(.A(KEYINPUT23), .B1(new_n210), .B2(G107), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT23), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n473), .A2(new_n226), .A3(G20), .ZN(new_n474));
  NAND2_X1  g0274(.A1(KEYINPUT87), .A2(KEYINPUT24), .ZN(new_n475));
  AND3_X1   g0275(.A1(new_n472), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n470), .A2(new_n471), .A3(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(KEYINPUT87), .A2(KEYINPUT24), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n254), .B1(new_n375), .B2(new_n252), .ZN(new_n479));
  INV_X1    g0279(.A(G87), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n468), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n479), .A2(new_n210), .A3(new_n481), .ZN(new_n482));
  AND3_X1   g0282(.A1(new_n477), .A2(new_n478), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n478), .B1(new_n477), .B2(new_n482), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n293), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n307), .A2(KEYINPUT25), .A3(new_n226), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(KEYINPUT25), .B1(new_n307), .B2(new_n226), .ZN(new_n488));
  INV_X1    g0288(.A(new_n293), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n213), .A2(G33), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n489), .A2(new_n306), .A3(new_n490), .ZN(new_n491));
  OAI22_X1  g0291(.A1(new_n487), .A2(new_n488), .B1(new_n491), .B2(new_n226), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n485), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n213), .A2(G45), .ZN(new_n495));
  OR2_X1    g0295(.A1(KEYINPUT5), .A2(G41), .ZN(new_n496));
  NAND2_X1  g0296(.A1(KEYINPUT5), .A2(G41), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n450), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n498), .A2(new_n263), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(G264), .ZN(new_n501));
  INV_X1    g0301(.A(G294), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n375), .A2(new_n502), .ZN(new_n503));
  MUX2_X1   g0303(.A(G250), .B(G257), .S(G1698), .Z(new_n504));
  AOI21_X1  g0304(.A(new_n503), .B1(new_n479), .B2(new_n504), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n499), .B(new_n501), .C1(new_n505), .C2(new_n269), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n506), .A2(G179), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n507), .B1(new_n337), .B2(new_n506), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n494), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n506), .A2(new_n424), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n510), .B1(G190), .B2(new_n506), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n511), .A2(new_n485), .A3(new_n493), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(G257), .A2(G1698), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n514), .B1(new_n227), .B2(G1698), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n515), .B1(new_n409), .B2(new_n379), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n444), .A2(G303), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n269), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n266), .A2(G1), .ZN(new_n519));
  INV_X1    g0319(.A(new_n497), .ZN(new_n520));
  NOR2_X1   g0320(.A1(KEYINPUT5), .A2(G41), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n522), .A2(G270), .A3(new_n269), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n499), .ZN(new_n524));
  OAI21_X1  g0324(.A(G200), .B1(new_n518), .B2(new_n524), .ZN(new_n525));
  AND2_X1   g0325(.A1(new_n523), .A2(new_n499), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n479), .A2(new_n515), .B1(G303), .B2(new_n444), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n526), .B(G190), .C1(new_n527), .C2(new_n269), .ZN(new_n528));
  INV_X1    g0328(.A(G116), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n307), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n489), .A2(G116), .A3(new_n306), .A4(new_n490), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n292), .A2(new_n209), .B1(G20), .B2(new_n529), .ZN(new_n532));
  NAND2_X1  g0332(.A1(G33), .A2(G283), .ZN(new_n533));
  INV_X1    g0333(.A(G97), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n533), .B(new_n210), .C1(G33), .C2(new_n534), .ZN(new_n535));
  AND3_X1   g0335(.A1(new_n532), .A2(KEYINPUT20), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(KEYINPUT20), .B1(new_n532), .B2(new_n535), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n530), .B(new_n531), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n525), .A2(new_n528), .A3(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT85), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n525), .A2(new_n528), .A3(KEYINPUT85), .A4(new_n539), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT21), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n538), .A2(G169), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n516), .A2(new_n517), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n524), .B1(new_n547), .B2(new_n263), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n545), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  NOR3_X1   g0349(.A1(new_n518), .A2(new_n288), .A3(new_n524), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n538), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n526), .B1(new_n527), .B2(new_n269), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n552), .A2(KEYINPUT21), .A3(G169), .A4(new_n538), .ZN(new_n553));
  AND3_X1   g0353(.A1(new_n549), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n544), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(KEYINPUT86), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT86), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n544), .A2(new_n557), .A3(new_n554), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n513), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT79), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT4), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n259), .A2(G244), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n561), .B1(new_n384), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n561), .A2(new_n225), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n564), .B(new_n259), .C1(new_n443), .C2(new_n379), .ZN(new_n565));
  OAI211_X1 g0365(.A(G250), .B(G1698), .C1(new_n443), .C2(new_n379), .ZN(new_n566));
  AND3_X1   g0366(.A1(new_n565), .A2(new_n566), .A3(new_n533), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n269), .B1(new_n563), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n500), .A2(G257), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n499), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n560), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n225), .A2(G1698), .ZN(new_n572));
  AOI21_X1  g0372(.A(KEYINPUT4), .B1(new_n479), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n565), .A2(new_n566), .A3(new_n533), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n263), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n500), .A2(G257), .B1(new_n498), .B2(new_n450), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n575), .A2(KEYINPUT79), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(G169), .B1(new_n571), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n294), .A2(G77), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT6), .ZN(new_n580));
  NOR3_X1   g0380(.A1(new_n580), .A2(new_n534), .A3(G107), .ZN(new_n581));
  XNOR2_X1  g0381(.A(G97), .B(G107), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n581), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n579), .B1(new_n583), .B2(new_n210), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n226), .B1(new_n392), .B2(new_n394), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n293), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n306), .A2(G97), .ZN(new_n587));
  INV_X1    g0387(.A(new_n491), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n587), .B1(new_n588), .B2(G97), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n575), .A2(new_n288), .A3(new_n576), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(KEYINPUT80), .B1(new_n578), .B2(new_n592), .ZN(new_n593));
  NOR3_X1   g0393(.A1(new_n568), .A2(new_n560), .A3(new_n570), .ZN(new_n594));
  AOI21_X1  g0394(.A(KEYINPUT79), .B1(new_n575), .B2(new_n576), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n337), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n592), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT80), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n571), .A2(G190), .A3(new_n577), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n424), .B1(new_n575), .B2(new_n576), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n601), .A2(new_n590), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n593), .A2(new_n599), .A3(new_n603), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n210), .B(G68), .C1(new_n409), .C2(new_n379), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT19), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n210), .B1(new_n258), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(G87), .A2(G97), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n608), .A2(KEYINPUT82), .A3(new_n226), .ZN(new_n609));
  AOI21_X1  g0409(.A(KEYINPUT82), .B1(new_n608), .B2(new_n226), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n607), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n606), .B1(new_n298), .B2(new_n534), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n605), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT83), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n605), .A2(KEYINPUT83), .A3(new_n611), .A4(new_n612), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n615), .A2(new_n293), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n436), .A2(new_n307), .ZN(new_n618));
  INV_X1    g0418(.A(new_n436), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n588), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n617), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT84), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n617), .A2(KEYINPUT84), .A3(new_n618), .A4(new_n620), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n269), .A2(G250), .A3(new_n495), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n269), .A2(G274), .A3(new_n519), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT81), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n450), .A2(KEYINPUT81), .A3(new_n519), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n626), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n375), .A2(new_n529), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n225), .A2(G1698), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n633), .B1(G238), .B2(G1698), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n632), .B1(new_n479), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n631), .B1(new_n636), .B2(new_n269), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(G169), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n638), .B1(new_n288), .B2(new_n637), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n623), .A2(new_n624), .A3(new_n639), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n631), .B(new_n314), .C1(new_n269), .C2(new_n636), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n479), .A2(new_n635), .ZN(new_n642));
  INV_X1    g0442(.A(new_n632), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n269), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n629), .A2(new_n630), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n625), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n641), .B1(new_n647), .B2(G200), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n588), .A2(G87), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n648), .A2(new_n649), .A3(new_n618), .A4(new_n617), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n640), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n604), .A2(new_n651), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n467), .A2(new_n559), .A3(new_n652), .ZN(G372));
  AND2_X1   g0453(.A1(new_n593), .A2(new_n599), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n621), .A2(new_n639), .ZN(new_n655));
  AND4_X1   g0455(.A1(new_n512), .A2(new_n603), .A3(new_n650), .A4(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n654), .A2(new_n656), .A3(KEYINPUT88), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n509), .A2(new_n554), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT88), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n593), .A2(new_n599), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n603), .A2(new_n512), .A3(new_n650), .A4(new_n655), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n659), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n657), .A2(new_n658), .A3(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT89), .ZN(new_n664));
  AND3_X1   g0464(.A1(new_n621), .A2(new_n639), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n664), .B1(new_n621), .B2(new_n639), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n571), .A2(new_n577), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n592), .B1(new_n668), .B2(new_n337), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT26), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n669), .A2(new_n670), .A3(new_n650), .A4(new_n655), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n647), .A2(G179), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n621), .A2(new_n622), .B1(new_n638), .B2(new_n673), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n617), .A2(new_n649), .A3(new_n618), .ZN(new_n675));
  AOI22_X1  g0475(.A1(new_n674), .A2(new_n624), .B1(new_n675), .B2(new_n648), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n660), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n672), .B1(new_n677), .B2(KEYINPUT26), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n663), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n467), .A2(new_n679), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n430), .A2(new_n431), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n465), .A2(new_n319), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n681), .B1(new_n313), .B2(new_n682), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n400), .A2(new_n422), .A3(new_n419), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n422), .B1(new_n400), .B2(new_n419), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n364), .A2(new_n370), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n354), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n680), .A2(new_n689), .ZN(G369));
  NAND2_X1  g0490(.A1(new_n556), .A2(new_n558), .ZN(new_n691));
  INV_X1    g0491(.A(new_n554), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n213), .A2(new_n210), .A3(G13), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(G213), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(G343), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n539), .A2(new_n699), .ZN(new_n700));
  MUX2_X1   g0500(.A(new_n691), .B(new_n692), .S(new_n700), .Z(new_n701));
  NAND2_X1  g0501(.A1(new_n494), .A2(new_n698), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n702), .A2(new_n509), .A3(new_n512), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n494), .A2(new_n508), .A3(new_n698), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n701), .A2(G330), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n692), .A2(new_n699), .ZN(new_n707));
  OAI22_X1  g0507(.A1(new_n703), .A2(new_n707), .B1(new_n509), .B2(new_n698), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n706), .A2(new_n709), .ZN(G399));
  INV_X1    g0510(.A(new_n216), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(G41), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n609), .A2(new_n610), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n529), .ZN(new_n714));
  NOR3_X1   g0514(.A1(new_n712), .A2(new_n213), .A3(new_n714), .ZN(new_n715));
  AOI22_X1  g0515(.A1(new_n715), .A2(KEYINPUT90), .B1(new_n208), .B2(new_n712), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n716), .B1(KEYINPUT90), .B2(new_n715), .ZN(new_n717));
  XOR2_X1   g0517(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n718));
  XNOR2_X1  g0518(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n679), .A2(new_n699), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT29), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n669), .A2(KEYINPUT26), .A3(new_n650), .A4(new_n655), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(KEYINPUT93), .ZN(new_n724));
  AOI22_X1  g0524(.A1(new_n675), .A2(new_n648), .B1(new_n621), .B2(new_n639), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT93), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n725), .A2(new_n726), .A3(KEYINPUT26), .A4(new_n669), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(KEYINPUT26), .B1(new_n676), .B2(new_n660), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n603), .A2(new_n512), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n731), .A2(new_n725), .A3(new_n593), .A4(new_n599), .ZN(new_n732));
  INV_X1    g0532(.A(new_n658), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n667), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  OAI211_X1 g0534(.A(KEYINPUT29), .B(new_n699), .C1(new_n730), .C2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(KEYINPUT94), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n660), .A2(new_n661), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n658), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n738), .B(new_n667), .C1(new_n729), .C2(new_n728), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT94), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n739), .A2(new_n740), .A3(KEYINPUT29), .A4(new_n699), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n722), .A2(new_n736), .A3(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(G330), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n501), .B1(new_n505), .B2(new_n269), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n637), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n571), .A2(new_n745), .A3(new_n550), .A4(new_n577), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT92), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT30), .ZN(new_n748));
  AND3_X1   g0548(.A1(new_n746), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n748), .B1(new_n746), .B2(new_n747), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n506), .B1(new_n568), .B2(new_n570), .ZN(new_n751));
  NOR4_X1   g0551(.A1(new_n751), .A2(new_n647), .A3(G179), .A4(new_n548), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n749), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT31), .ZN(new_n754));
  NOR3_X1   g0554(.A1(new_n753), .A2(new_n754), .A3(new_n699), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n746), .A2(new_n747), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n752), .B1(new_n756), .B2(KEYINPUT30), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n746), .A2(new_n747), .A3(new_n748), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(KEYINPUT31), .B1(new_n759), .B2(new_n698), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n755), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n559), .A2(new_n652), .A3(new_n699), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n743), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n742), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n719), .B1(new_n766), .B2(G1), .ZN(G364));
  INV_X1    g0567(.A(G13), .ZN(new_n768));
  NOR3_X1   g0568(.A1(new_n768), .A2(new_n266), .A3(G20), .ZN(new_n769));
  OR2_X1    g0569(.A1(new_n769), .A2(KEYINPUT95), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(KEYINPUT95), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n770), .A2(G1), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n712), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n773), .B1(new_n701), .B2(G330), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n774), .B1(G330), .B2(new_n701), .ZN(new_n775));
  OAI21_X1  g0575(.A(G20), .B1(KEYINPUT97), .B2(G169), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(KEYINPUT97), .A2(G169), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n209), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G13), .A2(G33), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(G20), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n247), .A2(new_n266), .ZN(new_n785));
  INV_X1    g0585(.A(KEYINPUT96), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n711), .A2(new_n479), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n788), .B1(new_n266), .B2(new_n208), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n785), .B1(new_n786), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n790), .B1(new_n786), .B2(new_n789), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n711), .A2(new_n444), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n792), .A2(G355), .B1(new_n529), .B2(new_n711), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n784), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n779), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n210), .A2(new_n314), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n796), .A2(G179), .A3(new_n424), .ZN(new_n797));
  INV_X1    g0597(.A(G322), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n424), .A2(G179), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(G303), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n797), .A2(new_n798), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n314), .A2(new_n424), .A3(G20), .A4(G179), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n256), .B(new_n802), .C1(G311), .C2(new_n804), .ZN(new_n805));
  NAND4_X1  g0605(.A1(G20), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n806), .A2(KEYINPUT98), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n806), .A2(KEYINPUT98), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(G326), .ZN(new_n811));
  NOR4_X1   g0611(.A1(new_n210), .A2(new_n288), .A3(new_n424), .A4(G190), .ZN(new_n812));
  XNOR2_X1  g0612(.A(KEYINPUT33), .B(G317), .ZN(new_n813));
  NOR2_X1   g0613(.A1(G179), .A2(G200), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n210), .B1(new_n814), .B2(G190), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n812), .A2(new_n813), .B1(new_n816), .B2(G294), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT99), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(new_n210), .B2(G190), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n314), .A2(KEYINPUT99), .A3(G20), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n819), .A2(new_n799), .A3(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n819), .A2(new_n814), .A3(new_n820), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  AOI22_X1  g0624(.A1(G283), .A2(new_n822), .B1(new_n824), .B2(G329), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n805), .A2(new_n811), .A3(new_n817), .A4(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n812), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n827), .A2(new_n302), .B1(new_n815), .B2(new_n534), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n256), .B1(new_n800), .B2(new_n480), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n797), .A2(new_n372), .B1(new_n803), .B2(new_n224), .ZN(new_n830));
  NOR3_X1   g0630(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n823), .A2(new_n389), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n832), .B(KEYINPUT32), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n810), .A2(G50), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n822), .A2(G107), .ZN(new_n835));
  NAND4_X1  g0635(.A1(new_n831), .A2(new_n833), .A3(new_n834), .A4(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n795), .B1(new_n826), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n773), .ZN(new_n838));
  NOR3_X1   g0638(.A1(new_n794), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n782), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n839), .B1(new_n701), .B2(new_n840), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n775), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(G396));
  NOR2_X1   g0643(.A1(new_n460), .A2(new_n699), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n459), .A2(new_n465), .A3(new_n845), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n462), .A2(new_n463), .A3(new_n464), .A4(new_n844), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n720), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n459), .A2(new_n465), .A3(new_n699), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(new_n663), .B2(new_n678), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n848), .A2(new_n763), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n838), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n853), .A2(KEYINPUT101), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n848), .A2(new_n851), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n764), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n853), .A2(KEYINPUT101), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n854), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n797), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n859), .A2(G143), .B1(G159), .B2(new_n804), .ZN(new_n860));
  INV_X1    g0660(.A(G150), .ZN(new_n861));
  INV_X1    g0661(.A(G137), .ZN(new_n862));
  OAI221_X1 g0662(.A(new_n860), .B1(new_n861), .B2(new_n827), .C1(new_n809), .C2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n864), .A2(KEYINPUT34), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n864), .A2(KEYINPUT34), .ZN(new_n866));
  OAI221_X1 g0666(.A(new_n479), .B1(new_n296), .B2(new_n800), .C1(new_n372), .C2(new_n815), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n822), .A2(G68), .ZN(new_n868));
  INV_X1    g0668(.A(G132), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n868), .B1(new_n869), .B2(new_n823), .ZN(new_n870));
  NOR4_X1   g0670(.A1(new_n865), .A2(new_n866), .A3(new_n867), .A4(new_n870), .ZN(new_n871));
  OAI22_X1  g0671(.A1(new_n800), .A2(new_n226), .B1(new_n529), .B2(new_n803), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n256), .B(new_n872), .C1(G294), .C2(new_n859), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n810), .A2(G303), .ZN(new_n874));
  AOI22_X1  g0674(.A1(G283), .A2(new_n812), .B1(new_n816), .B2(G97), .ZN(new_n875));
  AOI22_X1  g0675(.A1(G87), .A2(new_n822), .B1(new_n824), .B2(G311), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n873), .A2(new_n874), .A3(new_n875), .A4(new_n876), .ZN(new_n877));
  XNOR2_X1  g0677(.A(new_n877), .B(KEYINPUT100), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n779), .B1(new_n871), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n779), .A2(new_n780), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n838), .B1(new_n224), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n846), .A2(new_n847), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n879), .B(new_n881), .C1(new_n882), .C2(new_n781), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n858), .A2(new_n883), .ZN(G384));
  INV_X1    g0684(.A(new_n583), .ZN(new_n885));
  OR2_X1    g0685(.A1(new_n885), .A2(KEYINPUT35), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(KEYINPUT35), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n886), .A2(G116), .A3(new_n211), .A4(new_n887), .ZN(new_n888));
  XOR2_X1   g0688(.A(new_n888), .B(KEYINPUT36), .Z(new_n889));
  OAI211_X1 g0689(.A(new_n208), .B(G77), .C1(new_n302), .C2(new_n372), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n201), .A2(G68), .ZN(new_n891));
  AOI211_X1 g0691(.A(new_n213), .B(G13), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT38), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT37), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n397), .A2(new_n399), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n386), .A2(new_n293), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n384), .A2(new_n378), .A3(new_n210), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n376), .A2(KEYINPUT7), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n898), .A2(new_n899), .A3(G68), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT16), .B1(new_n900), .B2(new_n374), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n399), .B1(new_n897), .B2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n696), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n896), .A2(new_n427), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n902), .A2(new_n419), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n895), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n400), .A2(new_n903), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n420), .A2(new_n907), .A3(new_n895), .A4(new_n428), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n902), .A2(new_n903), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n681), .B2(new_n686), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n894), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n905), .A2(new_n911), .A3(new_n428), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(KEYINPUT37), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n908), .ZN(new_n916));
  INV_X1    g0716(.A(new_n911), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n432), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n916), .A2(new_n918), .A3(KEYINPUT38), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n913), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n311), .A2(new_n698), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n312), .A2(new_n318), .A3(new_n921), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n311), .B(new_n698), .C1(new_n291), .C2(new_n319), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n462), .A2(new_n463), .A3(new_n464), .A4(new_n699), .ZN(new_n925));
  XOR2_X1   g0725(.A(new_n925), .B(KEYINPUT102), .Z(new_n926));
  OAI211_X1 g0726(.A(new_n920), .B(new_n924), .C1(new_n850), .C2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n696), .B1(new_n684), .B2(new_n685), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n907), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n432), .A2(KEYINPUT103), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n420), .A2(new_n907), .A3(new_n428), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(KEYINPUT37), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n908), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT103), .B1(new_n432), .B2(new_n931), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n894), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n919), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT39), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n312), .A2(new_n698), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n913), .A2(KEYINPUT39), .A3(new_n919), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n930), .A2(new_n944), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n722), .A2(new_n736), .A3(new_n467), .A4(new_n741), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n689), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n945), .B(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  AND3_X1   g0749(.A1(new_n559), .A2(new_n652), .A3(new_n699), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n754), .B1(new_n753), .B2(new_n699), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n759), .A2(KEYINPUT31), .A3(new_n698), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n882), .B(new_n924), .C1(new_n950), .C2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT104), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT40), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(new_n938), .B2(new_n919), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n762), .A2(new_n951), .A3(new_n952), .ZN(new_n959));
  NAND4_X1  g0759(.A1(new_n959), .A2(KEYINPUT104), .A3(new_n882), .A4(new_n924), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n956), .A2(new_n958), .A3(new_n960), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n920), .A2(new_n959), .A3(new_n882), .A4(new_n924), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n957), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n467), .A2(new_n959), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n964), .A2(new_n965), .ZN(new_n967));
  NOR3_X1   g0767(.A1(new_n966), .A2(new_n967), .A3(new_n743), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n949), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(G1), .B1(new_n768), .B2(G20), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n949), .B2(new_n968), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n893), .B1(new_n969), .B2(new_n971), .ZN(G367));
  NOR2_X1   g0772(.A1(new_n788), .A2(new_n242), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n783), .B1(new_n216), .B2(new_n436), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n797), .A2(new_n861), .B1(new_n201), .B2(new_n803), .ZN(new_n975));
  INV_X1    g0775(.A(new_n800), .ZN(new_n976));
  AOI211_X1 g0776(.A(new_n444), .B(new_n975), .C1(new_n347), .C2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n810), .A2(G143), .ZN(new_n978));
  AOI22_X1  g0778(.A1(G159), .A2(new_n812), .B1(new_n816), .B2(G68), .ZN(new_n979));
  AOI22_X1  g0779(.A1(G77), .A2(new_n822), .B1(new_n824), .B2(G137), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n977), .A2(new_n978), .A3(new_n979), .A4(new_n980), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n859), .A2(G303), .B1(G283), .B2(new_n804), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n502), .B2(new_n827), .ZN(new_n983));
  OAI21_X1  g0783(.A(KEYINPUT105), .B1(new_n800), .B2(new_n529), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT46), .ZN(new_n985));
  AOI211_X1 g0785(.A(new_n983), .B(new_n985), .C1(G107), .C2(new_n816), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n810), .A2(G311), .ZN(new_n987));
  INV_X1    g0787(.A(G317), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n384), .B1(new_n821), .B2(new_n534), .C1(new_n988), .C2(new_n823), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n986), .B(new_n987), .C1(KEYINPUT106), .C2(new_n989), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n989), .A2(KEYINPUT106), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n981), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n992), .B(KEYINPUT47), .Z(new_n993));
  OAI221_X1 g0793(.A(new_n773), .B1(new_n973), .B2(new_n974), .C1(new_n993), .C2(new_n795), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT107), .Z(new_n995));
  OR2_X1    g0795(.A1(new_n675), .A2(new_n699), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n667), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(new_n725), .B2(new_n996), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n782), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n995), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n590), .A2(new_n698), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n654), .A2(new_n603), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n669), .A2(new_n698), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n708), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT44), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1004), .B(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n709), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT45), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1007), .A2(new_n709), .A3(KEYINPUT45), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1006), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n706), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1006), .A2(new_n1012), .A3(new_n706), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n701), .A2(G330), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n703), .A2(new_n707), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n705), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1019), .B1(new_n1020), .B2(new_n707), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1018), .B(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n766), .B1(new_n1017), .B2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n712), .B(KEYINPUT41), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n772), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1007), .A2(new_n1019), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT42), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1027), .B(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n509), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n699), .B1(new_n1030), .B2(new_n660), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT43), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n998), .A2(new_n1033), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n998), .A2(new_n1033), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1032), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1029), .A2(new_n1033), .A3(new_n998), .A4(new_n1031), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n706), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1036), .A2(new_n1039), .A3(new_n1037), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1000), .B1(new_n1026), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT108), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  OAI211_X1 g0846(.A(KEYINPUT108), .B(new_n1000), .C1(new_n1026), .C2(new_n1043), .ZN(new_n1047));
  AND2_X1   g0847(.A1(new_n1046), .A2(new_n1047), .ZN(G387));
  NAND2_X1  g0848(.A1(new_n765), .A2(new_n1023), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n742), .A2(new_n1022), .A3(new_n764), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1049), .A2(new_n712), .A3(new_n1050), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n797), .A2(new_n988), .B1(new_n803), .B2(new_n801), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(G311), .B2(new_n812), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n798), .B2(new_n809), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT48), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n976), .A2(G294), .B1(new_n816), .B2(G283), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT49), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n821), .A2(new_n529), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n479), .B(new_n1063), .C1(G326), .C2(new_n824), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1061), .A2(new_n1062), .A3(new_n1064), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n800), .A2(new_n224), .B1(new_n302), .B2(new_n803), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n816), .A2(new_n619), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n479), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n1066), .B(new_n1068), .C1(G50), .C2(new_n859), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n349), .A2(new_n827), .B1(new_n534), .B2(new_n821), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(G150), .B2(new_n824), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1069), .B(new_n1071), .C1(new_n389), .C2(new_n809), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n795), .B1(new_n1065), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT111), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n792), .A2(new_n714), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1075), .B1(G107), .B2(new_n216), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n239), .A2(G45), .ZN(new_n1077));
  XOR2_X1   g0877(.A(new_n1077), .B(KEYINPUT109), .Z(new_n1078));
  NAND2_X1  g0878(.A1(new_n434), .A2(new_n296), .ZN(new_n1079));
  XOR2_X1   g0879(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n1080));
  AND2_X1   g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n266), .B1(new_n302), .B2(new_n224), .ZN(new_n1083));
  NOR3_X1   g0883(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n714), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n788), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1076), .B1(new_n1078), .B2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n773), .B1(new_n1087), .B2(new_n784), .ZN(new_n1088));
  OR3_X1    g0888(.A1(new_n1073), .A2(new_n1074), .A3(new_n1088), .ZN(new_n1089));
  OR2_X1    g0889(.A1(new_n1073), .A2(new_n1088), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n1090), .A2(new_n1074), .B1(new_n1020), .B2(new_n782), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n1022), .A2(new_n772), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1051), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT112), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1051), .A2(KEYINPUT112), .A3(new_n1092), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1095), .A2(new_n1096), .ZN(G393));
  INV_X1    g0897(.A(KEYINPUT113), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1016), .A2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n706), .B1(new_n1006), .B2(new_n1012), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1015), .A2(new_n1098), .A3(new_n1016), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n772), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n783), .B1(new_n534), .B2(new_n216), .C1(new_n788), .C2(new_n250), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n773), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n810), .A2(G317), .B1(G311), .B2(new_n859), .ZN(new_n1107));
  XOR2_X1   g0907(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n444), .B1(new_n803), .B2(new_n502), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n827), .A2(new_n801), .B1(new_n815), .B2(new_n529), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n1110), .B(new_n1111), .C1(G283), .C2(new_n976), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n824), .A2(G322), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1109), .A2(new_n835), .A3(new_n1112), .A4(new_n1113), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n809), .A2(new_n861), .B1(new_n389), .B2(new_n797), .ZN(new_n1116));
  XOR2_X1   g0916(.A(new_n1116), .B(KEYINPUT51), .Z(new_n1117));
  AOI22_X1  g0917(.A1(G87), .A2(new_n822), .B1(new_n824), .B2(G143), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n976), .A2(G68), .B1(new_n434), .B2(new_n804), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n201), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n1120), .A2(new_n812), .B1(new_n816), .B2(G77), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1118), .A2(new_n479), .A3(new_n1119), .A4(new_n1121), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n1114), .A2(new_n1115), .B1(new_n1117), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1106), .B1(new_n1123), .B2(new_n779), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n1007), .B2(new_n840), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1050), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1103), .A2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n712), .B1(new_n1017), .B2(new_n1050), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1104), .B(new_n1125), .C1(new_n1127), .C2(new_n1128), .ZN(G390));
  NAND4_X1  g0929(.A1(new_n959), .A2(G330), .A3(new_n882), .A4(new_n924), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n924), .B1(new_n850), .B2(new_n926), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n942), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n941), .A2(new_n943), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n924), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n882), .B(new_n699), .C1(new_n730), .C2(new_n734), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1135), .B1(new_n1136), .B2(new_n925), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n939), .A2(new_n1133), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1131), .B1(new_n1134), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n467), .A2(new_n763), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n946), .A2(new_n689), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n924), .B1(new_n763), .B2(new_n882), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n1143), .A2(new_n1131), .B1(new_n850), .B2(new_n926), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n959), .A2(G330), .A3(new_n882), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n1135), .ZN(new_n1146));
  AND2_X1   g0946(.A1(new_n1136), .A2(new_n925), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1146), .A2(new_n1147), .A3(new_n1130), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1144), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1150));
  AND3_X1   g0950(.A1(new_n916), .A2(new_n918), .A3(KEYINPUT38), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n432), .A2(new_n931), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT103), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1154), .A2(new_n935), .A3(new_n932), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1151), .B1(new_n1155), .B2(new_n894), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n943), .B1(new_n1156), .B2(KEYINPUT39), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1150), .A2(new_n1157), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1156), .A2(new_n942), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1159), .B1(new_n1147), .B2(new_n1135), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1158), .A2(new_n1160), .A3(new_n1130), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1140), .A2(new_n1142), .A3(new_n1149), .A4(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n712), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT115), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1149), .A2(new_n1142), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1130), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1167));
  NOR3_X1   g0967(.A1(new_n1134), .A2(new_n1139), .A3(new_n1131), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1166), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1162), .A2(KEYINPUT115), .A3(new_n712), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1165), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1168), .A2(new_n1167), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(new_n772), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n838), .B1(new_n349), .B2(new_n880), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n868), .B1(new_n224), .B2(new_n815), .C1(new_n529), .C2(new_n797), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(G283), .B2(new_n810), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n812), .A2(G107), .B1(new_n804), .B2(G97), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT116), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n444), .B1(new_n800), .B2(new_n480), .ZN(new_n1179));
  OR2_X1    g0979(.A1(new_n1179), .A2(KEYINPUT117), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n1179), .A2(KEYINPUT117), .B1(new_n824), .B2(G294), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1176), .A2(new_n1178), .A3(new_n1180), .A4(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(KEYINPUT54), .B(G143), .ZN(new_n1183));
  OAI221_X1 g0983(.A(new_n256), .B1(new_n1183), .B2(new_n803), .C1(new_n797), .C2(new_n869), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n827), .A2(new_n862), .B1(new_n815), .B2(new_n389), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n1184), .B(new_n1185), .C1(new_n810), .C2(G128), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n824), .A2(G125), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n976), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT53), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n800), .B2(new_n861), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n1188), .A2(new_n1190), .B1(new_n1120), .B2(new_n822), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1186), .A2(new_n1187), .A3(new_n1191), .ZN(new_n1192));
  AND2_X1   g0992(.A1(new_n1182), .A2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1174), .B1(new_n1193), .B2(new_n795), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(new_n1157), .B2(new_n780), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1195), .B(KEYINPUT118), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1173), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1171), .A2(new_n1198), .ZN(G378));
  AOI21_X1  g0999(.A(new_n363), .B1(new_n357), .B2(new_n362), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n369), .A2(KEYINPUT10), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n353), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n351), .A2(new_n696), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n688), .B(new_n353), .C1(new_n351), .C2(new_n696), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1206));
  AND3_X1   g1006(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1206), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n743), .B1(new_n962), .B2(new_n957), .ZN(new_n1210));
  AND3_X1   g1010(.A1(new_n961), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1209), .B1(new_n961), .B2(new_n1210), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1157), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n929), .B1(new_n1213), .B2(new_n942), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT121), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n1211), .A2(new_n1212), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n961), .A2(new_n1210), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1209), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1215), .B1(new_n930), .B2(new_n944), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n961), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1219), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1216), .A2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1209), .A2(new_n780), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n880), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n773), .B1(new_n1225), .B2(new_n1120), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n409), .A2(G33), .ZN(new_n1227));
  AOI21_X1  g1027(.A(G50), .B1(new_n1227), .B2(new_n265), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n384), .B1(new_n302), .B2(new_n815), .C1(new_n827), .C2(new_n534), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(new_n810), .B2(G116), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n265), .B1(new_n436), .B2(new_n803), .C1(new_n800), .C2(new_n224), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(G283), .B2(new_n824), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n821), .A2(new_n372), .ZN(new_n1233));
  OR3_X1    g1033(.A1(new_n797), .A2(KEYINPUT119), .A3(new_n226), .ZN(new_n1234));
  OAI21_X1  g1034(.A(KEYINPUT119), .B1(new_n797), .B2(new_n226), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1233), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1230), .A2(new_n1232), .A3(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT58), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1228), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n824), .A2(G124), .ZN(new_n1240));
  AOI211_X1 g1040(.A(G33), .B(G41), .C1(new_n822), .C2(G159), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1183), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n976), .A2(new_n1242), .B1(G137), .B2(new_n804), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n859), .A2(G128), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1243), .B(new_n1244), .C1(new_n869), .C2(new_n827), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n810), .A2(G125), .B1(G150), .B2(new_n816), .ZN(new_n1246));
  OR2_X1    g1046(.A1(new_n1246), .A2(KEYINPUT120), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(KEYINPUT120), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1245), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT59), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1240), .B(new_n1241), .C1(new_n1249), .C2(new_n1250), .ZN(new_n1251));
  AND2_X1   g1051(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1252));
  OAI221_X1 g1052(.A(new_n1239), .B1(new_n1238), .B2(new_n1237), .C1(new_n1251), .C2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1226), .B1(new_n1253), .B2(new_n779), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n1223), .A2(new_n772), .B1(new_n1224), .B2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n946), .A2(new_n689), .A3(new_n1141), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(new_n1172), .B2(new_n1149), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n945), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1219), .A2(new_n1214), .A3(new_n1221), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1258), .A2(new_n1259), .A3(KEYINPUT57), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n712), .B1(new_n1257), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1162), .A2(new_n1142), .ZN(new_n1262));
  AOI21_X1  g1062(.A(KEYINPUT57), .B1(new_n1223), .B2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1255), .B1(new_n1261), .B2(new_n1263), .ZN(G375));
  INV_X1    g1064(.A(new_n772), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(new_n1144), .B2(new_n1148), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1135), .A2(new_n780), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n773), .B1(new_n1225), .B2(G68), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n827), .A2(new_n529), .B1(new_n803), .B2(new_n226), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT122), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(new_n1269), .A2(new_n1270), .B1(G294), .B2(new_n810), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1271), .B1(new_n1270), .B2(new_n1269), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(G77), .A2(new_n822), .B1(new_n824), .B2(G303), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n976), .A2(G97), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n256), .B1(new_n859), .B2(G283), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1273), .A2(new_n1067), .A3(new_n1274), .A4(new_n1275), .ZN(new_n1276));
  AOI22_X1  g1076(.A1(new_n859), .A2(G137), .B1(new_n976), .B2(G159), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1233), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n824), .A2(G128), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n804), .A2(G150), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1277), .A2(new_n1278), .A3(new_n1279), .A4(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n384), .B1(new_n812), .B2(new_n1242), .ZN(new_n1282));
  OAI221_X1 g1082(.A(new_n1282), .B1(new_n296), .B2(new_n815), .C1(new_n809), .C2(new_n869), .ZN(new_n1283));
  OAI22_X1  g1083(.A1(new_n1272), .A2(new_n1276), .B1(new_n1281), .B2(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1268), .B1(new_n1284), .B2(new_n779), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1267), .A2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(KEYINPUT123), .B1(new_n1266), .B2(new_n1287), .ZN(new_n1288));
  AND3_X1   g1088(.A1(new_n1146), .A2(new_n1147), .A3(new_n1130), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n850), .A2(new_n926), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1290), .B1(new_n1146), .B2(new_n1130), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n772), .B1(new_n1289), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT123), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1292), .A2(new_n1293), .A3(new_n1286), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1288), .A2(new_n1294), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1149), .A2(new_n1142), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1166), .A2(new_n1025), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1295), .B1(new_n1296), .B2(new_n1297), .ZN(G381));
  NAND3_X1  g1098(.A1(new_n1095), .A2(new_n842), .A3(new_n1096), .ZN(new_n1299));
  OR4_X1    g1099(.A1(G384), .A2(new_n1299), .A3(G381), .A4(G390), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1223), .A2(new_n772), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1224), .A2(new_n1254), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n712), .ZN(new_n1304));
  AND3_X1   g1104(.A1(new_n1258), .A2(new_n1259), .A3(KEYINPUT57), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1304), .B1(new_n1305), .B2(new_n1262), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1223), .A2(new_n1262), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT57), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1303), .B1(new_n1306), .B2(new_n1309), .ZN(new_n1310));
  AND2_X1   g1110(.A1(new_n1170), .A2(new_n1169), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1197), .B1(new_n1311), .B2(new_n1165), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1310), .A2(new_n1312), .ZN(new_n1313));
  OR3_X1    g1113(.A1(new_n1300), .A2(new_n1313), .A3(G387), .ZN(G407));
  OAI211_X1 g1114(.A(G407), .B(G213), .C1(G343), .C2(new_n1313), .ZN(G409));
  NAND2_X1  g1115(.A1(new_n697), .A2(G213), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1223), .A2(new_n1262), .A3(new_n1025), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1258), .A2(new_n1259), .A3(new_n772), .ZN(new_n1318));
  AND2_X1   g1118(.A1(new_n1318), .A2(new_n1302), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1171), .A2(new_n1198), .A3(new_n1317), .A4(new_n1319), .ZN(new_n1320));
  OAI211_X1 g1120(.A(new_n1316), .B(new_n1320), .C1(new_n1310), .C2(new_n1312), .ZN(new_n1321));
  AND2_X1   g1121(.A1(new_n858), .A2(new_n883), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1256), .A2(KEYINPUT60), .A3(new_n1144), .A4(new_n1148), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(new_n712), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1296), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(new_n1289), .A2(new_n1291), .ZN(new_n1326));
  OAI21_X1  g1126(.A(KEYINPUT60), .B1(new_n1326), .B2(new_n1256), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1324), .B1(new_n1325), .B2(new_n1327), .ZN(new_n1328));
  NOR3_X1   g1128(.A1(new_n1266), .A2(KEYINPUT123), .A3(new_n1287), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1293), .B1(new_n1292), .B2(new_n1286), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1322), .B1(new_n1328), .B2(new_n1331), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1296), .B1(KEYINPUT60), .B2(new_n1166), .ZN(new_n1333));
  OAI211_X1 g1133(.A(G384), .B(new_n1295), .C1(new_n1333), .C2(new_n1324), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n697), .A2(G213), .A3(G2897), .ZN(new_n1335));
  AND3_X1   g1135(.A1(new_n1332), .A2(new_n1334), .A3(new_n1335), .ZN(new_n1336));
  AOI21_X1  g1136(.A(new_n1335), .B1(new_n1332), .B2(new_n1334), .ZN(new_n1337));
  NOR2_X1   g1137(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1338));
  AOI21_X1  g1138(.A(KEYINPUT61), .B1(new_n1321), .B2(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(G375), .A2(G378), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1332), .A2(new_n1334), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1341), .ZN(new_n1342));
  NAND4_X1  g1142(.A1(new_n1340), .A2(new_n1316), .A3(new_n1342), .A4(new_n1320), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1343), .A2(KEYINPUT62), .ZN(new_n1344));
  AOI22_X1  g1144(.A1(G375), .A2(G378), .B1(G213), .B2(new_n697), .ZN(new_n1345));
  INV_X1    g1145(.A(KEYINPUT62), .ZN(new_n1346));
  NAND4_X1  g1146(.A1(new_n1345), .A2(new_n1346), .A3(new_n1342), .A4(new_n1320), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1339), .A2(new_n1344), .A3(new_n1347), .ZN(new_n1348));
  INV_X1    g1148(.A(G390), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1349), .A2(new_n1044), .ZN(new_n1350));
  OAI211_X1 g1150(.A(G390), .B(new_n1000), .C1(new_n1026), .C2(new_n1043), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1350), .A2(new_n1351), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(G393), .A2(G396), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1353), .A2(KEYINPUT125), .A3(new_n1299), .ZN(new_n1354));
  INV_X1    g1154(.A(KEYINPUT125), .ZN(new_n1355));
  INV_X1    g1155(.A(new_n1096), .ZN(new_n1356));
  AOI21_X1  g1156(.A(KEYINPUT112), .B1(new_n1051), .B2(new_n1092), .ZN(new_n1357));
  NOR3_X1   g1157(.A1(new_n1356), .A2(G396), .A3(new_n1357), .ZN(new_n1358));
  AOI21_X1  g1158(.A(new_n842), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1359));
  OAI21_X1  g1159(.A(new_n1355), .B1(new_n1358), .B2(new_n1359), .ZN(new_n1360));
  NAND3_X1  g1160(.A1(new_n1352), .A2(new_n1354), .A3(new_n1360), .ZN(new_n1361));
  NAND3_X1  g1161(.A1(new_n1046), .A2(new_n1047), .A3(new_n1349), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1353), .A2(new_n1299), .ZN(new_n1363));
  NAND3_X1  g1163(.A1(new_n1362), .A2(new_n1363), .A3(new_n1351), .ZN(new_n1364));
  AND3_X1   g1164(.A1(new_n1361), .A2(KEYINPUT126), .A3(new_n1364), .ZN(new_n1365));
  AOI21_X1  g1165(.A(KEYINPUT126), .B1(new_n1361), .B2(new_n1364), .ZN(new_n1366));
  NOR2_X1   g1166(.A1(new_n1365), .A2(new_n1366), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1348), .A2(new_n1367), .ZN(new_n1368));
  XOR2_X1   g1168(.A(KEYINPUT124), .B(KEYINPUT63), .Z(new_n1369));
  NAND2_X1  g1169(.A1(new_n1343), .A2(new_n1369), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1361), .A2(new_n1364), .ZN(new_n1371));
  NAND4_X1  g1171(.A1(new_n1345), .A2(KEYINPUT63), .A3(new_n1342), .A4(new_n1320), .ZN(new_n1372));
  NAND4_X1  g1172(.A1(new_n1339), .A2(new_n1370), .A3(new_n1371), .A4(new_n1372), .ZN(new_n1373));
  NAND2_X1  g1173(.A1(new_n1368), .A2(new_n1373), .ZN(G405));
  NAND2_X1  g1174(.A1(new_n1313), .A2(new_n1340), .ZN(new_n1375));
  NOR2_X1   g1175(.A1(new_n1341), .A2(KEYINPUT127), .ZN(new_n1376));
  NAND2_X1  g1176(.A1(new_n1375), .A2(new_n1376), .ZN(new_n1377));
  OAI211_X1 g1177(.A(new_n1313), .B(new_n1340), .C1(KEYINPUT127), .C2(new_n1341), .ZN(new_n1378));
  NAND2_X1  g1178(.A1(new_n1377), .A2(new_n1378), .ZN(new_n1379));
  OAI21_X1  g1179(.A(new_n1379), .B1(new_n1366), .B2(new_n1365), .ZN(new_n1380));
  INV_X1    g1180(.A(new_n1366), .ZN(new_n1381));
  NAND3_X1  g1181(.A1(new_n1361), .A2(KEYINPUT126), .A3(new_n1364), .ZN(new_n1382));
  NAND4_X1  g1182(.A1(new_n1381), .A2(new_n1377), .A3(new_n1382), .A4(new_n1378), .ZN(new_n1383));
  NAND2_X1  g1183(.A1(new_n1380), .A2(new_n1383), .ZN(G402));
endmodule


