//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 0 1 1 1 1 1 0 1 1 0 0 1 1 0 0 0 0 1 0 0 0 0 0 0 1 1 0 1 0 1 1 1 1 1 1 0 0 1 0 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:19 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n782, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n991, new_n992,
    new_n993, new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054;
  INV_X1    g000(.A(KEYINPUT11), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G137), .ZN(new_n189));
  INV_X1    g003(.A(G137), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT11), .A3(G134), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n188), .A2(G137), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G131), .ZN(new_n194));
  AND2_X1   g008(.A1(KEYINPUT65), .A2(G131), .ZN(new_n195));
  NOR2_X1   g009(.A1(KEYINPUT65), .A2(G131), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n197), .A2(new_n189), .A3(new_n191), .A4(new_n192), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n194), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT68), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n202), .A2(G143), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  XNOR2_X1  g018(.A(KEYINPUT64), .B(G143), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n204), .B1(new_n205), .B2(G146), .ZN(new_n206));
  AND2_X1   g020(.A1(KEYINPUT0), .A2(G128), .ZN(new_n207));
  NOR2_X1   g021(.A1(KEYINPUT0), .A2(G128), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n202), .A2(G143), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n211), .B1(new_n205), .B2(G146), .ZN(new_n212));
  AOI22_X1  g026(.A1(new_n206), .A2(new_n209), .B1(new_n212), .B2(new_n207), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n194), .A2(new_n198), .A3(KEYINPUT68), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n201), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G143), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT64), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT64), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G143), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n217), .A2(new_n219), .A3(G146), .ZN(new_n220));
  INV_X1    g034(.A(G128), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n220), .A2(new_n210), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n217), .A2(new_n219), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n203), .B1(new_n224), .B2(new_n202), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n221), .B1(new_n210), .B2(KEYINPUT1), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n223), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n189), .A2(new_n191), .A3(new_n192), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n229), .B1(new_n188), .B2(G137), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n190), .A2(KEYINPUT66), .A3(G134), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n230), .A2(new_n192), .A3(new_n231), .ZN(new_n232));
  AOI22_X1  g046(.A1(new_n228), .A2(new_n197), .B1(new_n232), .B2(G131), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n227), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n215), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT71), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  XOR2_X1   g051(.A(KEYINPUT2), .B(G113), .Z(new_n238));
  XNOR2_X1  g052(.A(G116), .B(G119), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT67), .ZN(new_n241));
  INV_X1    g055(.A(G119), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G116), .ZN(new_n243));
  INV_X1    g057(.A(G116), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G119), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT2), .B(G113), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n240), .A2(new_n241), .A3(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n246), .A2(new_n247), .A3(KEYINPUT67), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n215), .A2(KEYINPUT71), .A3(new_n234), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n237), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT28), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n215), .A2(new_n234), .A3(new_n251), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n251), .B1(new_n215), .B2(new_n234), .ZN(new_n258));
  OAI21_X1  g072(.A(KEYINPUT28), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  XOR2_X1   g073(.A(KEYINPUT69), .B(KEYINPUT27), .Z(new_n260));
  INV_X1    g074(.A(G237), .ZN(new_n261));
  INV_X1    g075(.A(G953), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n261), .A2(new_n262), .A3(G210), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n260), .B(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT26), .B(G101), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n264), .B(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT29), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n255), .A2(new_n259), .A3(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT72), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n255), .A2(KEYINPUT72), .A3(new_n259), .A4(new_n268), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  XOR2_X1   g087(.A(KEYINPUT73), .B(G902), .Z(new_n274));
  INV_X1    g088(.A(new_n251), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n275), .B1(new_n235), .B2(new_n236), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT28), .B1(new_n276), .B2(new_n252), .ZN(new_n277));
  AOI21_X1  g091(.A(G146), .B1(new_n217), .B2(new_n219), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n209), .B1(new_n278), .B2(new_n203), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n220), .A2(new_n210), .A3(new_n207), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n199), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n234), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n275), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n254), .B1(new_n256), .B2(new_n283), .ZN(new_n284));
  NOR3_X1   g098(.A1(new_n277), .A2(new_n284), .A3(new_n266), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n215), .A2(KEYINPUT30), .A3(new_n234), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT30), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n282), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n286), .A2(new_n288), .A3(new_n275), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n256), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n266), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n267), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n274), .B1(new_n285), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(G472), .B1(new_n273), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n266), .ZN(new_n295));
  INV_X1    g109(.A(new_n284), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n295), .B1(new_n255), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n232), .A2(G131), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(new_n198), .ZN(new_n299));
  INV_X1    g113(.A(new_n226), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n206), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n299), .B1(new_n301), .B2(new_n223), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n194), .A2(new_n198), .A3(KEYINPUT68), .ZN(new_n303));
  AOI21_X1  g117(.A(KEYINPUT68), .B1(new_n194), .B2(new_n198), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n302), .B1(new_n305), .B2(new_n213), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n266), .B1(new_n306), .B2(new_n251), .ZN(new_n307));
  AND3_X1   g121(.A1(new_n307), .A2(KEYINPUT70), .A3(new_n289), .ZN(new_n308));
  AOI21_X1  g122(.A(KEYINPUT70), .B1(new_n307), .B2(new_n289), .ZN(new_n309));
  OAI21_X1  g123(.A(KEYINPUT31), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(KEYINPUT31), .B1(new_n307), .B2(new_n289), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n297), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(G472), .A2(G902), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  NOR3_X1   g129(.A1(new_n313), .A2(KEYINPUT32), .A3(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT32), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n266), .B1(new_n277), .B2(new_n284), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT31), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT70), .ZN(new_n320));
  AND3_X1   g134(.A1(new_n286), .A2(new_n288), .A3(new_n275), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n295), .A2(new_n256), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n307), .A2(KEYINPUT70), .A3(new_n289), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n319), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n318), .B1(new_n325), .B2(new_n311), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n317), .B1(new_n326), .B2(new_n314), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n294), .B1(new_n316), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G217), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n329), .B1(new_n274), .B2(G234), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n221), .A2(G119), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n242), .A2(G128), .ZN(new_n333));
  AND2_X1   g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  XOR2_X1   g148(.A(KEYINPUT24), .B(G110), .Z(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OR2_X1    g150(.A1(new_n336), .A2(KEYINPUT74), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(KEYINPUT74), .ZN(new_n338));
  AND2_X1   g152(.A1(new_n333), .A2(KEYINPUT23), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n332), .A2(KEYINPUT75), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT75), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n341), .A2(KEYINPUT23), .ZN(new_n342));
  OAI22_X1  g156(.A1(new_n339), .A2(new_n340), .B1(new_n342), .B2(new_n332), .ZN(new_n343));
  AOI22_X1  g157(.A1(new_n337), .A2(new_n338), .B1(G110), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(G140), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(G125), .ZN(new_n346));
  INV_X1    g160(.A(G125), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G140), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n346), .A2(new_n348), .A3(KEYINPUT76), .ZN(new_n349));
  OR3_X1    g163(.A1(new_n347), .A2(KEYINPUT76), .A3(G140), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n349), .A2(new_n350), .A3(KEYINPUT16), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT16), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n346), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(G146), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n351), .A2(new_n202), .A3(new_n353), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n344), .A2(new_n357), .ZN(new_n358));
  OAI22_X1  g172(.A1(new_n343), .A2(G110), .B1(new_n334), .B2(new_n335), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n346), .A2(new_n348), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT77), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n346), .A2(new_n348), .A3(KEYINPUT77), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n359), .B(new_n355), .C1(G146), .C2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n358), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n262), .A2(G221), .A3(G234), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n367), .B(KEYINPUT78), .ZN(new_n368));
  XNOR2_X1  g182(.A(KEYINPUT22), .B(G137), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n368), .B(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n366), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n358), .A2(new_n365), .A3(new_n370), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n372), .A2(new_n274), .A3(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT25), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT79), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  OR2_X1    g191(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n374), .A2(new_n377), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n331), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n372), .A2(new_n373), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n330), .A2(G902), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n380), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(G107), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G104), .ZN(new_n387));
  INV_X1    g201(.A(G104), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(G107), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G101), .ZN(new_n391));
  OAI21_X1  g205(.A(KEYINPUT3), .B1(new_n388), .B2(G107), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT3), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(new_n386), .A3(G104), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n392), .A2(new_n394), .A3(new_n389), .ZN(new_n395));
  XNOR2_X1  g209(.A(KEYINPUT83), .B(G101), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n391), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n239), .A2(KEYINPUT5), .ZN(new_n399));
  INV_X1    g213(.A(G113), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n244), .A2(G119), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT5), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  AOI22_X1  g217(.A1(new_n399), .A2(new_n403), .B1(new_n238), .B2(new_n239), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n398), .A2(new_n404), .ZN(new_n405));
  AND3_X1   g219(.A1(new_n395), .A2(KEYINPUT82), .A3(G101), .ZN(new_n406));
  OAI21_X1  g220(.A(KEYINPUT4), .B1(new_n395), .B2(new_n396), .ZN(new_n407));
  AOI21_X1  g221(.A(KEYINPUT82), .B1(new_n395), .B2(G101), .ZN(new_n408));
  NOR3_X1   g222(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT4), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n395), .A2(new_n410), .A3(G101), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n249), .A2(new_n250), .A3(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n405), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(G110), .B(G122), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n405), .B(new_n414), .C1(new_n409), .C2(new_n412), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n416), .A2(KEYINPUT6), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n279), .A2(new_n280), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G125), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n420), .B1(G125), .B2(new_n227), .ZN(new_n421));
  INV_X1    g235(.A(G224), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n422), .A2(G953), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n421), .B(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT6), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n413), .A2(new_n425), .A3(new_n415), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n418), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n227), .A2(G125), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n347), .B1(new_n279), .B2(new_n280), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT7), .ZN(new_n430));
  OAI22_X1  g244(.A1(new_n428), .A2(new_n429), .B1(new_n430), .B2(new_n423), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n423), .A2(new_n430), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n420), .B(new_n432), .C1(G125), .C2(new_n227), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT8), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n414), .B(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n435), .B1(new_n397), .B2(new_n404), .ZN(new_n436));
  OAI21_X1  g250(.A(G113), .B1(new_n243), .B2(KEYINPUT5), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n437), .B1(new_n399), .B2(KEYINPUT87), .ZN(new_n438));
  OR3_X1    g252(.A1(new_n246), .A2(KEYINPUT87), .A3(new_n402), .ZN(new_n439));
  AOI22_X1  g253(.A1(new_n438), .A2(new_n439), .B1(new_n239), .B2(new_n238), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n436), .B1(new_n440), .B2(new_n397), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n431), .A2(new_n433), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(G902), .B1(new_n442), .B2(new_n417), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n427), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(G210), .B1(G237), .B2(G902), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n427), .A2(new_n443), .A3(new_n445), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n447), .A2(KEYINPUT88), .A3(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT88), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n444), .A2(new_n450), .A3(new_n446), .ZN(new_n451));
  OAI21_X1  g265(.A(G214), .B1(G237), .B2(G902), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n452), .B(KEYINPUT86), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n262), .A2(G952), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n455), .B1(G234), .B2(G237), .ZN(new_n456));
  AOI211_X1 g270(.A(new_n262), .B(new_n274), .C1(G234), .C2(G237), .ZN(new_n457));
  XNOR2_X1  g271(.A(KEYINPUT21), .B(G898), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n456), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n449), .A2(new_n451), .A3(new_n454), .A4(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT93), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT20), .ZN(new_n463));
  XOR2_X1   g277(.A(G113), .B(G122), .Z(new_n464));
  XOR2_X1   g278(.A(KEYINPUT90), .B(G104), .Z(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g280(.A(G113), .B(G122), .ZN(new_n467));
  XNOR2_X1  g281(.A(KEYINPUT90), .B(G104), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n261), .A2(new_n262), .A3(G143), .A4(G214), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n261), .A2(new_n262), .A3(G214), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n197), .B(new_n471), .C1(new_n224), .C2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(KEYINPUT89), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n471), .B1(new_n224), .B2(new_n472), .ZN(new_n475));
  INV_X1    g289(.A(new_n197), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n261), .A2(new_n262), .A3(G214), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n205), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT89), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n479), .A2(new_n480), .A3(new_n197), .A4(new_n471), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n474), .A2(new_n477), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n349), .A2(new_n350), .A3(KEYINPUT19), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n483), .B1(new_n364), .B2(KEYINPUT19), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n482), .B(new_n355), .C1(G146), .C2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT18), .ZN(new_n486));
  INV_X1    g300(.A(G131), .ZN(new_n487));
  NOR3_X1   g301(.A1(new_n475), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  AOI22_X1  g302(.A1(new_n479), .A2(new_n471), .B1(KEYINPUT18), .B2(G131), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n364), .A2(G146), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n349), .A2(G146), .A3(new_n350), .ZN(new_n491));
  OAI22_X1  g305(.A1(new_n488), .A2(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n470), .B1(new_n485), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT91), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n470), .B(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT17), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n474), .A2(new_n477), .A3(new_n481), .A4(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n475), .A2(KEYINPUT17), .A3(new_n476), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n355), .A2(new_n356), .A3(new_n499), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n492), .B(new_n495), .C1(new_n498), .C2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT92), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n497), .A2(new_n356), .A3(new_n355), .A4(new_n499), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n504), .A2(KEYINPUT92), .A3(new_n492), .A4(new_n495), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n493), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(G475), .A2(G902), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n462), .B(new_n463), .C1(new_n506), .C2(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n470), .B1(new_n504), .B2(new_n492), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n510), .B1(new_n503), .B2(new_n505), .ZN(new_n511));
  OAI21_X1  g325(.A(G475), .B1(new_n511), .B2(G902), .ZN(new_n512));
  AND2_X1   g326(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  XOR2_X1   g327(.A(KEYINPUT94), .B(KEYINPUT13), .Z(new_n514));
  NAND3_X1  g328(.A1(new_n217), .A2(new_n219), .A3(G128), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n221), .A2(G143), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(G134), .B1(new_n514), .B2(new_n515), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n515), .A2(new_n188), .A3(new_n516), .ZN(new_n520));
  XOR2_X1   g334(.A(G116), .B(G122), .Z(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n386), .ZN(new_n522));
  XNOR2_X1  g336(.A(G116), .B(G122), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(G107), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n520), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(KEYINPUT95), .B1(new_n519), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n527), .B(G134), .C1(new_n514), .C2(new_n515), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n520), .A2(new_n522), .A3(new_n524), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT95), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  OR2_X1    g346(.A1(new_n244), .A2(G122), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n386), .B1(new_n533), .B2(KEYINPUT14), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n534), .B(new_n523), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n515), .A2(new_n516), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(G134), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n520), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n532), .A2(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(KEYINPUT9), .B(G234), .ZN(new_n541));
  NOR3_X1   g355(.A1(new_n541), .A2(new_n329), .A3(G953), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  NOR3_X1   g358(.A1(new_n519), .A2(new_n525), .A3(KEYINPUT95), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n530), .B1(new_n528), .B2(new_n529), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n539), .B(new_n542), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n274), .ZN(new_n549));
  INV_X1    g363(.A(G478), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n550), .A2(KEYINPUT15), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n551), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n553), .B1(new_n548), .B2(new_n274), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n503), .A2(new_n505), .ZN(new_n556));
  INV_X1    g370(.A(new_n493), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n558), .A2(KEYINPUT93), .A3(new_n507), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n462), .B1(new_n506), .B2(new_n508), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(KEYINPUT20), .A3(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n513), .A2(new_n555), .A3(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n461), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(G221), .B1(new_n541), .B2(G902), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(G469), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n220), .A2(new_n210), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT1), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n278), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n567), .B1(new_n569), .B2(new_n221), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n397), .B1(new_n570), .B2(new_n223), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n398), .A2(new_n227), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n199), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(KEYINPUT1), .B1(new_n205), .B2(G146), .ZN(new_n574));
  AOI22_X1  g388(.A1(new_n574), .A2(G128), .B1(new_n210), .B2(new_n220), .ZN(new_n575));
  INV_X1    g389(.A(new_n223), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n398), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n577), .B1(new_n227), .B2(new_n398), .ZN(new_n578));
  NOR3_X1   g392(.A1(new_n303), .A2(new_n304), .A3(KEYINPUT12), .ZN(new_n579));
  AOI22_X1  g393(.A1(new_n573), .A2(KEYINPUT12), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT10), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n581), .B1(new_n301), .B2(new_n223), .ZN(new_n582));
  AOI22_X1  g396(.A1(new_n577), .A2(new_n581), .B1(new_n398), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n305), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT84), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n279), .A2(new_n411), .A3(new_n280), .ZN(new_n586));
  NOR3_X1   g400(.A1(new_n409), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n395), .ZN(new_n588));
  INV_X1    g402(.A(new_n396), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n410), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n395), .A2(G101), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT82), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n395), .A2(KEYINPUT82), .A3(G101), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n590), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n586), .ZN(new_n596));
  AOI21_X1  g410(.A(KEYINPUT84), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n583), .B(new_n584), .C1(new_n587), .C2(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(G110), .B(G140), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(KEYINPUT80), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n262), .A2(G227), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n600), .B(new_n601), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n580), .A2(new_n598), .A3(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n602), .ZN(new_n604));
  INV_X1    g418(.A(new_n598), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n585), .B1(new_n409), .B2(new_n586), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n595), .A2(new_n596), .A3(KEYINPUT84), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n584), .B1(new_n608), .B2(new_n583), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n604), .B1(new_n605), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT85), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n603), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n580), .A2(new_n598), .A3(new_n602), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n613), .A2(KEYINPUT85), .ZN(new_n614));
  OAI211_X1 g428(.A(new_n566), .B(new_n274), .C1(new_n612), .C2(new_n614), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n605), .A2(new_n609), .A3(new_n604), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n602), .B(KEYINPUT81), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n618), .B1(new_n580), .B2(new_n598), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g434(.A(G469), .B1(new_n620), .B2(G902), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n565), .B1(new_n615), .B2(new_n621), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n328), .A2(new_n385), .A3(new_n563), .A4(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(KEYINPUT96), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(new_n396), .ZN(G3));
  NAND2_X1  g439(.A1(new_n326), .A2(new_n274), .ZN(new_n626));
  AOI22_X1  g440(.A1(new_n626), .A2(G472), .B1(new_n314), .B2(new_n326), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n627), .A2(new_n385), .A3(new_n622), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT33), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n629), .B1(new_n547), .B2(KEYINPUT99), .ZN(new_n630));
  INV_X1    g444(.A(new_n547), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n542), .B1(new_n532), .B2(new_n539), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI211_X1 g447(.A(new_n544), .B(new_n547), .C1(KEYINPUT99), .C2(new_n629), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n274), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n636), .A2(new_n550), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n549), .A2(new_n550), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AND3_X1   g454(.A1(new_n559), .A2(KEYINPUT20), .A3(new_n560), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n509), .A2(new_n512), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT98), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n447), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n445), .B1(new_n427), .B2(new_n443), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(KEYINPUT98), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n448), .A2(KEYINPUT97), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT97), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n427), .A2(new_n443), .A3(new_n649), .A4(new_n445), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n645), .A2(new_n647), .A3(new_n648), .A4(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n651), .A2(new_n454), .A3(new_n460), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n628), .A2(new_n643), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G104), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT100), .B(KEYINPUT34), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G6));
  OAI211_X1 g470(.A(new_n513), .B(new_n561), .C1(new_n554), .C2(new_n552), .ZN(new_n657));
  NOR3_X1   g471(.A1(new_n628), .A2(new_n652), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G107), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT101), .B(KEYINPUT35), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G9));
  NOR2_X1   g475(.A1(new_n371), .A2(KEYINPUT36), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n366), .B(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n664), .A2(new_n383), .ZN(new_n665));
  OR2_X1    g479(.A1(new_n380), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n563), .A2(new_n627), .A3(new_n622), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT102), .ZN(new_n668));
  XOR2_X1   g482(.A(KEYINPUT37), .B(G110), .Z(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G12));
  NAND2_X1  g484(.A1(new_n615), .A2(new_n621), .ZN(new_n671));
  AND4_X1   g485(.A1(new_n564), .A2(new_n671), .A3(new_n454), .A4(new_n651), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n380), .A2(new_n665), .ZN(new_n673));
  OAI21_X1  g487(.A(KEYINPUT32), .B1(new_n313), .B2(new_n315), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n326), .A2(new_n317), .A3(new_n314), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n673), .B1(new_n676), .B2(new_n294), .ZN(new_n677));
  INV_X1    g491(.A(G900), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n456), .B1(new_n457), .B2(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n657), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n672), .A2(new_n677), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G128), .ZN(G30));
  OAI21_X1  g496(.A(new_n266), .B1(new_n257), .B2(new_n258), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n323), .A2(new_n324), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g498(.A(G472), .B1(new_n684), .B2(G902), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n685), .B1(new_n316), .B2(new_n327), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(KEYINPUT104), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT104), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n676), .A2(new_n688), .A3(new_n685), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g504(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n448), .A2(KEYINPUT88), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n693), .A2(new_n646), .ZN(new_n694));
  INV_X1    g508(.A(new_n451), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n692), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n555), .B1(new_n513), .B2(new_n561), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n380), .A2(new_n453), .A3(new_n665), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n449), .A2(new_n451), .A3(new_n691), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n696), .A2(new_n697), .A3(new_n698), .A4(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT40), .ZN(new_n701));
  XOR2_X1   g515(.A(new_n679), .B(KEYINPUT39), .Z(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  AOI211_X1 g517(.A(new_n565), .B(new_n703), .C1(new_n615), .C2(new_n621), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n700), .B1(new_n701), .B2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(new_n622), .ZN(new_n706));
  OAI21_X1  g520(.A(KEYINPUT40), .B1(new_n706), .B2(new_n703), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n690), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(new_n224), .ZN(G45));
  NOR2_X1   g523(.A1(new_n643), .A2(new_n679), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n672), .A2(new_n677), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G146), .ZN(G48));
  INV_X1    g526(.A(new_n385), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n713), .B1(new_n676), .B2(new_n294), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n652), .A2(new_n643), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n274), .B1(new_n612), .B2(new_n614), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(G469), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(new_n564), .A3(new_n615), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n714), .A2(new_n715), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(KEYINPUT41), .B(G113), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n720), .B(new_n721), .ZN(G15));
  NOR2_X1   g536(.A1(new_n652), .A2(new_n657), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n714), .A2(new_n723), .A3(new_n719), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G116), .ZN(G18));
  NAND2_X1  g539(.A1(new_n651), .A2(new_n454), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n718), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n562), .A2(new_n459), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n727), .A2(new_n677), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G119), .ZN(G21));
  AND4_X1   g544(.A1(new_n564), .A2(new_n717), .A3(new_n615), .A4(new_n460), .ZN(new_n731));
  OAI21_X1  g545(.A(G472), .B1(new_n313), .B2(new_n636), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT105), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n295), .B1(new_n255), .B2(new_n259), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n734), .B1(new_n310), .B2(new_n312), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n733), .B1(new_n735), .B2(new_n315), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n323), .A2(new_n324), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n311), .B1(new_n737), .B2(KEYINPUT31), .ZN(new_n738));
  OAI211_X1 g552(.A(KEYINPUT105), .B(new_n314), .C1(new_n738), .C2(new_n734), .ZN(new_n739));
  AND4_X1   g553(.A1(new_n385), .A2(new_n732), .A3(new_n736), .A4(new_n739), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n697), .A2(new_n454), .A3(new_n651), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n731), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  XOR2_X1   g556(.A(KEYINPUT106), .B(G122), .Z(new_n743));
  XNOR2_X1  g557(.A(new_n742), .B(new_n743), .ZN(G24));
  AND4_X1   g558(.A1(new_n732), .A2(new_n666), .A3(new_n736), .A4(new_n739), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n727), .A2(new_n745), .A3(new_n710), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G125), .ZN(G27));
  INV_X1    g561(.A(KEYINPUT108), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n748), .B1(new_n316), .B2(new_n327), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n674), .A2(KEYINPUT108), .A3(new_n675), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(new_n294), .A3(new_n750), .ZN(new_n751));
  AOI22_X1  g565(.A1(new_n513), .A2(new_n561), .B1(new_n639), .B2(new_n638), .ZN(new_n752));
  INV_X1    g566(.A(new_n679), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  OAI211_X1 g568(.A(new_n564), .B(new_n454), .C1(new_n694), .C2(new_n695), .ZN(new_n755));
  NAND2_X1  g569(.A1(G469), .A2(G902), .ZN(new_n756));
  XOR2_X1   g570(.A(new_n756), .B(KEYINPUT107), .Z(new_n757));
  NAND2_X1  g571(.A1(new_n580), .A2(new_n598), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n617), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n583), .B1(new_n587), .B2(new_n597), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n305), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(new_n598), .A3(new_n602), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n757), .B1(new_n763), .B2(new_n566), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n602), .B1(new_n761), .B2(new_n598), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n613), .B1(new_n765), .B2(KEYINPUT85), .ZN(new_n766));
  INV_X1    g580(.A(new_n614), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n636), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n764), .B1(new_n768), .B2(new_n566), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n754), .A2(new_n755), .A3(new_n769), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n751), .A2(new_n770), .A3(KEYINPUT42), .A4(new_n385), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n755), .A2(new_n769), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n772), .A2(new_n328), .A3(new_n710), .A4(new_n385), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT42), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT109), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n771), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n776), .B1(new_n771), .B2(new_n775), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G131), .ZN(G33));
  NAND3_X1  g595(.A1(new_n714), .A2(new_n680), .A3(new_n772), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G134), .ZN(G36));
  NAND2_X1  g597(.A1(new_n326), .A2(new_n314), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n673), .B1(new_n732), .B2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n640), .A2(new_n513), .A3(new_n561), .ZN(new_n786));
  AND2_X1   g600(.A1(KEYINPUT111), .A2(KEYINPUT43), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(KEYINPUT111), .A2(KEYINPUT43), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n640), .A2(new_n513), .A3(new_n561), .A4(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n785), .A2(KEYINPUT44), .A3(new_n788), .A4(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n453), .B1(new_n449), .B2(new_n451), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(KEYINPUT112), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT45), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n796), .B1(new_n616), .B2(new_n619), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n759), .A2(new_n762), .A3(KEYINPUT45), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n797), .A2(G469), .A3(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n799), .A2(KEYINPUT46), .A3(new_n757), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(KEYINPUT110), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT110), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n799), .A2(new_n802), .A3(KEYINPUT46), .A4(new_n757), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT46), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n759), .A2(new_n762), .A3(KEYINPUT45), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT45), .B1(new_n759), .B2(new_n762), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n805), .A2(new_n806), .A3(new_n566), .ZN(new_n807));
  INV_X1    g621(.A(new_n757), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n804), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n801), .A2(new_n615), .A3(new_n803), .A4(new_n809), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n810), .A2(new_n564), .A3(new_n702), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT112), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n792), .A2(new_n812), .A3(new_n793), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT44), .ZN(new_n814));
  INV_X1    g628(.A(new_n785), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n788), .A2(new_n791), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n795), .A2(new_n811), .A3(new_n813), .A4(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(G137), .ZN(G39));
  NAND2_X1  g633(.A1(new_n713), .A2(new_n793), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n328), .A2(new_n754), .A3(new_n820), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n810), .A2(KEYINPUT47), .A3(new_n564), .ZN(new_n822));
  AOI21_X1  g636(.A(KEYINPUT47), .B1(new_n810), .B2(new_n564), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(G140), .ZN(G42));
  NOR2_X1   g639(.A1(new_n768), .A2(new_n566), .ZN(new_n826));
  INV_X1    g640(.A(new_n615), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(KEYINPUT49), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n694), .A2(new_n695), .A3(new_n692), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n691), .B1(new_n449), .B2(new_n451), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n385), .A2(new_n564), .A3(new_n454), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n832), .A2(new_n786), .A3(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n829), .A2(new_n687), .A3(new_n689), .A4(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n461), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n627), .A2(new_n836), .A3(new_n622), .A4(new_n385), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n667), .B1(new_n837), .B2(new_n657), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n643), .A2(KEYINPUT113), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT113), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n752), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n837), .A2(new_n842), .ZN(new_n843));
  AND4_X1   g657(.A1(new_n328), .A2(new_n385), .A3(new_n622), .A4(new_n563), .ZN(new_n844));
  OAI21_X1  g658(.A(KEYINPUT114), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT114), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n623), .B(new_n846), .C1(new_n837), .C2(new_n842), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n838), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n729), .A2(new_n720), .A3(new_n724), .A4(new_n742), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n622), .A2(new_n793), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT115), .ZN(new_n851));
  OR3_X1    g665(.A1(new_n562), .A2(new_n851), .A3(new_n679), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n851), .B1(new_n562), .B2(new_n679), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n677), .A2(new_n850), .A3(new_n852), .A4(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n745), .A2(new_n710), .A3(new_n772), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n854), .A2(new_n782), .A3(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n849), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n771), .A2(new_n775), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(KEYINPUT109), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n848), .A2(new_n857), .A3(new_n859), .A4(new_n777), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n672), .B(new_n677), .C1(new_n680), .C2(new_n710), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n679), .A2(KEYINPUT116), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n564), .B1(new_n679), .B2(KEYINPUT116), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n666), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n769), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n741), .A2(new_n864), .A3(new_n686), .A4(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n861), .A2(new_n746), .A3(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT52), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n861), .A2(KEYINPUT52), .A3(new_n746), .A4(new_n866), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT53), .B1(new_n860), .B2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT117), .ZN(new_n873));
  AOI22_X1  g687(.A1(new_n869), .A2(new_n870), .B1(new_n873), .B2(new_n867), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n867), .A2(new_n873), .A3(KEYINPUT52), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT53), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n780), .A2(new_n877), .A3(new_n848), .A4(new_n857), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n872), .B(KEYINPUT54), .C1(new_n876), .C2(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n877), .B1(new_n860), .B2(new_n871), .ZN(new_n880));
  INV_X1    g694(.A(new_n849), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n877), .B1(new_n771), .B2(new_n775), .ZN(new_n882));
  INV_X1    g696(.A(new_n856), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n848), .B(new_n884), .C1(new_n874), .C2(new_n875), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT54), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n880), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n788), .A2(new_n791), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n717), .A2(new_n615), .A3(new_n456), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n889), .A2(new_n755), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n751), .A2(new_n888), .A3(new_n385), .A4(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(KEYINPUT48), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n816), .A2(new_n755), .A3(new_n889), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT48), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n893), .A2(new_n894), .A3(new_n385), .A4(new_n751), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n889), .A2(new_n713), .A3(new_n755), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n897), .A2(new_n687), .A3(new_n689), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n455), .B1(new_n898), .B2(new_n752), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n888), .A2(new_n727), .A3(new_n456), .A4(new_n740), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(KEYINPUT120), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n732), .A2(new_n736), .A3(new_n385), .A4(new_n739), .ZN(new_n902));
  INV_X1    g716(.A(new_n456), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n816), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT120), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n904), .A2(new_n905), .A3(new_n727), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n901), .A2(new_n906), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n896), .A2(new_n899), .A3(new_n907), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n826), .A2(new_n827), .A3(new_n564), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n822), .A2(new_n823), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n904), .A2(new_n793), .ZN(new_n911));
  OAI21_X1  g725(.A(KEYINPUT51), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n641), .A2(new_n640), .A3(new_n642), .ZN(new_n913));
  AOI22_X1  g727(.A1(new_n898), .A2(new_n913), .B1(new_n745), .B2(new_n893), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n453), .B1(new_n830), .B2(new_n831), .ZN(new_n915));
  OAI21_X1  g729(.A(KEYINPUT119), .B1(new_n915), .B2(new_n718), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n454), .B1(new_n696), .B2(new_n699), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT119), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n719), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n920), .A2(KEYINPUT50), .A3(new_n904), .ZN(new_n921));
  AOI21_X1  g735(.A(KEYINPUT50), .B1(new_n920), .B2(new_n904), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n914), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n908), .B1(new_n912), .B2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT51), .ZN(new_n925));
  INV_X1    g739(.A(new_n911), .ZN(new_n926));
  OR2_X1    g740(.A1(new_n822), .A2(new_n823), .ZN(new_n927));
  OAI211_X1 g741(.A(KEYINPUT118), .B(new_n926), .C1(new_n927), .C2(new_n909), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT118), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n929), .B1(new_n910), .B2(new_n911), .ZN(new_n930));
  INV_X1    g744(.A(new_n922), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n920), .A2(KEYINPUT50), .A3(new_n904), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n928), .A2(new_n930), .A3(new_n933), .A4(new_n914), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n924), .B1(new_n925), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n879), .A2(new_n887), .A3(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT121), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n879), .A2(new_n935), .A3(new_n887), .A4(KEYINPUT121), .ZN(new_n939));
  OR2_X1    g753(.A1(G952), .A2(G953), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n835), .B1(new_n938), .B2(new_n941), .ZN(G75));
  AOI21_X1  g756(.A(new_n274), .B1(new_n880), .B2(new_n885), .ZN(new_n943));
  AOI21_X1  g757(.A(KEYINPUT56), .B1(new_n943), .B2(new_n446), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n418), .A2(new_n426), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(new_n424), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT55), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n262), .A2(G952), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n950), .B1(new_n944), .B2(new_n947), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n948), .A2(new_n951), .ZN(G51));
  INV_X1    g766(.A(KEYINPUT122), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n880), .A2(new_n885), .ZN(new_n954));
  AND4_X1   g768(.A1(new_n953), .A2(new_n954), .A3(new_n636), .A4(new_n807), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n953), .B1(new_n943), .B2(new_n807), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n757), .B(KEYINPUT57), .Z(new_n958));
  AND3_X1   g772(.A1(new_n880), .A2(new_n885), .A3(new_n886), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n886), .B1(new_n880), .B2(new_n885), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n958), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n766), .A2(new_n767), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n949), .B1(new_n957), .B2(new_n963), .ZN(G54));
  AND2_X1   g778(.A1(KEYINPUT58), .A2(G475), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n943), .A2(new_n558), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n558), .B1(new_n943), .B2(new_n965), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n966), .A2(new_n967), .A3(new_n949), .ZN(G60));
  NAND2_X1  g782(.A1(G478), .A2(G902), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT59), .Z(new_n970));
  AOI21_X1  g784(.A(new_n970), .B1(new_n879), .B2(new_n887), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n971), .A2(new_n635), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n970), .B1(new_n633), .B2(new_n634), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n973), .B1(new_n959), .B2(new_n960), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(new_n950), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n972), .A2(new_n975), .ZN(G63));
  INV_X1    g790(.A(KEYINPUT61), .ZN(new_n977));
  NAND2_X1  g791(.A1(G217), .A2(G902), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT60), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n979), .B1(new_n880), .B2(new_n885), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n663), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(new_n381), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n950), .B1(new_n980), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n977), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n979), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n954), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n949), .B1(new_n987), .B2(new_n381), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n988), .A2(KEYINPUT61), .A3(new_n981), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n985), .A2(new_n989), .ZN(G66));
  OAI21_X1  g804(.A(G953), .B1(new_n458), .B2(new_n422), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n848), .A2(new_n881), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n991), .B1(new_n992), .B2(G953), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n945), .B1(G898), .B2(new_n262), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n993), .B(new_n994), .ZN(G69));
  NAND2_X1  g809(.A1(new_n286), .A2(new_n288), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n996), .B(new_n484), .ZN(new_n997));
  INV_X1    g811(.A(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT62), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n708), .A2(new_n999), .A3(new_n746), .A4(new_n861), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n842), .A2(new_n657), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n1001), .A2(new_n714), .A3(new_n704), .A4(new_n793), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n1000), .A2(new_n818), .A3(new_n824), .A4(new_n1002), .ZN(new_n1003));
  AND3_X1   g817(.A1(new_n676), .A2(new_n688), .A3(new_n685), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n688), .B1(new_n676), .B2(new_n685), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n707), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n704), .A2(new_n701), .ZN(new_n1007));
  NAND4_X1  g821(.A1(new_n1007), .A2(new_n832), .A3(new_n697), .A4(new_n698), .ZN(new_n1008));
  OAI211_X1 g822(.A(new_n746), .B(new_n861), .C1(new_n1006), .C2(new_n1008), .ZN(new_n1009));
  INV_X1    g823(.A(KEYINPUT123), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n1009), .A2(new_n1010), .A3(KEYINPUT62), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1009), .A2(KEYINPUT62), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1012), .A2(KEYINPUT123), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1003), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n998), .B1(new_n1014), .B2(G953), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n262), .B1(G227), .B2(G900), .ZN(new_n1016));
  AND3_X1   g830(.A1(new_n861), .A2(new_n746), .A3(new_n782), .ZN(new_n1017));
  AND2_X1   g831(.A1(new_n751), .A2(new_n385), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n811), .A2(new_n1018), .A3(new_n741), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n824), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g834(.A(new_n1020), .ZN(new_n1021));
  NAND4_X1  g835(.A1(new_n1021), .A2(new_n780), .A3(new_n262), .A4(new_n818), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n998), .B1(G900), .B2(G953), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1016), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1015), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g839(.A(KEYINPUT124), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n1022), .A2(new_n1026), .A3(new_n1023), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n859), .A2(new_n818), .A3(new_n777), .ZN(new_n1028));
  NOR3_X1   g842(.A1(new_n1028), .A2(new_n1020), .A3(G953), .ZN(new_n1029));
  INV_X1    g843(.A(new_n1023), .ZN(new_n1030));
  OAI21_X1  g844(.A(KEYINPUT124), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n1015), .A2(new_n1027), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g846(.A(KEYINPUT125), .ZN(new_n1033));
  AND3_X1   g847(.A1(new_n1032), .A2(new_n1033), .A3(new_n1016), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n1033), .B1(new_n1032), .B2(new_n1016), .ZN(new_n1035));
  OAI21_X1  g849(.A(new_n1025), .B1(new_n1034), .B2(new_n1035), .ZN(G72));
  NAND2_X1  g850(.A1(G472), .A2(G902), .ZN(new_n1037));
  XOR2_X1   g851(.A(new_n1037), .B(KEYINPUT63), .Z(new_n1038));
  INV_X1    g852(.A(new_n1038), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n1039), .B1(new_n1014), .B2(new_n992), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n290), .A2(new_n295), .ZN(new_n1041));
  OAI21_X1  g855(.A(new_n872), .B1(new_n876), .B2(new_n878), .ZN(new_n1042));
  INV_X1    g856(.A(new_n291), .ZN(new_n1043));
  AOI21_X1  g857(.A(new_n737), .B1(KEYINPUT127), .B2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g858(.A(new_n1044), .B1(KEYINPUT127), .B2(new_n1043), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n1045), .A2(new_n1038), .ZN(new_n1046));
  OAI22_X1  g860(.A1(new_n1040), .A2(new_n1041), .B1(new_n1042), .B2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g861(.A1(new_n1028), .A2(new_n1020), .ZN(new_n1048));
  AOI21_X1  g862(.A(new_n1039), .B1(new_n1048), .B2(new_n992), .ZN(new_n1049));
  NAND3_X1  g863(.A1(new_n289), .A2(new_n256), .A3(new_n266), .ZN(new_n1050));
  OAI21_X1  g864(.A(new_n950), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g865(.A(KEYINPUT126), .ZN(new_n1052));
  OR2_X1    g866(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g867(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1054));
  AOI21_X1  g868(.A(new_n1047), .B1(new_n1053), .B2(new_n1054), .ZN(G57));
endmodule


