//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 1 1 1 1 1 0 1 1 0 1 0 0 1 1 0 0 0 1 0 0 1 1 1 1 0 1 0 0 1 0 1 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:41 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n580, new_n581, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n594, new_n595,
    new_n597, new_n598, new_n599, new_n600, new_n602, new_n603, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n633, new_n634, new_n635, new_n636, new_n639,
    new_n641, new_n642, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1226,
    new_n1227, new_n1228, new_n1229;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT64), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  NAND3_X1  g034(.A1(new_n459), .A2(G101), .A3(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT66), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n462));
  NAND4_X1  g037(.A1(new_n462), .A2(new_n459), .A3(G101), .A4(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  OAI211_X1 g041(.A(G137), .B(new_n459), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g043(.A(G125), .B1(new_n465), .B2(new_n466), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n459), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n468), .A2(new_n471), .ZN(G160));
  OAI21_X1  g047(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n473));
  INV_X1    g048(.A(G112), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n473), .B1(new_n474), .B2(G2105), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  XNOR2_X1  g051(.A(KEYINPUT3), .B(G2104), .ZN(new_n477));
  AND2_X1   g052(.A1(new_n477), .A2(KEYINPUT67), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n477), .A2(KEYINPUT67), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n459), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(G136), .ZN(new_n481));
  INV_X1    g056(.A(G124), .ZN(new_n482));
  OAI21_X1  g057(.A(G2105), .B1(new_n478), .B2(new_n479), .ZN(new_n483));
  OAI221_X1 g058(.A(new_n476), .B1(new_n480), .B2(new_n481), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  AND2_X1   g060(.A1(G126), .A2(G2105), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(G114), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  AOI22_X1  g065(.A1(new_n477), .A2(new_n486), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n465), .A2(new_n466), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT68), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n494), .A2(new_n459), .A3(G138), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n492), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  AND3_X1   g071(.A1(new_n494), .A2(new_n459), .A3(G138), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n477), .A2(new_n497), .A3(KEYINPUT4), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n491), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G543), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  AND3_X1   g078(.A1(new_n503), .A2(KEYINPUT69), .A3(KEYINPUT5), .ZN(new_n504));
  AOI21_X1  g079(.A(KEYINPUT69), .B1(new_n503), .B2(KEYINPUT5), .ZN(new_n505));
  OAI211_X1 g080(.A(G62), .B(new_n502), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(G75), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G651), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT71), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n508), .A2(KEYINPUT71), .A3(G651), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT69), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n513), .B1(new_n501), .B2(G543), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n503), .A2(KEYINPUT69), .A3(KEYINPUT5), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT6), .B(G651), .ZN(new_n517));
  NAND4_X1  g092(.A1(new_n516), .A2(G88), .A3(new_n502), .A4(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n517), .A2(G50), .A3(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(KEYINPUT70), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT70), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n518), .A2(new_n522), .A3(new_n519), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n511), .A2(new_n512), .B1(new_n521), .B2(new_n523), .ZN(G166));
  AOI22_X1  g099(.A1(new_n514), .A2(new_n515), .B1(new_n501), .B2(G543), .ZN(new_n525));
  AND2_X1   g100(.A1(G63), .A2(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT72), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n528), .B1(new_n517), .B2(G543), .ZN(new_n529));
  AND2_X1   g104(.A1(KEYINPUT6), .A2(G651), .ZN(new_n530));
  NOR2_X1   g105(.A1(KEYINPUT6), .A2(G651), .ZN(new_n531));
  OAI211_X1 g106(.A(new_n528), .B(G543), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g109(.A(KEYINPUT73), .B(G51), .ZN(new_n535));
  OAI211_X1 g110(.A(KEYINPUT74), .B(new_n527), .C1(new_n534), .C2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT74), .ZN(new_n537));
  OAI21_X1  g112(.A(G543), .B1(new_n530), .B2(new_n531), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(KEYINPUT72), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n535), .B1(new_n539), .B2(new_n532), .ZN(new_n540));
  AND2_X1   g115(.A1(new_n525), .A2(new_n526), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n537), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND4_X1  g117(.A1(new_n516), .A2(G89), .A3(new_n502), .A4(new_n517), .ZN(new_n543));
  NAND3_X1  g118(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(KEYINPUT75), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT75), .ZN(new_n546));
  NAND4_X1  g121(.A1(new_n546), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n545), .A2(KEYINPUT7), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n545), .A2(new_n547), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT7), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n543), .A2(new_n548), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(KEYINPUT76), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT76), .ZN(new_n554));
  NAND4_X1  g129(.A1(new_n543), .A2(new_n551), .A3(new_n554), .A4(new_n548), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n536), .A2(new_n542), .B1(new_n553), .B2(new_n555), .ZN(G168));
  AOI22_X1  g131(.A1(new_n525), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G651), .ZN(new_n558));
  OR2_X1    g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n525), .A2(new_n517), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  XNOR2_X1  g136(.A(KEYINPUT78), .B(G90), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n539), .A2(new_n532), .ZN(new_n564));
  XOR2_X1   g139(.A(KEYINPUT77), .B(G52), .Z(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n559), .A2(new_n563), .A3(new_n566), .ZN(G301));
  INV_X1    g142(.A(G301), .ZN(G171));
  NAND2_X1  g143(.A1(G68), .A2(G543), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n516), .A2(new_n502), .ZN(new_n570));
  INV_X1    g145(.A(G56), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G651), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n561), .A2(G81), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n564), .A2(G43), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(G860), .ZN(G153));
  NAND4_X1  g153(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g154(.A1(G1), .A2(G3), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT8), .ZN(new_n581));
  NAND4_X1  g156(.A1(G319), .A2(G483), .A3(G661), .A4(new_n581), .ZN(G188));
  INV_X1    g157(.A(KEYINPUT79), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n561), .A2(new_n583), .A3(G91), .ZN(new_n584));
  NAND2_X1  g159(.A1(G78), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G65), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n570), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(G651), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n517), .A2(G53), .A3(G543), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n589), .B(KEYINPUT9), .ZN(new_n590));
  INV_X1    g165(.A(G91), .ZN(new_n591));
  OAI21_X1  g166(.A(KEYINPUT79), .B1(new_n560), .B2(new_n591), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n584), .A2(new_n588), .A3(new_n590), .A4(new_n592), .ZN(G299));
  NAND2_X1  g168(.A1(new_n536), .A2(new_n542), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n553), .A2(new_n555), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(G286));
  AOI21_X1  g171(.A(KEYINPUT71), .B1(new_n508), .B2(G651), .ZN(new_n597));
  AOI211_X1 g172(.A(new_n510), .B(new_n558), .C1(new_n506), .C2(new_n507), .ZN(new_n598));
  AND3_X1   g173(.A1(new_n518), .A2(new_n522), .A3(new_n519), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n522), .B1(new_n518), .B2(new_n519), .ZN(new_n600));
  OAI22_X1  g175(.A1(new_n597), .A2(new_n598), .B1(new_n599), .B2(new_n600), .ZN(G303));
  OAI21_X1  g176(.A(G651), .B1(new_n525), .B2(G74), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n517), .A2(G49), .A3(G543), .ZN(new_n603));
  INV_X1    g178(.A(G87), .ZN(new_n604));
  OAI211_X1 g179(.A(new_n602), .B(new_n603), .C1(new_n604), .C2(new_n560), .ZN(G288));
  NAND3_X1  g180(.A1(new_n516), .A2(G61), .A3(new_n502), .ZN(new_n606));
  NAND2_X1  g181(.A1(G73), .A2(G543), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G651), .ZN(new_n609));
  NAND4_X1  g184(.A1(new_n516), .A2(G86), .A3(new_n502), .A4(new_n517), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n517), .A2(G48), .A3(G543), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n609), .A2(new_n613), .ZN(G305));
  INV_X1    g189(.A(G47), .ZN(new_n615));
  INV_X1    g190(.A(G85), .ZN(new_n616));
  OAI22_X1  g191(.A1(new_n534), .A2(new_n615), .B1(new_n616), .B2(new_n560), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n525), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n618), .A2(new_n558), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(new_n620), .ZN(G290));
  NAND2_X1  g196(.A1(G301), .A2(G868), .ZN(new_n622));
  AND3_X1   g197(.A1(new_n525), .A2(G92), .A3(new_n517), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT10), .ZN(new_n624));
  NAND2_X1  g199(.A1(G79), .A2(G543), .ZN(new_n625));
  INV_X1    g200(.A(G66), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n570), .B2(new_n626), .ZN(new_n627));
  AOI22_X1  g202(.A1(new_n627), .A2(G651), .B1(G54), .B2(new_n564), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n622), .B1(new_n630), .B2(G868), .ZN(G284));
  OAI21_X1  g206(.A(new_n622), .B1(new_n630), .B2(G868), .ZN(G321));
  INV_X1    g207(.A(G868), .ZN(new_n633));
  OR3_X1    g208(.A1(G168), .A2(KEYINPUT80), .A3(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(KEYINPUT80), .B1(G168), .B2(new_n633), .ZN(new_n635));
  INV_X1    g210(.A(G299), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n634), .B(new_n635), .C1(G868), .C2(new_n636), .ZN(G297));
  OAI211_X1 g212(.A(new_n634), .B(new_n635), .C1(G868), .C2(new_n636), .ZN(G280));
  XNOR2_X1  g213(.A(KEYINPUT81), .B(G559), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n630), .B1(G860), .B2(new_n639), .ZN(G148));
  NAND2_X1  g215(.A1(new_n630), .A2(new_n639), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(G868), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n642), .B1(G868), .B2(new_n577), .ZN(G323));
  XNOR2_X1  g218(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g219(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n645));
  INV_X1    g220(.A(KEYINPUT82), .ZN(new_n646));
  INV_X1    g221(.A(G111), .ZN(new_n647));
  AOI22_X1  g222(.A1(new_n645), .A2(new_n646), .B1(new_n647), .B2(G2105), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n648), .B1(new_n646), .B2(new_n645), .ZN(new_n649));
  INV_X1    g224(.A(G135), .ZN(new_n650));
  INV_X1    g225(.A(G123), .ZN(new_n651));
  OAI221_X1 g226(.A(new_n649), .B1(new_n480), .B2(new_n650), .C1(new_n651), .C2(new_n483), .ZN(new_n652));
  INV_X1    g227(.A(G2096), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n459), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(KEYINPUT12), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT13), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(G2100), .Z(new_n658));
  NAND2_X1  g233(.A1(new_n654), .A2(new_n658), .ZN(G156));
  XNOR2_X1  g234(.A(G2427), .B(G2438), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2430), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT15), .B(G2435), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n663), .A2(KEYINPUT14), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1341), .B(G1348), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2443), .B(G2446), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n665), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2451), .B(G2454), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n670), .B(new_n671), .Z(new_n672));
  OR2_X1    g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n669), .A2(new_n672), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n673), .A2(G14), .A3(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(G401));
  INV_X1    g251(.A(KEYINPUT18), .ZN(new_n677));
  XOR2_X1   g252(.A(G2084), .B(G2090), .Z(new_n678));
  XNOR2_X1  g253(.A(G2067), .B(G2678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n680), .A2(KEYINPUT17), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n678), .A2(new_n679), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n677), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(G2100), .ZN(new_n684));
  XOR2_X1   g259(.A(G2072), .B(G2078), .Z(new_n685));
  AOI21_X1  g260(.A(new_n685), .B1(new_n680), .B2(KEYINPUT18), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(new_n653), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n684), .B(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(G227));
  XOR2_X1   g264(.A(G1971), .B(G1976), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT19), .ZN(new_n691));
  XOR2_X1   g266(.A(G1956), .B(G2474), .Z(new_n692));
  XOR2_X1   g267(.A(G1961), .B(G1966), .Z(new_n693));
  AND2_X1   g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT20), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n692), .A2(new_n693), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  MUX2_X1   g274(.A(new_n699), .B(new_n698), .S(new_n691), .Z(new_n700));
  NOR2_X1   g275(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1981), .B(G1986), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT84), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n703), .B(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(G1991), .B(G1996), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(G229));
  INV_X1    g283(.A(KEYINPUT91), .ZN(new_n709));
  INV_X1    g284(.A(G16), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G6), .ZN(new_n711));
  INV_X1    g286(.A(G305), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n711), .B1(new_n712), .B2(new_n710), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT89), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT32), .B(G1981), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n714), .B(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n710), .A2(G23), .ZN(new_n718));
  INV_X1    g293(.A(G288), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n718), .B1(new_n719), .B2(new_n710), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT90), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT33), .B(G1976), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT34), .ZN(new_n724));
  NOR2_X1   g299(.A1(G16), .A2(G22), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(G166), .B2(G16), .ZN(new_n726));
  INV_X1    g301(.A(G1971), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND4_X1  g303(.A1(new_n717), .A2(new_n723), .A3(new_n724), .A4(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n710), .A2(G24), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n620), .A2(KEYINPUT87), .ZN(new_n731));
  OAI21_X1  g306(.A(G16), .B1(new_n620), .B2(KEYINPUT87), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT88), .B(G1986), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n733), .B(new_n734), .Z(new_n735));
  OR2_X1    g310(.A1(G25), .A2(G29), .ZN(new_n736));
  OR2_X1    g311(.A1(G95), .A2(G2105), .ZN(new_n737));
  OAI211_X1 g312(.A(new_n737), .B(G2104), .C1(G107), .C2(new_n459), .ZN(new_n738));
  INV_X1    g313(.A(G131), .ZN(new_n739));
  INV_X1    g314(.A(G119), .ZN(new_n740));
  OAI221_X1 g315(.A(new_n738), .B1(new_n480), .B2(new_n739), .C1(new_n740), .C2(new_n483), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT85), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(new_n480), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G131), .ZN(new_n745));
  INV_X1    g320(.A(new_n483), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(G119), .ZN(new_n747));
  NAND4_X1  g322(.A1(new_n745), .A2(new_n747), .A3(KEYINPUT85), .A4(new_n738), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n743), .A2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(G29), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n736), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  XOR2_X1   g326(.A(KEYINPUT35), .B(G1991), .Z(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT86), .Z(new_n753));
  XNOR2_X1  g328(.A(new_n751), .B(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n735), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n709), .B1(new_n729), .B2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  AND2_X1   g332(.A1(KEYINPUT92), .A2(KEYINPUT36), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n729), .A2(new_n755), .A3(new_n709), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n723), .A2(new_n728), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n714), .B(new_n715), .ZN(new_n761));
  OAI21_X1  g336(.A(KEYINPUT34), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND4_X1  g337(.A1(new_n757), .A2(new_n758), .A3(new_n759), .A4(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(G16), .A2(G19), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n577), .B2(G16), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(G1341), .Z(new_n766));
  AND2_X1   g341(.A1(new_n750), .A2(G32), .ZN(new_n767));
  NAND3_X1  g342(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT26), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n768), .A2(new_n769), .ZN(new_n771));
  AND2_X1   g346(.A1(new_n459), .A2(G2104), .ZN(new_n772));
  AOI22_X1  g347(.A1(new_n770), .A2(new_n771), .B1(G105), .B2(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(G141), .ZN(new_n774));
  INV_X1    g349(.A(G129), .ZN(new_n775));
  OAI221_X1 g350(.A(new_n773), .B1(new_n480), .B2(new_n774), .C1(new_n775), .C2(new_n483), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n767), .B1(new_n776), .B2(G29), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT27), .B(G1996), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n766), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n710), .A2(G4), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(new_n630), .B2(new_n710), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G1348), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n750), .A2(G35), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n484), .B2(G29), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT29), .B(G2090), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(G34), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n787), .A2(KEYINPUT24), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n787), .A2(KEYINPUT24), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n750), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G160), .B2(new_n750), .ZN(new_n791));
  INV_X1    g366(.A(G2084), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n750), .A2(G27), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G164), .B2(new_n750), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n795), .A2(G2078), .ZN(new_n796));
  XOR2_X1   g371(.A(KEYINPUT30), .B(G28), .Z(new_n797));
  NOR2_X1   g372(.A1(KEYINPUT31), .A2(G11), .ZN(new_n798));
  AND2_X1   g373(.A1(KEYINPUT31), .A2(G11), .ZN(new_n799));
  OAI221_X1 g374(.A(new_n796), .B1(G29), .B2(new_n797), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  OAI22_X1  g375(.A1(new_n652), .A2(new_n750), .B1(new_n795), .B2(G2078), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n786), .A2(new_n793), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n777), .A2(new_n778), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT95), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NOR4_X1   g381(.A1(new_n779), .A2(new_n782), .A3(new_n803), .A4(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(G115), .A2(G2104), .ZN(new_n808));
  INV_X1    g383(.A(G127), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n808), .B1(new_n493), .B2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT25), .ZN(new_n811));
  NAND2_X1  g386(.A1(G103), .A2(G2104), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n811), .B1(new_n812), .B2(G2105), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n459), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n814));
  AOI22_X1  g389(.A1(new_n810), .A2(G2105), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g390(.A(KEYINPUT94), .B1(new_n744), .B2(G139), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT94), .ZN(new_n817));
  INV_X1    g392(.A(G139), .ZN(new_n818));
  NOR3_X1   g393(.A1(new_n480), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n815), .B1(new_n816), .B2(new_n819), .ZN(new_n820));
  MUX2_X1   g395(.A(G33), .B(new_n820), .S(G29), .Z(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(G2072), .ZN(new_n822));
  XNOR2_X1  g397(.A(KEYINPUT100), .B(KEYINPUT23), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n710), .A2(G20), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(G299), .B2(G16), .ZN(new_n826));
  INV_X1    g401(.A(G1956), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n750), .A2(G26), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(KEYINPUT28), .Z(new_n830));
  NAND2_X1  g405(.A1(new_n744), .A2(G140), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n746), .A2(G128), .ZN(new_n832));
  OR2_X1    g407(.A1(G104), .A2(G2105), .ZN(new_n833));
  OAI211_X1 g408(.A(new_n833), .B(G2104), .C1(G116), .C2(new_n459), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT93), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n831), .A2(new_n832), .A3(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n830), .B1(new_n836), .B2(G29), .ZN(new_n837));
  INV_X1    g412(.A(G2067), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(G5), .A2(G16), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT99), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(G301), .B2(new_n710), .ZN(new_n842));
  INV_X1    g417(.A(G1961), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  NOR4_X1   g419(.A1(new_n822), .A2(new_n828), .A3(new_n839), .A4(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(G1966), .ZN(new_n846));
  NOR3_X1   g421(.A1(G286), .A2(KEYINPUT96), .A3(new_n710), .ZN(new_n847));
  OAI21_X1  g422(.A(KEYINPUT96), .B1(G16), .B2(G21), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(G168), .B2(G16), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT97), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR3_X1   g427(.A1(new_n847), .A2(KEYINPUT97), .A3(new_n849), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n846), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n807), .A2(new_n845), .A3(new_n854), .ZN(new_n855));
  OR3_X1    g430(.A1(new_n852), .A2(new_n846), .A3(new_n853), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(KEYINPUT98), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n856), .A2(KEYINPUT98), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n855), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n759), .ZN(new_n860));
  INV_X1    g435(.A(new_n762), .ZN(new_n861));
  NOR3_X1   g436(.A1(new_n860), .A2(new_n756), .A3(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(KEYINPUT92), .B(KEYINPUT36), .ZN(new_n863));
  OAI211_X1 g438(.A(new_n763), .B(new_n859), .C1(new_n862), .C2(new_n863), .ZN(G150));
  INV_X1    g439(.A(G150), .ZN(G311));
  NAND2_X1  g440(.A1(new_n630), .A2(G559), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT38), .ZN(new_n867));
  INV_X1    g442(.A(G55), .ZN(new_n868));
  INV_X1    g443(.A(G93), .ZN(new_n869));
  OAI22_X1  g444(.A1(new_n534), .A2(new_n868), .B1(new_n869), .B2(new_n560), .ZN(new_n870));
  AOI22_X1  g445(.A1(new_n525), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n871), .A2(new_n558), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(new_n576), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n870), .A2(new_n872), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n577), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n867), .B(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT39), .ZN(new_n879));
  AOI21_X1  g454(.A(G860), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n880), .B1(new_n879), .B2(new_n878), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n873), .A2(G860), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n882), .B(KEYINPUT37), .Z(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(G145));
  NAND2_X1  g459(.A1(new_n836), .A2(new_n499), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n831), .A2(new_n832), .A3(G164), .A4(new_n835), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n885), .A2(new_n776), .A3(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n776), .B1(new_n885), .B2(new_n886), .ZN(new_n889));
  OAI211_X1 g464(.A(KEYINPUT101), .B(new_n820), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n889), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n820), .A2(KEYINPUT101), .ZN(new_n892));
  OR2_X1    g467(.A1(new_n820), .A2(KEYINPUT101), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n891), .A2(new_n892), .A3(new_n893), .A4(new_n887), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n743), .A2(new_n748), .A3(KEYINPUT102), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(KEYINPUT102), .B1(new_n743), .B2(new_n748), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n656), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n744), .A2(G142), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n746), .A2(G130), .ZN(new_n901));
  OR2_X1    g476(.A1(G106), .A2(G2105), .ZN(new_n902));
  OAI211_X1 g477(.A(new_n902), .B(G2104), .C1(G118), .C2(new_n459), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n900), .A2(new_n901), .A3(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT102), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n749), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n656), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n906), .A2(new_n907), .A3(new_n896), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n899), .A2(new_n904), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n904), .B1(new_n899), .B2(new_n908), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n895), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n904), .ZN(new_n913));
  NOR3_X1   g488(.A1(new_n897), .A2(new_n656), .A3(new_n898), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n907), .B1(new_n906), .B2(new_n896), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n916), .A2(new_n909), .A3(new_n890), .A4(new_n894), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n912), .A2(new_n917), .ZN(new_n918));
  XOR2_X1   g493(.A(new_n484), .B(new_n652), .Z(new_n919));
  XNOR2_X1  g494(.A(new_n919), .B(G160), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(G37), .ZN(new_n922));
  INV_X1    g497(.A(new_n920), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n912), .A2(new_n917), .A3(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n921), .A2(new_n922), .A3(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n925), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g501(.A(new_n641), .B(new_n877), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n630), .A2(new_n636), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n629), .A2(G299), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n930), .B(KEYINPUT41), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n931), .B1(new_n932), .B2(new_n927), .ZN(new_n933));
  OR2_X1    g508(.A1(new_n933), .A2(KEYINPUT42), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(KEYINPUT42), .ZN(new_n935));
  NAND2_X1  g510(.A1(G166), .A2(new_n712), .ZN(new_n936));
  NAND2_X1  g511(.A1(G303), .A2(G305), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n620), .B(G288), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT103), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n936), .B(new_n937), .C1(new_n938), .C2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n939), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n940), .B(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n934), .A2(new_n935), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n943), .B1(new_n934), .B2(new_n935), .ZN(new_n945));
  OAI21_X1  g520(.A(G868), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n946), .B1(G868), .B2(new_n875), .ZN(G295));
  OAI21_X1  g522(.A(new_n946), .B1(G868), .B2(new_n875), .ZN(G331));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n949));
  AND2_X1   g524(.A1(new_n928), .A2(new_n929), .ZN(new_n950));
  AOI21_X1  g525(.A(G301), .B1(new_n874), .B2(new_n876), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n874), .A2(new_n876), .A3(G301), .ZN(new_n953));
  AOI21_X1  g528(.A(G168), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n953), .ZN(new_n955));
  NOR3_X1   g530(.A1(new_n955), .A2(G286), .A3(new_n951), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n950), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n950), .A2(KEYINPUT41), .ZN(new_n958));
  OAI21_X1  g533(.A(G286), .B1(new_n955), .B2(new_n951), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n952), .A2(G168), .A3(new_n953), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT41), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n930), .A2(new_n961), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n958), .A2(new_n959), .A3(new_n960), .A4(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n957), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(G37), .B1(new_n964), .B2(new_n943), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT43), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n957), .A2(new_n942), .A3(new_n963), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n966), .B1(new_n965), .B2(new_n967), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n949), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n970), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n972), .A2(KEYINPUT44), .A3(new_n968), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n971), .A2(new_n973), .ZN(G397));
  XNOR2_X1  g549(.A(new_n836), .B(G2067), .ZN(new_n975));
  INV_X1    g550(.A(G1384), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n499), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT45), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G125), .ZN(new_n980));
  OR2_X1    g555(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n981));
  NAND2_X1  g556(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n980), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n470), .ZN(new_n984));
  OAI21_X1  g559(.A(G2105), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n985), .A2(G40), .A3(new_n464), .A4(new_n467), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n979), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n975), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT105), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n988), .B(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n987), .ZN(new_n991));
  INV_X1    g566(.A(new_n776), .ZN(new_n992));
  INV_X1    g567(.A(G1996), .ZN(new_n993));
  NOR3_X1   g568(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n987), .A2(new_n993), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n995), .B(KEYINPUT104), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n994), .B1(new_n996), .B2(new_n992), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n990), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(KEYINPUT106), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT106), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n990), .A2(new_n1000), .A3(new_n997), .ZN(new_n1001));
  INV_X1    g576(.A(new_n752), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n749), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n743), .A2(new_n748), .A3(new_n752), .ZN(new_n1004));
  AND2_X1   g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n999), .B(new_n1001), .C1(new_n991), .C2(new_n1005), .ZN(new_n1006));
  OR2_X1    g581(.A1(G290), .A2(G1986), .ZN(new_n1007));
  NAND2_X1  g582(.A1(G290), .A2(G1986), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n991), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(G8), .ZN(new_n1011));
  INV_X1    g586(.A(G40), .ZN(new_n1012));
  NOR3_X1   g587(.A1(new_n468), .A2(new_n471), .A3(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n499), .A2(KEYINPUT45), .A3(new_n976), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n979), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n846), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n986), .B1(new_n977), .B2(KEYINPUT50), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT50), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n499), .A2(new_n1018), .A3(new_n976), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1017), .A2(new_n792), .A3(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1011), .B1(new_n1016), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(G168), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g598(.A(KEYINPUT108), .B(G2090), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1017), .A2(new_n1024), .A3(new_n1019), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n986), .B1(new_n977), .B2(new_n978), .ZN(new_n1026));
  AOI21_X1  g601(.A(G1971), .B1(new_n1026), .B2(new_n1014), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT107), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1025), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  AND3_X1   g604(.A1(new_n499), .A2(KEYINPUT45), .A3(new_n976), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT45), .B1(new_n499), .B2(new_n976), .ZN(new_n1031));
  NOR3_X1   g606(.A1(new_n1030), .A2(new_n1031), .A3(new_n986), .ZN(new_n1032));
  NOR3_X1   g607(.A1(new_n1032), .A2(KEYINPUT107), .A3(G1971), .ZN(new_n1033));
  OAI21_X1  g608(.A(G8), .B1(new_n1029), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(KEYINPUT115), .ZN(new_n1035));
  AND3_X1   g610(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1036));
  AOI21_X1  g611(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(KEYINPUT107), .B1(new_n1032), .B2(G1971), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1015), .A2(new_n1028), .A3(new_n727), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1039), .A2(new_n1025), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT115), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1041), .A2(new_n1042), .A3(G8), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1035), .A2(new_n1038), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G1976), .ZN(new_n1045));
  NOR2_X1   g620(.A1(G288), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  OAI211_X1 g622(.A(KEYINPUT110), .B(G8), .C1(new_n977), .C2(new_n986), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  NAND4_X1  g624(.A1(G160), .A2(G40), .A3(new_n976), .A4(new_n499), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT110), .B1(new_n1050), .B2(G8), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1047), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(KEYINPUT52), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT49), .ZN(new_n1054));
  INV_X1    g629(.A(G1981), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1055), .B1(new_n609), .B2(new_n613), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n558), .B1(new_n606), .B2(new_n607), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n1057), .A2(new_n612), .A3(G1981), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1054), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT112), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  OR3_X1    g636(.A1(new_n1056), .A2(new_n1058), .A3(new_n1054), .ZN(new_n1062));
  OAI21_X1  g637(.A(G8), .B1(new_n977), .B2(new_n986), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT110), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(new_n1048), .ZN(new_n1066));
  OAI211_X1 g641(.A(KEYINPUT112), .B(new_n1054), .C1(new_n1056), .C2(new_n1058), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1061), .A2(new_n1062), .A3(new_n1066), .A4(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(KEYINPUT52), .B1(G288), .B2(new_n1045), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n1047), .B(new_n1069), .C1(new_n1049), .C2(new_n1051), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1070), .A2(KEYINPUT111), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT111), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1046), .B1(new_n1065), .B2(new_n1048), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1072), .B1(new_n1073), .B2(new_n1069), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1053), .B(new_n1068), .C1(new_n1071), .C2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1075), .A2(KEYINPUT113), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT113), .ZN(new_n1077));
  AND2_X1   g652(.A1(new_n1068), .A2(new_n1053), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1070), .A2(KEYINPUT111), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1073), .A2(new_n1072), .A3(new_n1069), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1077), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1023), .B(new_n1044), .C1(new_n1076), .C2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT63), .ZN(new_n1084));
  NOR2_X1   g659(.A1(G288), .A2(G1976), .ZN(new_n1085));
  XNOR2_X1  g660(.A(new_n1085), .B(KEYINPUT114), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1058), .B1(new_n1068), .B2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1087), .B1(new_n1048), .B2(new_n1065), .ZN(new_n1088));
  XNOR2_X1  g663(.A(new_n1075), .B(KEYINPUT113), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT109), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1090), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT55), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1092), .B1(G166), .B2(new_n1011), .ZN(new_n1093));
  NAND3_X1  g668(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1093), .A2(KEYINPUT109), .A3(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1041), .A2(new_n1091), .A3(G8), .A4(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1088), .B1(new_n1089), .B2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1022), .A2(KEYINPUT63), .ZN(new_n1099));
  INV_X1    g674(.A(G2078), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n979), .A2(new_n1100), .A3(new_n1013), .A4(new_n1014), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT53), .ZN(new_n1102));
  AND3_X1   g677(.A1(new_n1101), .A2(KEYINPUT123), .A3(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT123), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n843), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1107), .B1(new_n1102), .B2(new_n1101), .ZN(new_n1108));
  OAI21_X1  g683(.A(G171), .B1(new_n1105), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1016), .A2(new_n1020), .ZN(new_n1110));
  AOI21_X1  g685(.A(KEYINPUT121), .B1(G286), .B2(G8), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT121), .ZN(new_n1112));
  NOR3_X1   g687(.A1(G168), .A2(new_n1112), .A3(new_n1011), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1110), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT122), .ZN(new_n1115));
  NAND3_X1  g690(.A1(G286), .A2(KEYINPUT121), .A3(G8), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1112), .B1(G168), .B2(new_n1011), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT122), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1118), .A2(new_n1119), .A3(new_n1110), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1115), .A2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(KEYINPUT51), .B1(new_n1118), .B2(new_n1021), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n1017), .A2(new_n792), .A3(new_n1019), .ZN(new_n1123));
  AOI21_X1  g698(.A(G1966), .B1(new_n1026), .B2(new_n1014), .ZN(new_n1124));
  OAI21_X1  g699(.A(G8), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT51), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1125), .A2(new_n1126), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1122), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1121), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1109), .B1(new_n1129), .B2(KEYINPUT62), .ZN(new_n1130));
  AOI22_X1  g705(.A1(new_n1115), .A2(new_n1120), .B1(new_n1122), .B2(new_n1127), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT62), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1099), .B1(new_n1130), .B2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1025), .B1(new_n1032), .B2(G1971), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(G8), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(new_n1038), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1078), .A2(new_n1096), .A3(new_n1081), .A4(new_n1137), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1084), .B(new_n1098), .C1(new_n1134), .C2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1091), .A2(new_n1095), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1137), .B1(new_n1140), .B2(new_n1034), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1141), .A2(new_n1075), .ZN(new_n1142));
  OAI21_X1  g717(.A(KEYINPUT54), .B1(G301), .B2(KEYINPUT124), .ZN(new_n1143));
  NOR4_X1   g718(.A1(new_n1030), .A2(new_n1031), .A3(G2078), .A4(new_n986), .ZN(new_n1144));
  AOI22_X1  g719(.A1(new_n1144), .A2(KEYINPUT53), .B1(new_n843), .B2(new_n1106), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n1145), .B(G301), .C1(new_n1104), .C2(new_n1103), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT123), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1101), .A2(KEYINPUT123), .A3(new_n1102), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(G301), .B1(new_n1152), .B2(new_n1145), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1143), .B1(new_n1147), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1143), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1109), .A2(new_n1146), .A3(new_n1155), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1142), .A2(new_n1154), .A3(new_n1129), .A4(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT125), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  AND3_X1   g734(.A1(new_n1109), .A2(new_n1146), .A3(new_n1155), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1155), .B1(new_n1109), .B2(new_n1146), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1131), .A2(new_n1138), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1162), .A2(new_n1163), .A3(KEYINPUT125), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1013), .A2(new_n976), .A3(new_n838), .A4(new_n499), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n1165), .B(KEYINPUT118), .ZN(new_n1166));
  AOI21_X1  g741(.A(G1348), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1167));
  NOR4_X1   g742(.A1(new_n1166), .A2(new_n629), .A3(new_n1167), .A4(KEYINPUT60), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT60), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1169), .B1(new_n1170), .B2(new_n630), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n629), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1168), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g748(.A(KEYINPUT56), .B(G2072), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1032), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1106), .A2(new_n827), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1177), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n584), .A2(new_n588), .A3(KEYINPUT116), .A4(new_n592), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT57), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n1181), .B(new_n636), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1178), .A2(new_n1182), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1181), .B(G299), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1184), .A2(new_n1177), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1183), .A2(new_n1185), .A3(KEYINPUT61), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1032), .A2(KEYINPUT119), .A3(new_n993), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT119), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1188), .B1(new_n1015), .B2(G1996), .ZN(new_n1189));
  XOR2_X1   g764(.A(KEYINPUT58), .B(G1341), .Z(new_n1190));
  NAND2_X1  g765(.A1(new_n1050), .A2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1187), .A2(new_n1189), .A3(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1192), .A2(new_n577), .ZN(new_n1193));
  XNOR2_X1  g768(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(new_n1194), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1192), .A2(new_n577), .A3(new_n1196), .ZN(new_n1197));
  NAND4_X1  g772(.A1(new_n1173), .A2(new_n1186), .A3(new_n1195), .A4(new_n1197), .ZN(new_n1198));
  OAI21_X1  g773(.A(KEYINPUT117), .B1(new_n1184), .B2(new_n1177), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT117), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1178), .A2(new_n1182), .A3(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g777(.A(KEYINPUT61), .B1(new_n1202), .B2(new_n1185), .ZN(new_n1203));
  INV_X1    g778(.A(new_n1202), .ZN(new_n1204));
  NOR2_X1   g779(.A1(new_n1170), .A2(new_n629), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1205), .B1(new_n1184), .B2(new_n1177), .ZN(new_n1206));
  OAI22_X1  g781(.A1(new_n1198), .A2(new_n1203), .B1(new_n1204), .B2(new_n1206), .ZN(new_n1207));
  AND3_X1   g782(.A1(new_n1159), .A2(new_n1164), .A3(new_n1207), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n1010), .B1(new_n1139), .B2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n987), .B1(new_n975), .B2(new_n776), .ZN(new_n1210));
  INV_X1    g785(.A(new_n996), .ZN(new_n1211));
  AND2_X1   g786(.A1(new_n1211), .A2(KEYINPUT46), .ZN(new_n1212));
  NOR2_X1   g787(.A1(new_n1211), .A2(KEYINPUT46), .ZN(new_n1213));
  OAI21_X1  g788(.A(new_n1210), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  XNOR2_X1  g789(.A(new_n1214), .B(KEYINPUT47), .ZN(new_n1215));
  NOR2_X1   g790(.A1(new_n1007), .A2(new_n991), .ZN(new_n1216));
  XNOR2_X1  g791(.A(new_n1216), .B(KEYINPUT48), .ZN(new_n1217));
  OAI21_X1  g792(.A(new_n1215), .B1(new_n1006), .B2(new_n1217), .ZN(new_n1218));
  XOR2_X1   g793(.A(new_n1004), .B(KEYINPUT126), .Z(new_n1219));
  NAND3_X1  g794(.A1(new_n999), .A2(new_n1001), .A3(new_n1219), .ZN(new_n1220));
  OR2_X1    g795(.A1(new_n836), .A2(G2067), .ZN(new_n1221));
  AOI21_X1  g796(.A(new_n991), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  NOR2_X1   g797(.A1(new_n1218), .A2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1209), .A2(new_n1223), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g799(.A1(new_n688), .A2(G319), .ZN(new_n1226));
  XOR2_X1   g800(.A(new_n1226), .B(KEYINPUT127), .Z(new_n1227));
  NAND2_X1  g801(.A1(new_n1227), .A2(new_n675), .ZN(new_n1228));
  NOR2_X1   g802(.A1(G229), .A2(new_n1228), .ZN(new_n1229));
  OAI211_X1 g803(.A(new_n925), .B(new_n1229), .C1(new_n969), .C2(new_n970), .ZN(G225));
  INV_X1    g804(.A(G225), .ZN(G308));
endmodule


