

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779;

  OR2_X1 U374 ( .A1(n559), .A2(n417), .ZN(n499) );
  XNOR2_X1 U375 ( .A(n493), .B(n766), .ZN(n743) );
  XNOR2_X1 U376 ( .A(n485), .B(n484), .ZN(n415) );
  NAND2_X1 U377 ( .A1(n774), .A2(G234), .ZN(n485) );
  INV_X1 U378 ( .A(KEYINPUT64), .ZN(n461) );
  NAND2_X1 U379 ( .A1(n349), .A2(n574), .ZN(n575) );
  NOR2_X1 U380 ( .A1(n368), .A2(n649), .ZN(n349) );
  AND2_X2 U381 ( .A1(n438), .A2(n637), .ZN(n406) );
  AND2_X2 U382 ( .A1(n550), .A2(n549), .ZN(n571) );
  XNOR2_X2 U383 ( .A(n435), .B(n434), .ZN(n722) );
  NOR2_X2 U384 ( .A1(n387), .A2(n711), .ZN(n435) );
  NOR2_X2 U385 ( .A1(n562), .A2(n548), .ZN(n665) );
  XNOR2_X2 U386 ( .A(n579), .B(n578), .ZN(n748) );
  INV_X1 U387 ( .A(n540), .ZN(n542) );
  NAND2_X1 U388 ( .A1(n391), .A2(n390), .ZN(n389) );
  INV_X1 U389 ( .A(n748), .ZN(n750) );
  OR2_X1 U390 ( .A1(n607), .A2(n606), .ZN(n608) );
  BUF_X1 U391 ( .A(n551), .Z(n562) );
  AND2_X1 U392 ( .A1(n400), .A2(n398), .ZN(n375) );
  XNOR2_X1 U393 ( .A(n595), .B(KEYINPUT39), .ZN(n400) );
  NAND2_X1 U394 ( .A1(n542), .A2(n442), .ZN(n441) );
  AND2_X1 U395 ( .A1(n594), .A2(n593), .ZN(n602) );
  OR2_X1 U396 ( .A1(n612), .A2(n418), .ZN(n553) );
  INV_X1 U397 ( .A(n385), .ZN(n580) );
  OR2_X1 U398 ( .A1(n696), .A2(n623), .ZN(n592) );
  XNOR2_X1 U399 ( .A(n653), .B(KEYINPUT62), .ZN(n654) );
  XNOR2_X1 U400 ( .A(n452), .B(KEYINPUT3), .ZN(n454) );
  XNOR2_X1 U401 ( .A(n508), .B(n440), .ZN(n439) );
  INV_X1 U402 ( .A(KEYINPUT69), .ZN(n452) );
  XNOR2_X1 U403 ( .A(G119), .B(G116), .ZN(n453) );
  XNOR2_X1 U404 ( .A(KEYINPUT71), .B(KEYINPUT34), .ZN(n565) );
  XNOR2_X1 U405 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n487) );
  BUF_X1 U406 ( .A(n611), .Z(n350) );
  NOR2_X2 U407 ( .A1(n779), .A2(n649), .ZN(n410) );
  XNOR2_X2 U408 ( .A(n558), .B(n557), .ZN(n779) );
  NOR2_X2 U409 ( .A1(n562), .A2(n561), .ZN(n649) );
  INV_X1 U410 ( .A(n437), .ZN(n351) );
  BUF_X1 U411 ( .A(n709), .Z(n352) );
  XNOR2_X1 U412 ( .A(n580), .B(KEYINPUT38), .ZN(n709) );
  NAND2_X1 U413 ( .A1(n392), .A2(n360), .ZN(n391) );
  NAND2_X1 U414 ( .A1(n405), .A2(n406), .ZN(n392) );
  XNOR2_X1 U415 ( .A(n581), .B(n436), .ZN(n387) );
  XNOR2_X2 U416 ( .A(n457), .B(n456), .ZN(n755) );
  INV_X1 U417 ( .A(KEYINPUT33), .ZN(n563) );
  NOR2_X1 U418 ( .A1(n634), .A2(n404), .ZN(n403) );
  INV_X1 U419 ( .A(n637), .ZN(n404) );
  INV_X1 U420 ( .A(KEYINPUT44), .ZN(n430) );
  AND2_X1 U421 ( .A1(n433), .A2(n410), .ZN(n376) );
  INV_X1 U422 ( .A(G237), .ZN(n467) );
  XOR2_X1 U423 ( .A(KEYINPUT68), .B(G131), .Z(n520) );
  NOR2_X1 U424 ( .A1(G953), .A2(G237), .ZN(n523) );
  XNOR2_X1 U425 ( .A(G140), .B(G110), .ZN(n502) );
  XOR2_X1 U426 ( .A(G146), .B(G125), .Z(n482) );
  INV_X1 U427 ( .A(KEYINPUT6), .ZN(n411) );
  INV_X1 U428 ( .A(KEYINPUT48), .ZN(n420) );
  INV_X1 U429 ( .A(KEYINPUT41), .ZN(n434) );
  BUF_X1 U430 ( .A(n580), .Z(n408) );
  INV_X1 U431 ( .A(KEYINPUT28), .ZN(n395) );
  NAND2_X1 U432 ( .A1(n689), .A2(n358), .ZN(n396) );
  INV_X1 U433 ( .A(n412), .ZN(n612) );
  NAND2_X1 U434 ( .A1(n772), .A2(n634), .ZN(n438) );
  INV_X1 U435 ( .A(KEYINPUT86), .ZN(n373) );
  NAND2_X1 U436 ( .A1(n431), .A2(n428), .ZN(n422) );
  XNOR2_X1 U437 ( .A(KEYINPUT15), .B(G902), .ZN(n636) );
  NOR2_X1 U438 ( .A1(n711), .A2(n417), .ZN(n541) );
  XNOR2_X1 U439 ( .A(G137), .B(G134), .ZN(n471) );
  XOR2_X1 U440 ( .A(KEYINPUT18), .B(KEYINPUT81), .Z(n463) );
  XNOR2_X1 U441 ( .A(KEYINPUT66), .B(G101), .ZN(n460) );
  NAND2_X1 U442 ( .A1(G234), .A2(G237), .ZN(n444) );
  INV_X1 U443 ( .A(KEYINPUT107), .ZN(n436) );
  INV_X1 U444 ( .A(G902), .ZN(n531) );
  INV_X1 U445 ( .A(KEYINPUT1), .ZN(n382) );
  XNOR2_X1 U446 ( .A(KEYINPUT5), .B(G113), .ZN(n473) );
  XNOR2_X1 U447 ( .A(n477), .B(n455), .ZN(n457) );
  XOR2_X1 U448 ( .A(G110), .B(KEYINPUT16), .Z(n455) );
  XNOR2_X1 U449 ( .A(n483), .B(KEYINPUT10), .ZN(n766) );
  INV_X1 U450 ( .A(KEYINPUT8), .ZN(n484) );
  XNOR2_X1 U451 ( .A(G116), .B(G134), .ZN(n512) );
  XNOR2_X1 U452 ( .A(G107), .B(G104), .ZN(n503) );
  INV_X1 U453 ( .A(KEYINPUT31), .ZN(n440) );
  XOR2_X1 U454 ( .A(n658), .B(KEYINPUT59), .Z(n659) );
  NAND2_X1 U455 ( .A1(n750), .A2(n437), .ZN(n687) );
  NAND2_X1 U456 ( .A1(n629), .A2(n408), .ZN(n686) );
  XNOR2_X1 U457 ( .A(n388), .B(n365), .ZN(n778) );
  INV_X1 U458 ( .A(n682), .ZN(n399) );
  NOR2_X1 U459 ( .A1(n600), .A2(n408), .ZN(n601) );
  NAND2_X1 U460 ( .A1(n356), .A2(n605), .ZN(n676) );
  AND2_X1 U461 ( .A1(n363), .A2(n696), .ZN(n353) );
  INV_X1 U462 ( .A(n694), .ZN(n417) );
  OR2_X1 U463 ( .A1(n587), .A2(n586), .ZN(n354) );
  XOR2_X1 U464 ( .A(n505), .B(n504), .Z(n355) );
  AND2_X1 U465 ( .A1(n394), .A2(n370), .ZN(n356) );
  XOR2_X1 U466 ( .A(n464), .B(KEYINPUT17), .Z(n357) );
  AND2_X1 U467 ( .A1(n588), .A2(n694), .ZN(n358) );
  AND2_X1 U468 ( .A1(n370), .A2(n354), .ZN(n359) );
  NAND2_X1 U469 ( .A1(n371), .A2(n372), .ZN(n360) );
  XOR2_X1 U470 ( .A(n495), .B(KEYINPUT25), .Z(n361) );
  AND2_X1 U471 ( .A1(n648), .A2(n686), .ZN(n362) );
  AND2_X1 U472 ( .A1(n691), .A2(n370), .ZN(n363) );
  NOR2_X1 U473 ( .A1(n712), .A2(n387), .ZN(n364) );
  XOR2_X1 U474 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n365) );
  XOR2_X1 U475 ( .A(n641), .B(n640), .Z(n366) );
  OR2_X1 U476 ( .A1(n568), .A2(n536), .ZN(n679) );
  INV_X1 U477 ( .A(n679), .ZN(n398) );
  NAND2_X1 U478 ( .A1(n572), .A2(KEYINPUT44), .ZN(n367) );
  XNOR2_X1 U479 ( .A(n575), .B(KEYINPUT70), .ZN(n576) );
  XNOR2_X1 U480 ( .A(n570), .B(KEYINPUT35), .ZN(n368) );
  XNOR2_X1 U481 ( .A(n389), .B(KEYINPUT65), .ZN(n369) );
  XNOR2_X1 U482 ( .A(n506), .B(G469), .ZN(n370) );
  XNOR2_X1 U483 ( .A(n570), .B(KEYINPUT35), .ZN(n650) );
  XNOR2_X1 U484 ( .A(n389), .B(KEYINPUT65), .ZN(n738) );
  XNOR2_X1 U485 ( .A(n506), .B(G469), .ZN(n589) );
  NAND2_X1 U486 ( .A1(n772), .A2(n374), .ZN(n371) );
  OR2_X1 U487 ( .A1(n373), .A2(n403), .ZN(n372) );
  AND2_X1 U488 ( .A1(n634), .A2(KEYINPUT86), .ZN(n374) );
  NAND2_X1 U489 ( .A1(n433), .A2(n410), .ZN(n432) );
  XNOR2_X1 U490 ( .A(n611), .B(KEYINPUT19), .ZN(n605) );
  NAND2_X1 U491 ( .A1(n385), .A2(n708), .ZN(n611) );
  NAND2_X1 U492 ( .A1(n400), .A2(n398), .ZN(n377) );
  NAND2_X1 U493 ( .A1(n377), .A2(n597), .ZN(n379) );
  NAND2_X1 U494 ( .A1(n375), .A2(n378), .ZN(n380) );
  NAND2_X1 U495 ( .A1(n380), .A2(n379), .ZN(n652) );
  INV_X1 U496 ( .A(n597), .ZN(n378) );
  BUF_X1 U497 ( .A(n559), .Z(n416) );
  XNOR2_X1 U498 ( .A(n696), .B(n411), .ZN(n412) );
  NAND2_X1 U499 ( .A1(n589), .A2(KEYINPUT1), .ZN(n383) );
  NAND2_X1 U500 ( .A1(n381), .A2(n382), .ZN(n384) );
  NAND2_X1 U501 ( .A1(n384), .A2(n383), .ZN(n546) );
  INV_X1 U502 ( .A(n589), .ZN(n381) );
  XNOR2_X2 U503 ( .A(n414), .B(n468), .ZN(n385) );
  NAND2_X1 U504 ( .A1(n653), .A2(n531), .ZN(n401) );
  XNOR2_X1 U505 ( .A(n393), .B(n355), .ZN(n734) );
  XNOR2_X1 U506 ( .A(n413), .B(n507), .ZN(n386) );
  XNOR2_X1 U507 ( .A(n413), .B(n507), .ZN(n688) );
  BUF_X1 U508 ( .A(n546), .Z(n692) );
  XNOR2_X1 U509 ( .A(n466), .B(n465), .ZN(n638) );
  NOR2_X2 U510 ( .A1(n778), .A2(n652), .ZN(n598) );
  NAND2_X1 U511 ( .A1(n722), .A2(n356), .ZN(n388) );
  NAND2_X1 U512 ( .A1(n750), .A2(n407), .ZN(n390) );
  XNOR2_X1 U513 ( .A(n393), .B(n479), .ZN(n653) );
  XNOR2_X2 U514 ( .A(n402), .B(n472), .ZN(n393) );
  XNOR2_X2 U515 ( .A(n765), .B(n460), .ZN(n402) );
  XNOR2_X2 U516 ( .A(n515), .B(KEYINPUT4), .ZN(n765) );
  XNOR2_X1 U517 ( .A(n396), .B(n395), .ZN(n394) );
  NAND2_X1 U518 ( .A1(n707), .A2(n397), .ZN(n566) );
  NAND2_X1 U519 ( .A1(n397), .A2(n353), .ZN(n668) );
  XNOR2_X1 U520 ( .A(n540), .B(KEYINPUT93), .ZN(n397) );
  NAND2_X1 U521 ( .A1(n400), .A2(n399), .ZN(n648) );
  XNOR2_X2 U522 ( .A(n401), .B(n481), .ZN(n696) );
  XNOR2_X1 U523 ( .A(n755), .B(n402), .ZN(n466) );
  INV_X1 U524 ( .A(n748), .ZN(n405) );
  INV_X1 U525 ( .A(n772), .ZN(n437) );
  NOR2_X1 U526 ( .A1(n772), .A2(n631), .ZN(n407) );
  XNOR2_X1 U527 ( .A(n421), .B(n420), .ZN(n419) );
  BUF_X2 U528 ( .A(n369), .Z(n742) );
  XNOR2_X2 U529 ( .A(n409), .B(KEYINPUT0), .ZN(n540) );
  NAND2_X1 U530 ( .A1(n605), .A2(n470), .ZN(n409) );
  NAND2_X1 U531 ( .A1(n546), .A2(n691), .ZN(n413) );
  NOR2_X2 U532 ( .A1(n688), .A2(n412), .ZN(n564) );
  NAND2_X1 U533 ( .A1(n638), .A2(n636), .ZN(n414) );
  NAND2_X1 U534 ( .A1(n415), .A2(G221), .ZN(n492) );
  NAND2_X1 U535 ( .A1(n415), .A2(G217), .ZN(n510) );
  XNOR2_X1 U536 ( .A(n496), .B(n361), .ZN(n559) );
  AND2_X1 U537 ( .A1(n416), .A2(n354), .ZN(n588) );
  AND2_X1 U538 ( .A1(n416), .A2(n417), .ZN(n695) );
  INV_X1 U539 ( .A(n416), .ZN(n418) );
  NAND2_X2 U540 ( .A1(n419), .A2(n362), .ZN(n772) );
  NAND2_X1 U541 ( .A1(n622), .A2(n621), .ZN(n421) );
  NAND2_X1 U542 ( .A1(n691), .A2(n359), .ZN(n590) );
  NAND2_X1 U543 ( .A1(n376), .A2(n427), .ZN(n425) );
  NAND2_X1 U544 ( .A1(n423), .A2(n422), .ZN(n577) );
  NAND2_X1 U545 ( .A1(n425), .A2(n424), .ZN(n423) );
  NAND2_X1 U546 ( .A1(n432), .A2(n367), .ZN(n424) );
  NAND2_X1 U547 ( .A1(n426), .A2(KEYINPUT88), .ZN(n431) );
  INV_X1 U548 ( .A(n571), .ZN(n426) );
  NAND2_X1 U549 ( .A1(n571), .A2(KEYINPUT88), .ZN(n427) );
  NAND2_X1 U550 ( .A1(n571), .A2(n429), .ZN(n428) );
  NAND2_X1 U551 ( .A1(KEYINPUT88), .A2(n430), .ZN(n429) );
  INV_X1 U552 ( .A(n650), .ZN(n433) );
  XNOR2_X2 U553 ( .A(n441), .B(n439), .ZN(n681) );
  NOR2_X1 U554 ( .A1(n386), .A2(n696), .ZN(n442) );
  NAND2_X1 U555 ( .A1(n542), .A2(n541), .ZN(n545) );
  OR2_X1 U556 ( .A1(n774), .A2(G952), .ZN(n661) );
  XOR2_X1 U557 ( .A(n491), .B(n490), .Z(n443) );
  BUF_X1 U558 ( .A(n638), .Z(n639) );
  INV_X1 U559 ( .A(n616), .ZN(n552) );
  NOR2_X1 U560 ( .A1(n553), .A2(n552), .ZN(n554) );
  INV_X1 U561 ( .A(KEYINPUT56), .ZN(n644) );
  XOR2_X1 U562 ( .A(KEYINPUT91), .B(KEYINPUT14), .Z(n445) );
  XNOR2_X1 U563 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U564 ( .A(KEYINPUT76), .B(n446), .ZN(n448) );
  NAND2_X1 U565 ( .A1(n448), .A2(G952), .ZN(n447) );
  XNOR2_X1 U566 ( .A(n447), .B(KEYINPUT92), .ZN(n721) );
  NOR2_X1 U567 ( .A1(G953), .A2(n721), .ZN(n587) );
  INV_X1 U568 ( .A(n587), .ZN(n451) );
  NAND2_X1 U569 ( .A1(G902), .A2(n448), .ZN(n582) );
  INV_X1 U570 ( .A(n582), .ZN(n449) );
  INV_X1 U571 ( .A(G953), .ZN(n749) );
  NOR2_X1 U572 ( .A1(G898), .A2(n749), .ZN(n759) );
  NAND2_X1 U573 ( .A1(n449), .A2(n759), .ZN(n450) );
  NAND2_X1 U574 ( .A1(n451), .A2(n450), .ZN(n470) );
  XNOR2_X2 U575 ( .A(n454), .B(n453), .ZN(n477) );
  XOR2_X1 U576 ( .A(G113), .B(G104), .Z(n527) );
  XOR2_X1 U577 ( .A(G122), .B(G107), .Z(n509) );
  XNOR2_X1 U578 ( .A(n527), .B(n509), .ZN(n456) );
  XNOR2_X2 U579 ( .A(G143), .B(KEYINPUT83), .ZN(n459) );
  INV_X1 U580 ( .A(G128), .ZN(n458) );
  XNOR2_X2 U581 ( .A(n459), .B(n458), .ZN(n515) );
  XNOR2_X2 U582 ( .A(n461), .B(G953), .ZN(n774) );
  NAND2_X1 U583 ( .A1(G224), .A2(n774), .ZN(n462) );
  XNOR2_X1 U584 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U585 ( .A(n357), .B(n482), .ZN(n465) );
  NAND2_X1 U586 ( .A1(n531), .A2(n467), .ZN(n469) );
  AND2_X1 U587 ( .A1(n469), .A2(G210), .ZN(n468) );
  NAND2_X1 U588 ( .A1(n469), .A2(G214), .ZN(n708) );
  INV_X1 U589 ( .A(n708), .ZN(n623) );
  XNOR2_X1 U590 ( .A(n520), .B(n471), .ZN(n767) );
  XNOR2_X1 U591 ( .A(n767), .B(G146), .ZN(n472) );
  NAND2_X1 U592 ( .A1(n523), .A2(G210), .ZN(n474) );
  XNOR2_X1 U593 ( .A(n474), .B(n473), .ZN(n476) );
  XNOR2_X1 U594 ( .A(KEYINPUT78), .B(KEYINPUT96), .ZN(n475) );
  XNOR2_X1 U595 ( .A(n476), .B(n475), .ZN(n478) );
  XNOR2_X1 U596 ( .A(n477), .B(n478), .ZN(n479) );
  INV_X1 U597 ( .A(KEYINPUT72), .ZN(n480) );
  XNOR2_X1 U598 ( .A(n480), .B(G472), .ZN(n481) );
  INV_X1 U599 ( .A(n696), .ZN(n689) );
  XNOR2_X1 U600 ( .A(n482), .B(G140), .ZN(n483) );
  XNOR2_X1 U601 ( .A(G119), .B(G110), .ZN(n486) );
  XNOR2_X1 U602 ( .A(n486), .B(KEYINPUT95), .ZN(n491) );
  INV_X1 U603 ( .A(n487), .ZN(n489) );
  XNOR2_X1 U604 ( .A(G128), .B(G137), .ZN(n488) );
  XNOR2_X1 U605 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U606 ( .A(n492), .B(n443), .ZN(n493) );
  NOR2_X1 U607 ( .A1(G902), .A2(n743), .ZN(n496) );
  NAND2_X1 U608 ( .A1(G234), .A2(n636), .ZN(n494) );
  XNOR2_X1 U609 ( .A(KEYINPUT20), .B(n494), .ZN(n497) );
  NAND2_X1 U610 ( .A1(G217), .A2(n497), .ZN(n495) );
  NAND2_X1 U611 ( .A1(n497), .A2(G221), .ZN(n498) );
  XOR2_X1 U612 ( .A(KEYINPUT21), .B(n498), .Z(n694) );
  XNOR2_X2 U613 ( .A(n499), .B(KEYINPUT67), .ZN(n691) );
  NAND2_X1 U614 ( .A1(n774), .A2(G227), .ZN(n501) );
  XNOR2_X1 U615 ( .A(KEYINPUT80), .B(KEYINPUT94), .ZN(n500) );
  XNOR2_X1 U616 ( .A(n501), .B(n500), .ZN(n505) );
  XNOR2_X1 U617 ( .A(n503), .B(n502), .ZN(n504) );
  NAND2_X1 U618 ( .A1(n734), .A2(n531), .ZN(n506) );
  INV_X1 U619 ( .A(KEYINPUT77), .ZN(n507) );
  INV_X1 U620 ( .A(KEYINPUT97), .ZN(n508) );
  NAND2_X1 U621 ( .A1(n681), .A2(n668), .ZN(n538) );
  XOR2_X1 U622 ( .A(n509), .B(KEYINPUT102), .Z(n511) );
  XNOR2_X1 U623 ( .A(n511), .B(n510), .ZN(n517) );
  XOR2_X1 U624 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n513) );
  XNOR2_X1 U625 ( .A(n513), .B(n512), .ZN(n514) );
  XOR2_X1 U626 ( .A(n515), .B(n514), .Z(n516) );
  XNOR2_X1 U627 ( .A(n517), .B(n516), .ZN(n739) );
  NOR2_X1 U628 ( .A1(G902), .A2(n739), .ZN(n518) );
  XNOR2_X1 U629 ( .A(n518), .B(KEYINPUT103), .ZN(n519) );
  XNOR2_X1 U630 ( .A(n519), .B(G478), .ZN(n568) );
  XNOR2_X1 U631 ( .A(G143), .B(n520), .ZN(n521) );
  XNOR2_X1 U632 ( .A(n521), .B(G122), .ZN(n522) );
  XNOR2_X1 U633 ( .A(n766), .B(n522), .ZN(n530) );
  XOR2_X1 U634 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n525) );
  NAND2_X1 U635 ( .A1(G214), .A2(n523), .ZN(n524) );
  XNOR2_X1 U636 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U637 ( .A(KEYINPUT98), .B(n526), .ZN(n528) );
  XNOR2_X1 U638 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U639 ( .A(n530), .B(n529), .ZN(n658) );
  NAND2_X1 U640 ( .A1(n658), .A2(n531), .ZN(n535) );
  XOR2_X1 U641 ( .A(KEYINPUT13), .B(KEYINPUT100), .Z(n533) );
  XNOR2_X1 U642 ( .A(KEYINPUT99), .B(G475), .ZN(n532) );
  XOR2_X1 U643 ( .A(n533), .B(n532), .Z(n534) );
  XNOR2_X1 U644 ( .A(n535), .B(n534), .ZN(n567) );
  XNOR2_X1 U645 ( .A(n567), .B(KEYINPUT101), .ZN(n536) );
  NAND2_X1 U646 ( .A1(n536), .A2(n568), .ZN(n682) );
  AND2_X1 U647 ( .A1(n679), .A2(n682), .ZN(n712) );
  INV_X1 U648 ( .A(n712), .ZN(n537) );
  NAND2_X1 U649 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U650 ( .A(n539), .B(KEYINPUT104), .ZN(n550) );
  OR2_X1 U651 ( .A1(n568), .A2(n567), .ZN(n711) );
  XOR2_X1 U652 ( .A(KEYINPUT73), .B(KEYINPUT74), .Z(n543) );
  XNOR2_X1 U653 ( .A(KEYINPUT22), .B(n543), .ZN(n544) );
  XNOR2_X1 U654 ( .A(n545), .B(n544), .ZN(n551) );
  OR2_X1 U655 ( .A1(n692), .A2(n416), .ZN(n547) );
  OR2_X1 U656 ( .A1(n547), .A2(n612), .ZN(n548) );
  INV_X1 U657 ( .A(n665), .ZN(n549) );
  INV_X1 U658 ( .A(n551), .ZN(n555) );
  XNOR2_X1 U659 ( .A(n692), .B(KEYINPUT90), .ZN(n616) );
  NAND2_X1 U660 ( .A1(n555), .A2(n554), .ZN(n558) );
  INV_X1 U661 ( .A(KEYINPUT82), .ZN(n556) );
  XNOR2_X1 U662 ( .A(n556), .B(KEYINPUT32), .ZN(n557) );
  NAND2_X1 U663 ( .A1(n416), .A2(n696), .ZN(n560) );
  OR2_X1 U664 ( .A1(n692), .A2(n560), .ZN(n561) );
  XNOR2_X1 U665 ( .A(n564), .B(n563), .ZN(n707) );
  XNOR2_X1 U666 ( .A(n566), .B(n565), .ZN(n569) );
  AND2_X1 U667 ( .A1(n568), .A2(n567), .ZN(n599) );
  NAND2_X1 U668 ( .A1(n569), .A2(n599), .ZN(n570) );
  INV_X1 U669 ( .A(KEYINPUT88), .ZN(n572) );
  NOR2_X1 U670 ( .A1(n779), .A2(KEYINPUT44), .ZN(n574) );
  NAND2_X1 U671 ( .A1(n577), .A2(n576), .ZN(n579) );
  INV_X1 U672 ( .A(KEYINPUT45), .ZN(n578) );
  NAND2_X1 U673 ( .A1(n708), .A2(n709), .ZN(n581) );
  NOR2_X1 U674 ( .A1(G900), .A2(n582), .ZN(n584) );
  INV_X1 U675 ( .A(n774), .ZN(n583) );
  NAND2_X1 U676 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U677 ( .A(KEYINPUT105), .B(n585), .ZN(n586) );
  XNOR2_X1 U678 ( .A(n590), .B(KEYINPUT79), .ZN(n594) );
  INV_X1 U679 ( .A(KEYINPUT30), .ZN(n591) );
  XNOR2_X1 U680 ( .A(n592), .B(n591), .ZN(n593) );
  NAND2_X1 U681 ( .A1(n602), .A2(n352), .ZN(n595) );
  INV_X1 U682 ( .A(KEYINPUT106), .ZN(n596) );
  XNOR2_X1 U683 ( .A(n596), .B(KEYINPUT40), .ZN(n597) );
  XNOR2_X1 U684 ( .A(n598), .B(KEYINPUT46), .ZN(n622) );
  INV_X1 U685 ( .A(n599), .ZN(n600) );
  NAND2_X1 U686 ( .A1(n602), .A2(n601), .ZN(n647) );
  NAND2_X1 U687 ( .A1(KEYINPUT47), .A2(n712), .ZN(n603) );
  NAND2_X1 U688 ( .A1(n647), .A2(n603), .ZN(n604) );
  XNOR2_X1 U689 ( .A(n604), .B(KEYINPUT84), .ZN(n607) );
  AND2_X1 U690 ( .A1(n676), .A2(KEYINPUT47), .ZN(n606) );
  XNOR2_X1 U691 ( .A(n608), .B(KEYINPUT85), .ZN(n620) );
  OR2_X1 U692 ( .A1(KEYINPUT47), .A2(n712), .ZN(n609) );
  OR2_X1 U693 ( .A1(n676), .A2(n609), .ZN(n610) );
  XNOR2_X1 U694 ( .A(n610), .B(KEYINPUT75), .ZN(n618) );
  NOR2_X1 U695 ( .A1(n350), .A2(n679), .ZN(n613) );
  AND2_X1 U696 ( .A1(n358), .A2(n612), .ZN(n626) );
  NAND2_X1 U697 ( .A1(n613), .A2(n626), .ZN(n615) );
  INV_X1 U698 ( .A(KEYINPUT36), .ZN(n614) );
  XNOR2_X1 U699 ( .A(n615), .B(n614), .ZN(n617) );
  AND2_X1 U700 ( .A1(n617), .A2(n616), .ZN(n684) );
  NOR2_X1 U701 ( .A1(n618), .A2(n684), .ZN(n619) );
  AND2_X1 U702 ( .A1(n620), .A2(n619), .ZN(n621) );
  INV_X1 U703 ( .A(n692), .ZN(n625) );
  NOR2_X1 U704 ( .A1(n679), .A2(n623), .ZN(n624) );
  AND2_X1 U705 ( .A1(n625), .A2(n624), .ZN(n627) );
  NAND2_X1 U706 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U707 ( .A(n628), .B(KEYINPUT43), .ZN(n629) );
  NOR2_X1 U708 ( .A1(n636), .A2(KEYINPUT86), .ZN(n630) );
  NOR2_X1 U709 ( .A1(n630), .A2(KEYINPUT2), .ZN(n631) );
  INV_X1 U710 ( .A(KEYINPUT2), .ZN(n632) );
  NOR2_X1 U711 ( .A1(n632), .A2(KEYINPUT87), .ZN(n633) );
  NOR2_X1 U712 ( .A1(n636), .A2(n633), .ZN(n634) );
  NAND2_X1 U713 ( .A1(KEYINPUT2), .A2(KEYINPUT87), .ZN(n635) );
  NAND2_X1 U714 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U715 ( .A1(n369), .A2(G210), .ZN(n642) );
  XOR2_X1 U716 ( .A(KEYINPUT89), .B(KEYINPUT55), .Z(n641) );
  XNOR2_X1 U717 ( .A(n639), .B(KEYINPUT54), .ZN(n640) );
  XNOR2_X1 U718 ( .A(n642), .B(n366), .ZN(n643) );
  INV_X1 U719 ( .A(n661), .ZN(n747) );
  NAND2_X1 U720 ( .A1(n643), .A2(n661), .ZN(n645) );
  XNOR2_X1 U721 ( .A(n645), .B(n644), .ZN(G51) );
  XNOR2_X1 U722 ( .A(G143), .B(KEYINPUT112), .ZN(n646) );
  XNOR2_X1 U723 ( .A(n647), .B(n646), .ZN(G45) );
  XNOR2_X1 U724 ( .A(n648), .B(G134), .ZN(G36) );
  XOR2_X1 U725 ( .A(G110), .B(n649), .Z(G12) );
  XOR2_X1 U726 ( .A(G122), .B(KEYINPUT127), .Z(n651) );
  XOR2_X1 U727 ( .A(n651), .B(n368), .Z(G24) );
  XOR2_X1 U728 ( .A(G131), .B(n652), .Z(G33) );
  NAND2_X1 U729 ( .A1(n738), .A2(G472), .ZN(n655) );
  XNOR2_X1 U730 ( .A(n655), .B(n654), .ZN(n656) );
  NAND2_X1 U731 ( .A1(n656), .A2(n661), .ZN(n657) );
  XNOR2_X1 U732 ( .A(n657), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U733 ( .A1(n738), .A2(G475), .ZN(n660) );
  XNOR2_X1 U734 ( .A(n660), .B(n659), .ZN(n662) );
  NAND2_X1 U735 ( .A1(n662), .A2(n661), .ZN(n664) );
  INV_X1 U736 ( .A(KEYINPUT60), .ZN(n663) );
  XNOR2_X1 U737 ( .A(n664), .B(n663), .ZN(G60) );
  XOR2_X1 U738 ( .A(G101), .B(n665), .Z(G3) );
  NOR2_X1 U739 ( .A1(n668), .A2(n679), .ZN(n667) );
  XNOR2_X1 U740 ( .A(G104), .B(KEYINPUT109), .ZN(n666) );
  XNOR2_X1 U741 ( .A(n667), .B(n666), .ZN(G6) );
  NOR2_X1 U742 ( .A1(n668), .A2(n682), .ZN(n670) );
  XNOR2_X1 U743 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n669) );
  XNOR2_X1 U744 ( .A(n670), .B(n669), .ZN(n671) );
  XNOR2_X1 U745 ( .A(G107), .B(n671), .ZN(G9) );
  NOR2_X1 U746 ( .A1(n676), .A2(n682), .ZN(n675) );
  XOR2_X1 U747 ( .A(KEYINPUT110), .B(KEYINPUT29), .Z(n673) );
  XNOR2_X1 U748 ( .A(G128), .B(KEYINPUT111), .ZN(n672) );
  XNOR2_X1 U749 ( .A(n673), .B(n672), .ZN(n674) );
  XNOR2_X1 U750 ( .A(n675), .B(n674), .ZN(G30) );
  INV_X1 U751 ( .A(n676), .ZN(n677) );
  NAND2_X1 U752 ( .A1(n677), .A2(n398), .ZN(n678) );
  XNOR2_X1 U753 ( .A(n678), .B(G146), .ZN(G48) );
  NOR2_X1 U754 ( .A1(n679), .A2(n681), .ZN(n680) );
  XOR2_X1 U755 ( .A(G113), .B(n680), .Z(G15) );
  NOR2_X1 U756 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U757 ( .A(G116), .B(n683), .Z(G18) );
  XNOR2_X1 U758 ( .A(G125), .B(n684), .ZN(n685) );
  XNOR2_X1 U759 ( .A(n685), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U760 ( .A(G140), .B(n686), .ZN(G42) );
  XNOR2_X1 U761 ( .A(n687), .B(KEYINPUT2), .ZN(n727) );
  INV_X1 U762 ( .A(n386), .ZN(n690) );
  NAND2_X1 U763 ( .A1(n690), .A2(n689), .ZN(n702) );
  NOR2_X1 U764 ( .A1(n691), .A2(n692), .ZN(n693) );
  XOR2_X1 U765 ( .A(KEYINPUT50), .B(n693), .Z(n700) );
  XNOR2_X1 U766 ( .A(KEYINPUT49), .B(n695), .ZN(n697) );
  NAND2_X1 U767 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U768 ( .A(n698), .B(KEYINPUT113), .ZN(n699) );
  NAND2_X1 U769 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U770 ( .A1(n702), .A2(n701), .ZN(n704) );
  XOR2_X1 U771 ( .A(KEYINPUT114), .B(KEYINPUT51), .Z(n703) );
  XNOR2_X1 U772 ( .A(n704), .B(n703), .ZN(n705) );
  NAND2_X1 U773 ( .A1(n722), .A2(n705), .ZN(n706) );
  XNOR2_X1 U774 ( .A(n706), .B(KEYINPUT115), .ZN(n717) );
  BUF_X1 U775 ( .A(n707), .Z(n723) );
  INV_X1 U776 ( .A(n723), .ZN(n715) );
  NOR2_X1 U777 ( .A1(n352), .A2(n708), .ZN(n710) );
  NOR2_X1 U778 ( .A1(n711), .A2(n710), .ZN(n713) );
  NOR2_X1 U779 ( .A1(n713), .A2(n364), .ZN(n714) );
  NOR2_X1 U780 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U781 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U782 ( .A(n718), .B(KEYINPUT52), .ZN(n719) );
  XNOR2_X1 U783 ( .A(KEYINPUT116), .B(n719), .ZN(n720) );
  NOR2_X1 U784 ( .A1(n721), .A2(n720), .ZN(n725) );
  AND2_X1 U785 ( .A1(n723), .A2(n722), .ZN(n724) );
  OR2_X1 U786 ( .A1(n725), .A2(n724), .ZN(n726) );
  OR2_X1 U787 ( .A1(n727), .A2(n726), .ZN(n728) );
  NOR2_X1 U788 ( .A1(n728), .A2(G953), .ZN(n729) );
  XNOR2_X1 U789 ( .A(n729), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U790 ( .A1(n742), .A2(G469), .ZN(n736) );
  XOR2_X1 U791 ( .A(KEYINPUT117), .B(KEYINPUT119), .Z(n730) );
  XNOR2_X1 U792 ( .A(n730), .B(KEYINPUT118), .ZN(n732) );
  XOR2_X1 U793 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(n731) );
  XNOR2_X1 U794 ( .A(n732), .B(n731), .ZN(n733) );
  XNOR2_X1 U795 ( .A(n734), .B(n733), .ZN(n735) );
  XNOR2_X1 U796 ( .A(n736), .B(n735), .ZN(n737) );
  NOR2_X1 U797 ( .A1(n747), .A2(n737), .ZN(G54) );
  NAND2_X1 U798 ( .A1(n742), .A2(G478), .ZN(n740) );
  XNOR2_X1 U799 ( .A(n740), .B(n739), .ZN(n741) );
  NOR2_X1 U800 ( .A1(n747), .A2(n741), .ZN(G63) );
  NAND2_X1 U801 ( .A1(n742), .A2(G217), .ZN(n745) );
  XNOR2_X1 U802 ( .A(n743), .B(KEYINPUT120), .ZN(n744) );
  XNOR2_X1 U803 ( .A(n745), .B(n744), .ZN(n746) );
  NOR2_X1 U804 ( .A1(n747), .A2(n746), .ZN(G66) );
  NAND2_X1 U805 ( .A1(n750), .A2(n749), .ZN(n754) );
  NAND2_X1 U806 ( .A1(G953), .A2(G224), .ZN(n751) );
  XNOR2_X1 U807 ( .A(KEYINPUT61), .B(n751), .ZN(n752) );
  NAND2_X1 U808 ( .A1(n752), .A2(G898), .ZN(n753) );
  NAND2_X1 U809 ( .A1(n754), .A2(n753), .ZN(n762) );
  XOR2_X1 U810 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n756) );
  XNOR2_X1 U811 ( .A(n755), .B(n756), .ZN(n757) );
  XOR2_X1 U812 ( .A(G101), .B(n757), .Z(n758) );
  NOR2_X1 U813 ( .A1(n759), .A2(n758), .ZN(n760) );
  XOR2_X1 U814 ( .A(KEYINPUT124), .B(n760), .Z(n761) );
  XNOR2_X1 U815 ( .A(n762), .B(n761), .ZN(n764) );
  XOR2_X1 U816 ( .A(KEYINPUT121), .B(KEYINPUT125), .Z(n763) );
  XNOR2_X1 U817 ( .A(n764), .B(n763), .ZN(G69) );
  XNOR2_X1 U818 ( .A(n766), .B(n765), .ZN(n768) );
  XNOR2_X1 U819 ( .A(n768), .B(n767), .ZN(n773) );
  XOR2_X1 U820 ( .A(KEYINPUT126), .B(n773), .Z(n769) );
  XNOR2_X1 U821 ( .A(G227), .B(n769), .ZN(n770) );
  NAND2_X1 U822 ( .A1(n770), .A2(G900), .ZN(n771) );
  NAND2_X1 U823 ( .A1(n771), .A2(G953), .ZN(n777) );
  XOR2_X1 U824 ( .A(n773), .B(n351), .Z(n775) );
  NAND2_X1 U825 ( .A1(n775), .A2(n774), .ZN(n776) );
  NAND2_X1 U826 ( .A1(n777), .A2(n776), .ZN(G72) );
  XOR2_X1 U827 ( .A(G137), .B(n778), .Z(G39) );
  XOR2_X1 U828 ( .A(G119), .B(n779), .Z(G21) );
endmodule

