//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 1 1 1 0 0 0 0 1 1 1 1 1 1 0 1 0 0 1 1 1 1 0 1 1 1 1 1 0 1 0 0 0 1 0 0 1 0 1 0 1 0 1 0 0 1 1 1 0 1 0 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n770, new_n771, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n866, new_n867, new_n868, new_n870, new_n871,
    new_n872, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n985, new_n986, new_n987, new_n988,
    new_n989;
  INV_X1    g000(.A(KEYINPUT85), .ZN(new_n202));
  XNOR2_X1  g001(.A(G78gat), .B(G106gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT31), .B(G50gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  XOR2_X1   g004(.A(new_n205), .B(KEYINPUT81), .Z(new_n206));
  INV_X1    g005(.A(G228gat), .ZN(new_n207));
  INV_X1    g006(.A(G233gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  AND2_X1   g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT77), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G155gat), .ZN(new_n214));
  INV_X1    g013(.A(G162gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT77), .ZN(new_n217));
  NAND2_X1  g016(.A1(G155gat), .A2(G162gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n213), .A2(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(KEYINPUT78), .B1(new_n218), .B2(KEYINPUT2), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n218), .A2(KEYINPUT78), .A3(KEYINPUT2), .ZN(new_n223));
  AND2_X1   g022(.A1(G141gat), .A2(G148gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(G141gat), .A2(G148gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n222), .A2(new_n223), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n216), .A2(new_n218), .ZN(new_n228));
  AND2_X1   g027(.A1(new_n228), .A2(new_n226), .ZN(new_n229));
  AND2_X1   g028(.A1(KEYINPUT79), .A2(G155gat), .ZN(new_n230));
  NOR2_X1   g029(.A1(KEYINPUT79), .A2(G155gat), .ZN(new_n231));
  OAI21_X1  g030(.A(G162gat), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT2), .ZN(new_n233));
  AOI22_X1  g032(.A1(new_n220), .A2(new_n227), .B1(new_n229), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT29), .ZN(new_n235));
  XNOR2_X1  g034(.A(G211gat), .B(G218gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(G197gat), .B(G204gat), .ZN(new_n237));
  INV_X1    g036(.A(G211gat), .ZN(new_n238));
  INV_X1    g037(.A(G218gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT73), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT73), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(G218gat), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n238), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n236), .B(new_n237), .C1(new_n243), .C2(KEYINPUT22), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT22), .ZN(new_n246));
  XNOR2_X1  g045(.A(KEYINPUT73), .B(G218gat), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n246), .B1(new_n247), .B2(new_n238), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n236), .B1(new_n248), .B2(new_n237), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n235), .B1(new_n245), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n234), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n236), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n240), .A2(new_n242), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT22), .B1(new_n254), .B2(G211gat), .ZN(new_n255));
  INV_X1    g054(.A(new_n237), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n253), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT74), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n257), .A2(new_n258), .A3(new_n244), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n249), .A2(KEYINPUT74), .ZN(new_n260));
  OR2_X1    g059(.A1(KEYINPUT79), .A2(G155gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(KEYINPUT79), .A2(G155gat), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n215), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT2), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n226), .B(new_n228), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n223), .ZN(new_n266));
  XNOR2_X1  g065(.A(G141gat), .B(G148gat), .ZN(new_n267));
  NOR3_X1   g066(.A1(new_n266), .A2(new_n267), .A3(new_n221), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n213), .A2(new_n219), .ZN(new_n269));
  OAI211_X1 g068(.A(new_n265), .B(new_n251), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  AOI22_X1  g069(.A1(new_n259), .A2(new_n260), .B1(new_n270), .B2(new_n235), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n210), .B1(new_n252), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n261), .A2(new_n262), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n264), .B1(new_n273), .B2(G162gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n228), .A2(new_n226), .ZN(new_n275));
  OAI22_X1  g074(.A1(new_n268), .A2(new_n269), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT80), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n265), .B(KEYINPUT80), .C1(new_n268), .C2(new_n269), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n259), .A2(new_n235), .A3(new_n260), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n280), .B1(new_n251), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n259), .A2(new_n260), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n270), .A2(new_n235), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(new_n209), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n272), .B1(new_n282), .B2(new_n286), .ZN(new_n287));
  XOR2_X1   g086(.A(KEYINPUT82), .B(G22gat), .Z(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  AND3_X1   g088(.A1(new_n287), .A2(KEYINPUT84), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(KEYINPUT84), .B1(new_n287), .B2(new_n289), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n272), .B(new_n288), .C1(new_n282), .C2(new_n286), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT83), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n281), .A2(new_n251), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n295), .A2(new_n278), .A3(new_n279), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n271), .A2(new_n210), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT83), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n298), .A2(new_n299), .A3(new_n272), .A4(new_n288), .ZN(new_n300));
  AND2_X1   g099(.A1(new_n294), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n206), .B1(new_n292), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n205), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n293), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n304), .B1(G22gat), .B2(new_n287), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n202), .B1(new_n302), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT84), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT29), .B1(new_n257), .B2(new_n244), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n276), .B1(new_n308), .B2(KEYINPUT3), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n285), .A2(new_n309), .ZN(new_n310));
  AOI22_X1  g109(.A1(new_n296), .A2(new_n297), .B1(new_n310), .B2(new_n210), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n307), .B1(new_n311), .B2(new_n288), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n287), .A2(KEYINPUT84), .A3(new_n289), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n312), .A2(new_n313), .A3(new_n294), .A4(new_n300), .ZN(new_n314));
  INV_X1    g113(.A(new_n206), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n305), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(KEYINPUT85), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT5), .ZN(new_n318));
  INV_X1    g117(.A(G127gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G134gat), .ZN(new_n320));
  INV_X1    g119(.A(G134gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(G127gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT1), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n325), .B1(G113gat), .B2(G120gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(G113gat), .A2(G120gat), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n324), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT71), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n323), .A2(new_n331), .ZN(new_n332));
  OAI22_X1  g131(.A1(new_n326), .A2(new_n328), .B1(new_n320), .B2(KEYINPUT71), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n330), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n278), .A2(new_n279), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n324), .A2(KEYINPUT71), .ZN(new_n336));
  INV_X1    g135(.A(new_n333), .ZN(new_n337));
  AOI22_X1  g136(.A1(new_n336), .A2(new_n337), .B1(new_n329), .B2(new_n324), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n234), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n335), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(G225gat), .A2(G233gat), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n318), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n278), .A2(KEYINPUT3), .A3(new_n279), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n338), .B1(new_n234), .B2(new_n251), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT4), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n347), .B1(new_n276), .B2(new_n334), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n234), .A2(KEYINPUT4), .A3(new_n338), .ZN(new_n349));
  AND2_X1   g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n346), .A2(new_n350), .A3(new_n341), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n343), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n348), .A2(new_n349), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n353), .B1(new_n344), .B2(new_n345), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n354), .A2(new_n318), .A3(new_n341), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(G1gat), .B(G29gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n357), .B(KEYINPUT0), .ZN(new_n358));
  XNOR2_X1  g157(.A(G57gat), .B(G85gat), .ZN(new_n359));
  XOR2_X1   g158(.A(new_n358), .B(new_n359), .Z(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n356), .A2(KEYINPUT6), .A3(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n352), .A2(new_n360), .A3(new_n355), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT6), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n360), .B1(new_n352), .B2(new_n355), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n362), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(G8gat), .B(G36gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(G64gat), .B(G92gat), .ZN(new_n369));
  XOR2_X1   g168(.A(new_n368), .B(new_n369), .Z(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(G169gat), .A2(G176gat), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT23), .ZN(new_n374));
  NOR3_X1   g173(.A1(new_n374), .A2(G169gat), .A3(G176gat), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n373), .B1(new_n375), .B2(KEYINPUT66), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT65), .ZN(new_n377));
  INV_X1    g176(.A(G183gat), .ZN(new_n378));
  INV_X1    g177(.A(G190gat), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(G183gat), .A2(G190gat), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT24), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n384));
  OAI21_X1  g183(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n380), .A2(new_n383), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(G169gat), .ZN(new_n387));
  INV_X1    g186(.A(G176gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT67), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n390), .A2(KEYINPUT23), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n374), .A2(KEYINPUT67), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n389), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NOR2_X1   g192(.A1(G169gat), .A2(G176gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT23), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT66), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n376), .A2(new_n386), .A3(new_n393), .A4(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT25), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n383), .B(new_n384), .C1(G183gat), .C2(G190gat), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n395), .A2(KEYINPUT25), .A3(new_n372), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n374), .A2(KEYINPUT67), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n390), .A2(KEYINPUT23), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n394), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  AOI22_X1  g204(.A1(new_n398), .A2(new_n399), .B1(new_n400), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n407));
  AOI22_X1  g206(.A1(new_n407), .A2(KEYINPUT69), .B1(G169gat), .B2(G176gat), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT69), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n389), .A2(new_n409), .A3(KEYINPUT26), .ZN(new_n410));
  NOR4_X1   g209(.A1(KEYINPUT70), .A2(KEYINPUT26), .A3(G169gat), .A4(G176gat), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT70), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT26), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n412), .B1(new_n394), .B2(new_n413), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n408), .B(new_n410), .C1(new_n411), .C2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n378), .A2(KEYINPUT27), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT27), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(G183gat), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n416), .A2(new_n418), .A3(new_n379), .ZN(new_n419));
  XNOR2_X1  g218(.A(KEYINPUT68), .B(KEYINPUT28), .ZN(new_n420));
  OR2_X1    g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI22_X1  g220(.A1(new_n419), .A2(new_n420), .B1(G183gat), .B2(G190gat), .ZN(new_n422));
  AND3_X1   g221(.A1(new_n415), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n235), .B1(new_n406), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(G226gat), .A2(G233gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n283), .ZN(new_n427));
  INV_X1    g226(.A(new_n425), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n428), .B1(new_n406), .B2(new_n423), .ZN(new_n429));
  AND3_X1   g228(.A1(new_n426), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n427), .B1(new_n426), .B2(new_n429), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n371), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n415), .A2(new_n421), .A3(new_n422), .ZN(new_n433));
  AND2_X1   g232(.A1(new_n398), .A2(new_n399), .ZN(new_n434));
  AND2_X1   g233(.A1(new_n405), .A2(new_n400), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n428), .B1(new_n436), .B2(new_n235), .ZN(new_n437));
  INV_X1    g236(.A(new_n429), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n283), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n426), .A2(new_n427), .A3(new_n429), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n439), .A2(new_n440), .A3(new_n370), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT30), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n432), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT75), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT76), .ZN(new_n446));
  NOR3_X1   g245(.A1(new_n430), .A2(new_n431), .A3(new_n371), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n446), .B1(new_n447), .B2(KEYINPUT30), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n441), .A2(KEYINPUT76), .A3(new_n442), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n432), .B(KEYINPUT75), .C1(new_n441), .C2(new_n442), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n367), .A2(new_n445), .A3(new_n450), .A4(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n306), .A2(new_n317), .A3(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT72), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n454), .B(new_n433), .C1(new_n434), .C2(new_n435), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT72), .B1(new_n406), .B2(new_n423), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n455), .A2(new_n456), .A3(new_n334), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n436), .A2(KEYINPUT72), .A3(new_n338), .ZN(new_n458));
  NAND2_X1  g257(.A1(G227gat), .A2(G233gat), .ZN(new_n459));
  XOR2_X1   g258(.A(new_n459), .B(KEYINPUT64), .Z(new_n460));
  NAND3_X1  g259(.A1(new_n457), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT32), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT33), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  XOR2_X1   g263(.A(G15gat), .B(G43gat), .Z(new_n465));
  XNOR2_X1  g264(.A(G71gat), .B(G99gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n465), .B(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n462), .A2(new_n464), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n457), .A2(new_n458), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n459), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n460), .A2(KEYINPUT34), .ZN(new_n471));
  AOI22_X1  g270(.A1(new_n470), .A2(KEYINPUT34), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n467), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n461), .B(KEYINPUT32), .C1(new_n463), .C2(new_n473), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n468), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n472), .B1(new_n468), .B2(new_n474), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT36), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n468), .A2(new_n474), .ZN(new_n479));
  INV_X1    g278(.A(new_n472), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n468), .A2(new_n472), .A3(new_n474), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT36), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n478), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n366), .A2(KEYINPUT88), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT88), .ZN(new_n488));
  AOI211_X1 g287(.A(new_n488), .B(new_n360), .C1(new_n352), .C2(new_n355), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n341), .B1(new_n346), .B2(new_n350), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT39), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n361), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n335), .A2(new_n341), .A3(new_n339), .ZN(new_n494));
  OAI211_X1 g293(.A(KEYINPUT39), .B(new_n494), .C1(new_n354), .C2(new_n341), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n493), .A2(KEYINPUT40), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT89), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT89), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n493), .A2(new_n495), .A3(new_n498), .A4(KEYINPUT40), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n493), .A2(new_n495), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT87), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT40), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n493), .A2(KEYINPUT87), .A3(new_n495), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n500), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n370), .B1(new_n439), .B2(new_n440), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n508), .B1(KEYINPUT30), .B2(new_n447), .ZN(new_n509));
  AND3_X1   g308(.A1(new_n441), .A2(KEYINPUT76), .A3(new_n442), .ZN(new_n510));
  AOI21_X1  g309(.A(KEYINPUT76), .B1(new_n441), .B2(new_n442), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT86), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n450), .A2(KEYINPUT86), .A3(new_n509), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n507), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AND4_X1   g315(.A1(new_n318), .A2(new_n346), .A3(new_n341), .A4(new_n350), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n517), .B1(new_n351), .B2(new_n343), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n488), .B1(new_n518), .B2(new_n360), .ZN(new_n519));
  AND2_X1   g318(.A1(new_n363), .A2(new_n364), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n366), .A2(KEYINPUT88), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n439), .B1(new_n430), .B2(KEYINPUT90), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT90), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n440), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g324(.A(KEYINPUT37), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(KEYINPUT91), .B(KEYINPUT38), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n371), .A2(KEYINPUT37), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n526), .B(new_n527), .C1(new_n508), .C2(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT37), .B1(new_n430), .B2(new_n431), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n531), .B1(new_n508), .B2(new_n529), .ZN(new_n532));
  INV_X1    g331(.A(new_n527), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n447), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n522), .A2(new_n362), .A3(new_n530), .A4(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n314), .A2(new_n315), .ZN(new_n536));
  INV_X1    g335(.A(new_n305), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  OAI211_X1 g338(.A(new_n453), .B(new_n486), .C1(new_n516), .C2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT92), .ZN(new_n541));
  NOR3_X1   g340(.A1(new_n452), .A2(new_n316), .A3(new_n483), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT35), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n538), .A2(new_n514), .A3(new_n515), .A4(new_n477), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n522), .A2(new_n362), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(new_n543), .ZN(new_n546));
  OAI22_X1  g345(.A1(new_n542), .A2(new_n543), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  AND3_X1   g346(.A1(new_n540), .A2(new_n541), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n541), .B1(new_n540), .B2(new_n547), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(G29gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT14), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT14), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(G29gat), .ZN(new_n554));
  INV_X1    g353(.A(G36gat), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n552), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n556), .B1(new_n555), .B2(new_n552), .ZN(new_n557));
  XNOR2_X1  g356(.A(G43gat), .B(G50gat), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n557), .B1(KEYINPUT15), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT93), .ZN(new_n560));
  OR2_X1    g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n558), .A2(new_n560), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n561), .A2(KEYINPUT15), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n561), .A2(new_n557), .A3(KEYINPUT15), .A4(new_n562), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT94), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT17), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT94), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n564), .A2(new_n569), .A3(new_n565), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n567), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G15gat), .B(G22gat), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT16), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n572), .B1(new_n573), .B2(G1gat), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n574), .B1(G1gat), .B2(new_n572), .ZN(new_n575));
  INV_X1    g374(.A(G8gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n566), .A2(KEYINPUT17), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n571), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(G229gat), .A2(G233gat), .ZN(new_n580));
  INV_X1    g379(.A(new_n577), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n567), .A2(new_n581), .A3(new_n570), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n579), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT18), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n579), .A2(KEYINPUT18), .A3(new_n580), .A4(new_n582), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n567), .A2(new_n570), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(new_n577), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(new_n582), .ZN(new_n589));
  XOR2_X1   g388(.A(new_n580), .B(KEYINPUT13), .Z(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n585), .A2(new_n586), .A3(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G113gat), .B(G141gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(G197gat), .ZN(new_n594));
  XOR2_X1   g393(.A(KEYINPUT11), .B(G169gat), .Z(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(KEYINPUT12), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n592), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n585), .A2(new_n591), .A3(new_n586), .A4(new_n597), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  OR2_X1    g401(.A1(G57gat), .A2(G64gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(G57gat), .A2(G64gat), .ZN(new_n604));
  AND2_X1   g403(.A1(G71gat), .A2(G78gat), .ZN(new_n605));
  OAI211_X1 g404(.A(new_n603), .B(new_n604), .C1(new_n605), .C2(KEYINPUT9), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n606), .B1(KEYINPUT95), .B2(new_n605), .ZN(new_n607));
  NOR2_X1   g406(.A1(G71gat), .A2(G78gat), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  AND2_X1   g408(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n607), .A2(new_n609), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT21), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G231gat), .A2(G233gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  OR2_X1    g415(.A1(new_n616), .A2(new_n319), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n319), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n577), .B1(new_n612), .B2(new_n613), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n617), .A2(new_n620), .A3(new_n618), .ZN(new_n623));
  XNOR2_X1  g422(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT96), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(G155gat), .ZN(new_n626));
  XOR2_X1   g425(.A(G183gat), .B(G211gat), .Z(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  AND3_X1   g427(.A1(new_n622), .A2(new_n623), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n628), .B1(new_n622), .B2(new_n623), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g430(.A(G190gat), .B(G218gat), .Z(new_n632));
  XNOR2_X1  g431(.A(KEYINPUT97), .B(KEYINPUT7), .ZN(new_n633));
  NAND2_X1  g432(.A1(G85gat), .A2(G92gat), .ZN(new_n634));
  OR2_X1    g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND2_X1  g435(.A1(G99gat), .A2(G106gat), .ZN(new_n637));
  INV_X1    g436(.A(G85gat), .ZN(new_n638));
  INV_X1    g437(.A(G92gat), .ZN(new_n639));
  AOI22_X1  g438(.A1(KEYINPUT8), .A2(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n635), .A2(new_n636), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g440(.A(G99gat), .B(G106gat), .Z(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  AND3_X1   g442(.A1(new_n571), .A2(new_n578), .A3(new_n643), .ZN(new_n644));
  OR2_X1    g443(.A1(new_n641), .A2(new_n642), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n641), .A2(new_n642), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n567), .A2(new_n570), .A3(new_n645), .A4(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(G232gat), .A2(G233gat), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(KEYINPUT41), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n632), .B1(new_n644), .B2(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n649), .A2(KEYINPUT41), .ZN(new_n653));
  XNOR2_X1  g452(.A(G134gat), .B(G162gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n571), .A2(new_n578), .A3(new_n643), .ZN(new_n656));
  INV_X1    g455(.A(new_n632), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n656), .A2(new_n657), .A3(new_n647), .A4(new_n650), .ZN(new_n658));
  AND3_X1   g457(.A1(new_n652), .A2(new_n655), .A3(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n655), .B1(new_n652), .B2(new_n658), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(G230gat), .A2(G233gat), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n643), .A2(new_n612), .ZN(new_n665));
  OAI211_X1 g464(.A(new_n645), .B(new_n646), .C1(new_n610), .C2(new_n611), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT10), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  OR3_X1    g467(.A1(new_n643), .A2(new_n667), .A3(new_n612), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n664), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n663), .B1(new_n665), .B2(new_n666), .ZN(new_n671));
  XNOR2_X1  g470(.A(G120gat), .B(G148gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(G176gat), .B(G204gat), .ZN(new_n673));
  XOR2_X1   g472(.A(new_n672), .B(new_n673), .Z(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  OR3_X1    g474(.A1(new_n670), .A2(new_n671), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n675), .B1(new_n670), .B2(new_n671), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n631), .A2(new_n662), .A3(new_n679), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n550), .A2(new_n602), .A3(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n367), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(KEYINPUT98), .B(G1gat), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(G1324gat));
  NAND2_X1  g484(.A1(new_n514), .A2(new_n515), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT99), .B(KEYINPUT16), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(G8gat), .ZN(new_n688));
  AND3_X1   g487(.A1(new_n681), .A2(new_n686), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n576), .B1(new_n681), .B2(new_n686), .ZN(new_n690));
  OAI21_X1  g489(.A(KEYINPUT42), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n691), .B1(KEYINPUT42), .B2(new_n689), .ZN(G1325gat));
  INV_X1    g491(.A(G15gat), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n681), .A2(new_n693), .A3(new_n477), .ZN(new_n694));
  INV_X1    g493(.A(new_n486), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n681), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n694), .B1(new_n697), .B2(new_n693), .ZN(G1326gat));
  NAND2_X1  g497(.A1(new_n306), .A2(new_n317), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n681), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(KEYINPUT43), .B(G22gat), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(G1327gat));
  NOR3_X1   g502(.A1(new_n631), .A2(new_n602), .A3(new_n678), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n705), .A2(new_n662), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n706), .B1(new_n548), .B2(new_n549), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n708), .A2(new_n551), .A3(new_n682), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT45), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n662), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n712), .B1(new_n548), .B2(new_n549), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n540), .A2(new_n547), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n661), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(new_n711), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n713), .A2(new_n716), .A3(new_n704), .ZN(new_n717));
  OAI21_X1  g516(.A(G29gat), .B1(new_n717), .B2(new_n367), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n710), .A2(new_n718), .ZN(G1328gat));
  NAND3_X1  g518(.A1(new_n708), .A2(new_n555), .A3(new_n686), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n720), .B(KEYINPUT46), .Z(new_n721));
  INV_X1    g520(.A(new_n686), .ZN(new_n722));
  OAI21_X1  g521(.A(G36gat), .B1(new_n717), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n723), .ZN(G1329gat));
  OAI21_X1  g523(.A(G43gat), .B1(new_n717), .B2(new_n486), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n483), .A2(G43gat), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n708), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g526(.A(KEYINPUT100), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT47), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(G1330gat));
  INV_X1    g529(.A(KEYINPUT103), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n713), .A2(new_n316), .A3(new_n716), .A4(new_n704), .ZN(new_n732));
  AND2_X1   g531(.A1(KEYINPUT48), .A2(G50gat), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT101), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n707), .A2(new_n735), .ZN(new_n736));
  OAI211_X1 g535(.A(KEYINPUT101), .B(new_n706), .C1(new_n548), .C2(new_n549), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n699), .A2(G50gat), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n736), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT48), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(KEYINPUT102), .ZN(new_n741));
  AND3_X1   g540(.A1(new_n734), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n713), .A2(new_n700), .A3(new_n716), .A4(new_n704), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(G50gat), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n736), .A2(KEYINPUT102), .A3(new_n737), .A4(new_n738), .ZN(new_n745));
  AOI21_X1  g544(.A(KEYINPUT48), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n731), .B1(new_n742), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n744), .A2(new_n745), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n740), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n734), .A2(new_n739), .A3(new_n741), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n749), .A2(KEYINPUT103), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n747), .A2(new_n751), .ZN(G1331gat));
  INV_X1    g551(.A(new_n631), .ZN(new_n753));
  NOR4_X1   g552(.A1(new_n753), .A2(new_n601), .A3(new_n661), .A4(new_n679), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n714), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT104), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n682), .ZN(new_n757));
  XNOR2_X1  g556(.A(KEYINPUT105), .B(G57gat), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n757), .B(new_n758), .ZN(G1332gat));
  NAND2_X1  g558(.A1(new_n756), .A2(new_n686), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n760), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n761));
  XOR2_X1   g560(.A(KEYINPUT49), .B(G64gat), .Z(new_n762));
  OAI21_X1  g561(.A(new_n761), .B1(new_n760), .B2(new_n762), .ZN(G1333gat));
  INV_X1    g562(.A(G71gat), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n756), .A2(new_n764), .A3(new_n477), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n756), .A2(new_n695), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n765), .B1(new_n766), .B2(new_n764), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT50), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n767), .B(new_n768), .ZN(G1334gat));
  NAND2_X1  g568(.A1(new_n756), .A2(new_n700), .ZN(new_n770));
  XOR2_X1   g569(.A(KEYINPUT106), .B(G78gat), .Z(new_n771));
  XNOR2_X1  g570(.A(new_n770), .B(new_n771), .ZN(G1335gat));
  NOR2_X1   g571(.A1(new_n631), .A2(new_n601), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(new_n678), .ZN(new_n774));
  XOR2_X1   g573(.A(new_n774), .B(KEYINPUT107), .Z(new_n775));
  NAND3_X1  g574(.A1(new_n713), .A2(new_n716), .A3(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(G85gat), .B1(new_n776), .B2(new_n367), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n714), .A2(new_n661), .A3(new_n773), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT51), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n778), .B(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n682), .A2(new_n638), .A3(new_n678), .ZN(new_n782));
  XOR2_X1   g581(.A(new_n782), .B(KEYINPUT108), .Z(new_n783));
  OAI21_X1  g582(.A(new_n777), .B1(new_n781), .B2(new_n783), .ZN(G1336gat));
  NOR3_X1   g583(.A1(new_n722), .A2(G92gat), .A3(new_n679), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(new_n778), .ZN(new_n787));
  XNOR2_X1  g586(.A(KEYINPUT109), .B(KEYINPUT51), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT110), .ZN(new_n790));
  AOI22_X1  g589(.A1(new_n789), .A2(new_n790), .B1(KEYINPUT51), .B2(new_n787), .ZN(new_n791));
  OAI21_X1  g590(.A(KEYINPUT110), .B1(new_n787), .B2(new_n788), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n786), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n713), .A2(new_n686), .A3(new_n716), .A4(new_n775), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(G92gat), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(KEYINPUT52), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT111), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT52), .B1(new_n780), .B2(new_n785), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n798), .B1(new_n799), .B2(new_n795), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n799), .A2(new_n798), .A3(new_n795), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n797), .B1(new_n800), .B2(new_n801), .ZN(G1337gat));
  OAI21_X1  g601(.A(G99gat), .B1(new_n776), .B2(new_n486), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n483), .A2(G99gat), .A3(new_n679), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n804), .B(KEYINPUT112), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n803), .B1(new_n781), .B2(new_n805), .ZN(G1338gat));
  NOR3_X1   g605(.A1(new_n538), .A2(G106gat), .A3(new_n679), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n808), .B1(new_n791), .B2(new_n792), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n776), .A2(new_n699), .ZN(new_n810));
  INV_X1    g609(.A(G106gat), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(KEYINPUT53), .B1(new_n809), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(KEYINPUT53), .B1(new_n780), .B2(new_n807), .ZN(new_n814));
  OAI21_X1  g613(.A(G106gat), .B1(new_n776), .B2(new_n538), .ZN(new_n815));
  AOI21_X1  g614(.A(KEYINPUT113), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AND3_X1   g615(.A1(new_n814), .A2(KEYINPUT113), .A3(new_n815), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n813), .B1(new_n816), .B2(new_n817), .ZN(G1339gat));
  NAND2_X1  g617(.A1(new_n668), .A2(new_n669), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n663), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n668), .A2(new_n669), .A3(new_n664), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n820), .A2(KEYINPUT54), .A3(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n674), .B1(new_n670), .B2(new_n823), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n822), .A2(KEYINPUT55), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(KEYINPUT55), .B1(new_n822), .B2(new_n824), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n670), .A2(new_n671), .A3(new_n675), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n825), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT115), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n589), .A2(new_n590), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n580), .B1(new_n579), .B2(new_n582), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n596), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n678), .A2(new_n600), .A3(new_n832), .ZN(new_n833));
  AOI22_X1  g632(.A1(new_n828), .A2(new_n601), .B1(new_n829), .B2(new_n833), .ZN(new_n834));
  AND3_X1   g633(.A1(new_n678), .A2(new_n600), .A3(new_n832), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(KEYINPUT115), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n661), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n600), .A2(new_n832), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n824), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT55), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n827), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n822), .A2(KEYINPUT55), .A3(new_n824), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n838), .A2(new_n661), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT114), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n828), .A2(KEYINPUT114), .A3(new_n661), .A4(new_n838), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n753), .B1(new_n837), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n680), .A2(new_n601), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  AOI211_X1 g649(.A(new_n367), .B(new_n544), .C1(new_n848), .C2(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(G113gat), .B1(new_n851), .B2(new_n601), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n848), .A2(new_n850), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n700), .A2(new_n483), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n686), .A2(new_n367), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n601), .A2(G113gat), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n852), .B1(new_n858), .B2(new_n859), .ZN(G1340gat));
  INV_X1    g659(.A(G120gat), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n861), .B1(new_n858), .B2(new_n678), .ZN(new_n862));
  XOR2_X1   g661(.A(new_n862), .B(KEYINPUT116), .Z(new_n863));
  NAND3_X1  g662(.A1(new_n851), .A2(new_n861), .A3(new_n678), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(G1341gat));
  INV_X1    g664(.A(new_n858), .ZN(new_n866));
  OAI21_X1  g665(.A(G127gat), .B1(new_n866), .B2(new_n753), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n851), .A2(new_n319), .A3(new_n631), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(G1342gat));
  NAND3_X1  g668(.A1(new_n851), .A2(new_n321), .A3(new_n661), .ZN(new_n870));
  XOR2_X1   g669(.A(new_n870), .B(KEYINPUT56), .Z(new_n871));
  OAI21_X1  g670(.A(G134gat), .B1(new_n866), .B2(new_n662), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(G1343gat));
  NOR2_X1   g672(.A1(new_n857), .A2(new_n695), .ZN(new_n874));
  INV_X1    g673(.A(G141gat), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n602), .A2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT117), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n699), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n835), .B1(new_n828), .B2(new_n601), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n845), .B(new_n846), .C1(new_n880), .C2(new_n661), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n881), .A2(new_n753), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n877), .B(new_n879), .C1(new_n882), .C2(new_n849), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n849), .B1(new_n881), .B2(new_n753), .ZN(new_n884));
  INV_X1    g683(.A(new_n879), .ZN(new_n885));
  OAI21_X1  g684(.A(KEYINPUT117), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n538), .B1(new_n848), .B2(new_n850), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n888), .A2(KEYINPUT57), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n874), .B(new_n876), .C1(new_n887), .C2(new_n889), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n695), .A2(new_n538), .A3(new_n686), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n853), .A2(new_n682), .A3(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n875), .B1(new_n892), .B2(new_n602), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  XOR2_X1   g693(.A(KEYINPUT118), .B(KEYINPUT58), .Z(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(KEYINPUT119), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT119), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n894), .A2(new_n898), .A3(new_n895), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n890), .A2(KEYINPUT58), .A3(new_n893), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n897), .A2(new_n899), .A3(new_n900), .ZN(G1344gat));
  INV_X1    g700(.A(KEYINPUT59), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n874), .B1(new_n887), .B2(new_n889), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n902), .B(G148gat), .C1(new_n903), .C2(new_n679), .ZN(new_n904));
  INV_X1    g703(.A(G148gat), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n828), .A2(new_n601), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n661), .B1(new_n906), .B2(new_n833), .ZN(new_n907));
  INV_X1    g706(.A(new_n843), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n753), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n850), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(KEYINPUT120), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n700), .B1(new_n910), .B2(KEYINPUT120), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n878), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n888), .A2(KEYINPUT57), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n857), .A2(new_n695), .A3(new_n679), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n905), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n904), .B1(new_n918), .B2(new_n902), .ZN(new_n919));
  AND3_X1   g718(.A1(new_n853), .A2(new_n682), .A3(new_n891), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n920), .A2(new_n905), .A3(new_n678), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n919), .A2(new_n921), .ZN(G1345gat));
  OAI21_X1  g721(.A(new_n273), .B1(new_n903), .B2(new_n753), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n631), .A2(new_n261), .A3(new_n262), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n923), .B1(new_n892), .B2(new_n924), .ZN(G1346gat));
  OAI21_X1  g724(.A(G162gat), .B1(new_n903), .B2(new_n662), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n920), .A2(new_n215), .A3(new_n661), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(G1347gat));
  NOR2_X1   g727(.A1(new_n722), .A2(new_n682), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n853), .A2(new_n854), .A3(new_n929), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n930), .A2(new_n387), .A3(new_n602), .ZN(new_n931));
  INV_X1    g730(.A(new_n929), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n932), .B1(new_n848), .B2(new_n850), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n316), .A2(new_n483), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n933), .A2(new_n934), .A3(new_n601), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n931), .B1(new_n935), .B2(new_n387), .ZN(G1348gat));
  OAI21_X1  g735(.A(G176gat), .B1(new_n930), .B2(new_n679), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n933), .A2(new_n934), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n678), .A2(new_n388), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(G1349gat));
  OAI21_X1  g739(.A(G183gat), .B1(new_n930), .B2(new_n753), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n631), .A2(new_n416), .A3(new_n418), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n941), .B1(new_n938), .B2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT60), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n944), .A2(KEYINPUT121), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n943), .B(new_n945), .ZN(G1350gat));
  NOR3_X1   g745(.A1(new_n938), .A2(G190gat), .A3(new_n662), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT122), .ZN(new_n948));
  OAI21_X1  g747(.A(G190gat), .B1(new_n930), .B2(new_n662), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(KEYINPUT61), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n948), .A2(new_n950), .ZN(G1351gat));
  NAND4_X1  g750(.A1(new_n853), .A2(new_n316), .A3(new_n486), .A4(new_n929), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT123), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  XOR2_X1   g753(.A(KEYINPUT124), .B(G197gat), .Z(new_n955));
  NAND3_X1  g754(.A1(new_n954), .A2(new_n601), .A3(new_n955), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n932), .A2(new_n695), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n916), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n958), .A2(new_n602), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n956), .B1(new_n959), .B2(new_n955), .ZN(G1352gat));
  AND2_X1   g759(.A1(new_n909), .A2(new_n850), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT120), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n699), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g762(.A(KEYINPUT57), .B1(new_n963), .B2(new_n911), .ZN(new_n964));
  INV_X1    g763(.A(new_n915), .ZN(new_n965));
  OAI211_X1 g764(.A(new_n678), .B(new_n957), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(KEYINPUT126), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT126), .ZN(new_n968));
  NAND4_X1  g767(.A1(new_n916), .A2(new_n968), .A3(new_n678), .A4(new_n957), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n967), .A2(G204gat), .A3(new_n969), .ZN(new_n970));
  OR3_X1    g769(.A1(new_n952), .A2(G204gat), .A3(new_n679), .ZN(new_n971));
  AND3_X1   g770(.A1(new_n971), .A2(KEYINPUT125), .A3(KEYINPUT62), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT125), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT62), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n973), .A2(new_n974), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n975), .B1(new_n971), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n972), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n970), .A2(new_n978), .ZN(G1353gat));
  NAND3_X1  g778(.A1(new_n954), .A2(new_n238), .A3(new_n631), .ZN(new_n980));
  OAI211_X1 g779(.A(new_n631), .B(new_n957), .C1(new_n964), .C2(new_n965), .ZN(new_n981));
  AND3_X1   g780(.A1(new_n981), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n982));
  AOI21_X1  g781(.A(KEYINPUT63), .B1(new_n981), .B2(G211gat), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n980), .B1(new_n982), .B2(new_n983), .ZN(G1354gat));
  NOR3_X1   g783(.A1(new_n958), .A2(new_n247), .A3(new_n662), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n239), .B1(new_n953), .B2(new_n662), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n986), .A2(KEYINPUT127), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT127), .ZN(new_n988));
  OAI211_X1 g787(.A(new_n988), .B(new_n239), .C1(new_n953), .C2(new_n662), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n985), .B1(new_n987), .B2(new_n989), .ZN(G1355gat));
endmodule


