

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U560 ( .A(n707), .ZN(n743) );
  NOR2_X1 U561 ( .A1(n732), .A2(n731), .ZN(n733) );
  INV_X1 U562 ( .A(KEYINPUT101), .ZN(n766) );
  NAND2_X1 U563 ( .A1(n826), .A2(n815), .ZN(n816) );
  NOR2_X1 U564 ( .A1(G164), .A2(G1384), .ZN(n785) );
  OR2_X1 U565 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U566 ( .A(n591), .B(KEYINPUT15), .ZN(n999) );
  NOR2_X1 U567 ( .A1(n655), .A2(G651), .ZN(n653) );
  XNOR2_X1 U568 ( .A(KEYINPUT85), .B(n541), .ZN(G164) );
  XNOR2_X1 U569 ( .A(KEYINPUT17), .B(KEYINPUT65), .ZN(n530) );
  NOR2_X1 U570 ( .A1(G2105), .A2(G2104), .ZN(n529) );
  XNOR2_X2 U571 ( .A(n530), .B(n529), .ZN(n897) );
  NAND2_X1 U572 ( .A1(n897), .A2(G138), .ZN(n540) );
  AND2_X1 U573 ( .A1(G2105), .A2(G2104), .ZN(n900) );
  NAND2_X1 U574 ( .A1(G114), .A2(n900), .ZN(n534) );
  INV_X1 U575 ( .A(G2105), .ZN(n531) );
  NOR2_X1 U576 ( .A1(n531), .A2(G2104), .ZN(n532) );
  XNOR2_X2 U577 ( .A(n532), .B(KEYINPUT64), .ZN(n901) );
  NAND2_X1 U578 ( .A1(G126), .A2(n901), .ZN(n533) );
  NAND2_X1 U579 ( .A1(n534), .A2(n533), .ZN(n538) );
  AND2_X1 U580 ( .A1(G2104), .A2(G102), .ZN(n535) );
  NAND2_X1 U581 ( .A1(n531), .A2(n535), .ZN(n536) );
  XOR2_X1 U582 ( .A(n536), .B(KEYINPUT84), .Z(n537) );
  NOR2_X1 U583 ( .A1(n538), .A2(n537), .ZN(n539) );
  NAND2_X1 U584 ( .A1(n540), .A2(n539), .ZN(n541) );
  NAND2_X1 U585 ( .A1(G137), .A2(n897), .ZN(n542) );
  XNOR2_X1 U586 ( .A(n542), .B(KEYINPUT66), .ZN(n549) );
  AND2_X1 U587 ( .A1(n531), .A2(G2104), .ZN(n896) );
  NAND2_X1 U588 ( .A1(G101), .A2(n896), .ZN(n543) );
  XNOR2_X1 U589 ( .A(KEYINPUT23), .B(n543), .ZN(n547) );
  NAND2_X1 U590 ( .A1(G113), .A2(n900), .ZN(n545) );
  NAND2_X1 U591 ( .A1(G125), .A2(n901), .ZN(n544) );
  NAND2_X1 U592 ( .A1(n545), .A2(n544), .ZN(n546) );
  NOR2_X1 U593 ( .A1(n547), .A2(n546), .ZN(n548) );
  AND2_X1 U594 ( .A1(n549), .A2(n548), .ZN(G160) );
  AND2_X1 U595 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U596 ( .A(G57), .ZN(G237) );
  INV_X1 U597 ( .A(G132), .ZN(G219) );
  INV_X1 U598 ( .A(G82), .ZN(G220) );
  NOR2_X1 U599 ( .A1(G543), .A2(G651), .ZN(n644) );
  NAND2_X1 U600 ( .A1(n644), .A2(G89), .ZN(n550) );
  XNOR2_X1 U601 ( .A(n550), .B(KEYINPUT4), .ZN(n552) );
  XOR2_X1 U602 ( .A(KEYINPUT0), .B(G543), .Z(n655) );
  INV_X1 U603 ( .A(G651), .ZN(n554) );
  NOR2_X1 U604 ( .A1(n655), .A2(n554), .ZN(n647) );
  NAND2_X1 U605 ( .A1(G76), .A2(n647), .ZN(n551) );
  NAND2_X1 U606 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U607 ( .A(n553), .B(KEYINPUT5), .ZN(n560) );
  NAND2_X1 U608 ( .A1(G51), .A2(n653), .ZN(n557) );
  NOR2_X1 U609 ( .A1(G543), .A2(n554), .ZN(n555) );
  XOR2_X2 U610 ( .A(KEYINPUT1), .B(n555), .Z(n659) );
  NAND2_X1 U611 ( .A1(G63), .A2(n659), .ZN(n556) );
  NAND2_X1 U612 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U613 ( .A(KEYINPUT6), .B(n558), .Z(n559) );
  NAND2_X1 U614 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U615 ( .A(n561), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U616 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U617 ( .A1(G7), .A2(G661), .ZN(n562) );
  XNOR2_X1 U618 ( .A(n562), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U619 ( .A(G223), .B(KEYINPUT70), .Z(n835) );
  NAND2_X1 U620 ( .A1(n835), .A2(G567), .ZN(n563) );
  XOR2_X1 U621 ( .A(KEYINPUT11), .B(n563), .Z(G234) );
  NAND2_X1 U622 ( .A1(G81), .A2(n644), .ZN(n564) );
  XNOR2_X1 U623 ( .A(n564), .B(KEYINPUT72), .ZN(n565) );
  XNOR2_X1 U624 ( .A(n565), .B(KEYINPUT12), .ZN(n567) );
  NAND2_X1 U625 ( .A1(G68), .A2(n647), .ZN(n566) );
  NAND2_X1 U626 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U627 ( .A(KEYINPUT13), .B(n568), .Z(n572) );
  NAND2_X1 U628 ( .A1(G56), .A2(n659), .ZN(n569) );
  XNOR2_X1 U629 ( .A(n569), .B(KEYINPUT14), .ZN(n570) );
  XNOR2_X1 U630 ( .A(n570), .B(KEYINPUT71), .ZN(n571) );
  NOR2_X1 U631 ( .A1(n572), .A2(n571), .ZN(n574) );
  NAND2_X1 U632 ( .A1(n653), .A2(G43), .ZN(n573) );
  NAND2_X1 U633 ( .A1(n574), .A2(n573), .ZN(n982) );
  INV_X1 U634 ( .A(G860), .ZN(n603) );
  OR2_X1 U635 ( .A1(n982), .A2(n603), .ZN(G153) );
  NAND2_X1 U636 ( .A1(G52), .A2(n653), .ZN(n576) );
  NAND2_X1 U637 ( .A1(G64), .A2(n659), .ZN(n575) );
  NAND2_X1 U638 ( .A1(n576), .A2(n575), .ZN(n581) );
  NAND2_X1 U639 ( .A1(G90), .A2(n644), .ZN(n578) );
  NAND2_X1 U640 ( .A1(G77), .A2(n647), .ZN(n577) );
  NAND2_X1 U641 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U642 ( .A(KEYINPUT9), .B(n579), .Z(n580) );
  NOR2_X1 U643 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U644 ( .A(KEYINPUT69), .B(n582), .Z(G171) );
  INV_X1 U645 ( .A(G171), .ZN(G301) );
  NAND2_X1 U646 ( .A1(G868), .A2(G301), .ZN(n593) );
  NAND2_X1 U647 ( .A1(G54), .A2(n653), .ZN(n584) );
  NAND2_X1 U648 ( .A1(G79), .A2(n647), .ZN(n583) );
  NAND2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n590) );
  NAND2_X1 U650 ( .A1(n659), .A2(G66), .ZN(n585) );
  XOR2_X1 U651 ( .A(KEYINPUT73), .B(n585), .Z(n587) );
  NAND2_X1 U652 ( .A1(n644), .A2(G92), .ZN(n586) );
  NAND2_X1 U653 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U654 ( .A(KEYINPUT74), .B(n588), .ZN(n589) );
  NOR2_X1 U655 ( .A1(n590), .A2(n589), .ZN(n591) );
  INV_X1 U656 ( .A(G868), .ZN(n600) );
  NAND2_X1 U657 ( .A1(n999), .A2(n600), .ZN(n592) );
  NAND2_X1 U658 ( .A1(n593), .A2(n592), .ZN(G284) );
  NAND2_X1 U659 ( .A1(G53), .A2(n653), .ZN(n595) );
  NAND2_X1 U660 ( .A1(G65), .A2(n659), .ZN(n594) );
  NAND2_X1 U661 ( .A1(n595), .A2(n594), .ZN(n599) );
  NAND2_X1 U662 ( .A1(G91), .A2(n644), .ZN(n597) );
  NAND2_X1 U663 ( .A1(G78), .A2(n647), .ZN(n596) );
  NAND2_X1 U664 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U665 ( .A1(n599), .A2(n598), .ZN(n981) );
  INV_X1 U666 ( .A(n981), .ZN(G299) );
  NOR2_X1 U667 ( .A1(G286), .A2(n600), .ZN(n602) );
  NOR2_X1 U668 ( .A1(G868), .A2(G299), .ZN(n601) );
  NOR2_X1 U669 ( .A1(n602), .A2(n601), .ZN(G297) );
  NAND2_X1 U670 ( .A1(n603), .A2(G559), .ZN(n604) );
  INV_X1 U671 ( .A(n999), .ZN(n620) );
  NAND2_X1 U672 ( .A1(n604), .A2(n620), .ZN(n605) );
  XNOR2_X1 U673 ( .A(n605), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U674 ( .A1(G868), .A2(n982), .ZN(n608) );
  NAND2_X1 U675 ( .A1(n620), .A2(G868), .ZN(n606) );
  NOR2_X1 U676 ( .A1(G559), .A2(n606), .ZN(n607) );
  NOR2_X1 U677 ( .A1(n608), .A2(n607), .ZN(G282) );
  XNOR2_X1 U678 ( .A(G2100), .B(KEYINPUT77), .ZN(n619) );
  NAND2_X1 U679 ( .A1(G99), .A2(n896), .ZN(n610) );
  NAND2_X1 U680 ( .A1(G111), .A2(n900), .ZN(n609) );
  NAND2_X1 U681 ( .A1(n610), .A2(n609), .ZN(n617) );
  NAND2_X1 U682 ( .A1(G135), .A2(n897), .ZN(n611) );
  XNOR2_X1 U683 ( .A(n611), .B(KEYINPUT76), .ZN(n615) );
  XOR2_X1 U684 ( .A(KEYINPUT18), .B(KEYINPUT75), .Z(n613) );
  NAND2_X1 U685 ( .A1(G123), .A2(n901), .ZN(n612) );
  XNOR2_X1 U686 ( .A(n613), .B(n612), .ZN(n614) );
  NAND2_X1 U687 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U688 ( .A1(n617), .A2(n616), .ZN(n935) );
  XNOR2_X1 U689 ( .A(n935), .B(G2096), .ZN(n618) );
  NAND2_X1 U690 ( .A1(n619), .A2(n618), .ZN(G156) );
  NAND2_X1 U691 ( .A1(G559), .A2(n620), .ZN(n621) );
  XNOR2_X1 U692 ( .A(n621), .B(n982), .ZN(n671) );
  NOR2_X1 U693 ( .A1(n671), .A2(G860), .ZN(n628) );
  NAND2_X1 U694 ( .A1(G55), .A2(n653), .ZN(n623) );
  NAND2_X1 U695 ( .A1(G67), .A2(n659), .ZN(n622) );
  NAND2_X1 U696 ( .A1(n623), .A2(n622), .ZN(n627) );
  NAND2_X1 U697 ( .A1(G93), .A2(n644), .ZN(n625) );
  NAND2_X1 U698 ( .A1(G80), .A2(n647), .ZN(n624) );
  NAND2_X1 U699 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U700 ( .A1(n627), .A2(n626), .ZN(n668) );
  XNOR2_X1 U701 ( .A(n628), .B(n668), .ZN(G145) );
  NAND2_X1 U702 ( .A1(G88), .A2(n644), .ZN(n630) );
  NAND2_X1 U703 ( .A1(G75), .A2(n647), .ZN(n629) );
  NAND2_X1 U704 ( .A1(n630), .A2(n629), .ZN(n634) );
  NAND2_X1 U705 ( .A1(G50), .A2(n653), .ZN(n632) );
  NAND2_X1 U706 ( .A1(G62), .A2(n659), .ZN(n631) );
  NAND2_X1 U707 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U708 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U709 ( .A(KEYINPUT79), .B(n635), .Z(G166) );
  NAND2_X1 U710 ( .A1(n653), .A2(G47), .ZN(n636) );
  XOR2_X1 U711 ( .A(KEYINPUT67), .B(n636), .Z(n638) );
  NAND2_X1 U712 ( .A1(n659), .A2(G60), .ZN(n637) );
  NAND2_X1 U713 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U714 ( .A(KEYINPUT68), .B(n639), .Z(n643) );
  NAND2_X1 U715 ( .A1(G85), .A2(n644), .ZN(n641) );
  NAND2_X1 U716 ( .A1(G72), .A2(n647), .ZN(n640) );
  AND2_X1 U717 ( .A1(n641), .A2(n640), .ZN(n642) );
  NAND2_X1 U718 ( .A1(n643), .A2(n642), .ZN(G290) );
  NAND2_X1 U719 ( .A1(G61), .A2(n659), .ZN(n646) );
  NAND2_X1 U720 ( .A1(G86), .A2(n644), .ZN(n645) );
  NAND2_X1 U721 ( .A1(n646), .A2(n645), .ZN(n650) );
  NAND2_X1 U722 ( .A1(n647), .A2(G73), .ZN(n648) );
  XOR2_X1 U723 ( .A(KEYINPUT2), .B(n648), .Z(n649) );
  NOR2_X1 U724 ( .A1(n650), .A2(n649), .ZN(n652) );
  NAND2_X1 U725 ( .A1(n653), .A2(G48), .ZN(n651) );
  NAND2_X1 U726 ( .A1(n652), .A2(n651), .ZN(G305) );
  NAND2_X1 U727 ( .A1(G49), .A2(n653), .ZN(n654) );
  XNOR2_X1 U728 ( .A(n654), .B(KEYINPUT78), .ZN(n661) );
  NAND2_X1 U729 ( .A1(G74), .A2(G651), .ZN(n657) );
  NAND2_X1 U730 ( .A1(G87), .A2(n655), .ZN(n656) );
  NAND2_X1 U731 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U732 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U733 ( .A1(n661), .A2(n660), .ZN(G288) );
  NOR2_X1 U734 ( .A1(G868), .A2(n668), .ZN(n662) );
  XOR2_X1 U735 ( .A(n662), .B(KEYINPUT82), .Z(n674) );
  XOR2_X1 U736 ( .A(KEYINPUT81), .B(KEYINPUT19), .Z(n664) );
  XNOR2_X1 U737 ( .A(n981), .B(KEYINPUT80), .ZN(n663) );
  XNOR2_X1 U738 ( .A(n664), .B(n663), .ZN(n667) );
  XNOR2_X1 U739 ( .A(G166), .B(G290), .ZN(n665) );
  XNOR2_X1 U740 ( .A(n665), .B(G305), .ZN(n666) );
  XNOR2_X1 U741 ( .A(n667), .B(n666), .ZN(n670) );
  XNOR2_X1 U742 ( .A(G288), .B(n668), .ZN(n669) );
  XNOR2_X1 U743 ( .A(n670), .B(n669), .ZN(n918) );
  XNOR2_X1 U744 ( .A(n918), .B(n671), .ZN(n672) );
  NAND2_X1 U745 ( .A1(G868), .A2(n672), .ZN(n673) );
  NAND2_X1 U746 ( .A1(n674), .A2(n673), .ZN(G295) );
  NAND2_X1 U747 ( .A1(G2078), .A2(G2084), .ZN(n675) );
  XOR2_X1 U748 ( .A(KEYINPUT20), .B(n675), .Z(n676) );
  NAND2_X1 U749 ( .A1(G2090), .A2(n676), .ZN(n677) );
  XNOR2_X1 U750 ( .A(KEYINPUT21), .B(n677), .ZN(n678) );
  NAND2_X1 U751 ( .A1(n678), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U752 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U753 ( .A1(G220), .A2(G219), .ZN(n679) );
  XOR2_X1 U754 ( .A(KEYINPUT22), .B(n679), .Z(n680) );
  NOR2_X1 U755 ( .A1(G218), .A2(n680), .ZN(n681) );
  NAND2_X1 U756 ( .A1(G96), .A2(n681), .ZN(n839) );
  NAND2_X1 U757 ( .A1(G2106), .A2(n839), .ZN(n685) );
  NAND2_X1 U758 ( .A1(G69), .A2(G120), .ZN(n682) );
  NOR2_X1 U759 ( .A1(G237), .A2(n682), .ZN(n683) );
  NAND2_X1 U760 ( .A1(G108), .A2(n683), .ZN(n840) );
  NAND2_X1 U761 ( .A1(G567), .A2(n840), .ZN(n684) );
  NAND2_X1 U762 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U763 ( .A(KEYINPUT83), .B(n686), .ZN(G319) );
  INV_X1 U764 ( .A(G319), .ZN(n688) );
  NAND2_X1 U765 ( .A1(G661), .A2(G483), .ZN(n687) );
  NOR2_X1 U766 ( .A1(n688), .A2(n687), .ZN(n838) );
  NAND2_X1 U767 ( .A1(n838), .A2(G36), .ZN(G176) );
  XOR2_X1 U768 ( .A(KEYINPUT86), .B(G166), .Z(G303) );
  NOR2_X1 U769 ( .A1(G1981), .A2(G305), .ZN(n689) );
  XNOR2_X1 U770 ( .A(KEYINPUT24), .B(n689), .ZN(n691) );
  INV_X1 U771 ( .A(n785), .ZN(n690) );
  NAND2_X1 U772 ( .A1(G160), .A2(G40), .ZN(n784) );
  NOR2_X2 U773 ( .A1(n690), .A2(n784), .ZN(n707) );
  NAND2_X1 U774 ( .A1(n743), .A2(G8), .ZN(n756) );
  INV_X1 U775 ( .A(n756), .ZN(n771) );
  NAND2_X1 U776 ( .A1(n691), .A2(n771), .ZN(n758) );
  NOR2_X1 U777 ( .A1(G2084), .A2(n743), .ZN(n726) );
  NAND2_X1 U778 ( .A1(G8), .A2(n726), .ZN(n741) );
  NOR2_X1 U779 ( .A1(G1966), .A2(n756), .ZN(n739) );
  XOR2_X1 U780 ( .A(G2078), .B(KEYINPUT25), .Z(n961) );
  NOR2_X1 U781 ( .A1(n961), .A2(n743), .ZN(n692) );
  XOR2_X1 U782 ( .A(KEYINPUT94), .B(n692), .Z(n695) );
  NOR2_X1 U783 ( .A1(n707), .A2(G1961), .ZN(n693) );
  XNOR2_X1 U784 ( .A(KEYINPUT93), .B(n693), .ZN(n694) );
  NAND2_X1 U785 ( .A1(n695), .A2(n694), .ZN(n730) );
  NAND2_X1 U786 ( .A1(n730), .A2(G171), .ZN(n725) );
  XNOR2_X1 U787 ( .A(G1996), .B(KEYINPUT98), .ZN(n960) );
  NAND2_X1 U788 ( .A1(n960), .A2(n707), .ZN(n696) );
  XNOR2_X1 U789 ( .A(n696), .B(KEYINPUT26), .ZN(n698) );
  NAND2_X1 U790 ( .A1(n743), .A2(G1341), .ZN(n697) );
  NAND2_X1 U791 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U792 ( .A1(n982), .A2(n699), .ZN(n703) );
  NAND2_X1 U793 ( .A1(G1348), .A2(n743), .ZN(n701) );
  NAND2_X1 U794 ( .A1(G2067), .A2(n707), .ZN(n700) );
  NAND2_X1 U795 ( .A1(n701), .A2(n700), .ZN(n704) );
  NOR2_X1 U796 ( .A1(n999), .A2(n704), .ZN(n702) );
  OR2_X1 U797 ( .A1(n703), .A2(n702), .ZN(n706) );
  NAND2_X1 U798 ( .A1(n999), .A2(n704), .ZN(n705) );
  NAND2_X1 U799 ( .A1(n706), .A2(n705), .ZN(n716) );
  NAND2_X1 U800 ( .A1(G2072), .A2(n707), .ZN(n708) );
  XNOR2_X1 U801 ( .A(n708), .B(KEYINPUT95), .ZN(n710) );
  INV_X1 U802 ( .A(KEYINPUT27), .ZN(n709) );
  XNOR2_X1 U803 ( .A(n710), .B(n709), .ZN(n714) );
  INV_X1 U804 ( .A(KEYINPUT96), .ZN(n712) );
  NAND2_X1 U805 ( .A1(G1956), .A2(n743), .ZN(n711) );
  XNOR2_X1 U806 ( .A(n712), .B(n711), .ZN(n713) );
  NOR2_X1 U807 ( .A1(n714), .A2(n713), .ZN(n717) );
  NAND2_X1 U808 ( .A1(n981), .A2(n717), .ZN(n715) );
  NAND2_X1 U809 ( .A1(n716), .A2(n715), .ZN(n721) );
  NOR2_X1 U810 ( .A1(n717), .A2(n981), .ZN(n719) );
  XNOR2_X1 U811 ( .A(KEYINPUT97), .B(KEYINPUT28), .ZN(n718) );
  XNOR2_X1 U812 ( .A(n719), .B(n718), .ZN(n720) );
  NAND2_X1 U813 ( .A1(n721), .A2(n720), .ZN(n723) );
  XNOR2_X1 U814 ( .A(KEYINPUT29), .B(KEYINPUT99), .ZN(n722) );
  XNOR2_X1 U815 ( .A(n723), .B(n722), .ZN(n724) );
  NAND2_X1 U816 ( .A1(n725), .A2(n724), .ZN(n736) );
  INV_X1 U817 ( .A(KEYINPUT31), .ZN(n734) );
  NOR2_X1 U818 ( .A1(n739), .A2(n726), .ZN(n727) );
  NAND2_X1 U819 ( .A1(G8), .A2(n727), .ZN(n728) );
  XNOR2_X1 U820 ( .A(n728), .B(KEYINPUT30), .ZN(n729) );
  NOR2_X1 U821 ( .A1(G168), .A2(n729), .ZN(n732) );
  NOR2_X1 U822 ( .A1(G171), .A2(n730), .ZN(n731) );
  XNOR2_X1 U823 ( .A(n734), .B(n733), .ZN(n735) );
  NAND2_X1 U824 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U825 ( .A(n737), .B(KEYINPUT100), .ZN(n742) );
  INV_X1 U826 ( .A(n742), .ZN(n738) );
  NOR2_X1 U827 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U828 ( .A1(n741), .A2(n740), .ZN(n759) );
  NAND2_X1 U829 ( .A1(n742), .A2(G286), .ZN(n750) );
  INV_X1 U830 ( .A(G8), .ZN(n748) );
  NOR2_X1 U831 ( .A1(G1971), .A2(n756), .ZN(n745) );
  NOR2_X1 U832 ( .A1(G2090), .A2(n743), .ZN(n744) );
  NOR2_X1 U833 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U834 ( .A1(G303), .A2(n746), .ZN(n747) );
  OR2_X1 U835 ( .A1(n748), .A2(n747), .ZN(n749) );
  AND2_X1 U836 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U837 ( .A(n751), .B(KEYINPUT32), .ZN(n761) );
  NAND2_X1 U838 ( .A1(n759), .A2(n761), .ZN(n754) );
  NOR2_X1 U839 ( .A1(G2090), .A2(G303), .ZN(n752) );
  NAND2_X1 U840 ( .A1(G8), .A2(n752), .ZN(n753) );
  NAND2_X1 U841 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U842 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U843 ( .A1(n758), .A2(n757), .ZN(n783) );
  NAND2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n992) );
  AND2_X1 U845 ( .A1(n759), .A2(n992), .ZN(n760) );
  NAND2_X1 U846 ( .A1(n761), .A2(n760), .ZN(n765) );
  INV_X1 U847 ( .A(n992), .ZN(n763) );
  NOR2_X1 U848 ( .A1(G1976), .A2(G288), .ZN(n768) );
  NOR2_X1 U849 ( .A1(G303), .A2(G1971), .ZN(n762) );
  NOR2_X1 U850 ( .A1(n768), .A2(n762), .ZN(n993) );
  OR2_X1 U851 ( .A1(n763), .A2(n993), .ZN(n764) );
  NAND2_X1 U852 ( .A1(n765), .A2(n764), .ZN(n767) );
  XNOR2_X1 U853 ( .A(n767), .B(n766), .ZN(n775) );
  INV_X1 U854 ( .A(KEYINPUT33), .ZN(n777) );
  NAND2_X1 U855 ( .A1(n771), .A2(n768), .ZN(n769) );
  NOR2_X1 U856 ( .A1(n777), .A2(n769), .ZN(n770) );
  XOR2_X1 U857 ( .A(n770), .B(KEYINPUT102), .Z(n776) );
  AND2_X1 U858 ( .A1(n771), .A2(n776), .ZN(n773) );
  XNOR2_X1 U859 ( .A(G1981), .B(G305), .ZN(n990) );
  INV_X1 U860 ( .A(n990), .ZN(n772) );
  AND2_X1 U861 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U862 ( .A1(n775), .A2(n774), .ZN(n781) );
  INV_X1 U863 ( .A(n776), .ZN(n778) );
  OR2_X1 U864 ( .A1(n778), .A2(n777), .ZN(n779) );
  OR2_X1 U865 ( .A1(n990), .A2(n779), .ZN(n780) );
  NAND2_X1 U866 ( .A1(n781), .A2(n780), .ZN(n782) );
  NOR2_X1 U867 ( .A1(n783), .A2(n782), .ZN(n817) );
  NOR2_X1 U868 ( .A1(n785), .A2(n784), .ZN(n830) );
  NAND2_X1 U869 ( .A1(G104), .A2(n896), .ZN(n787) );
  NAND2_X1 U870 ( .A1(G140), .A2(n897), .ZN(n786) );
  NAND2_X1 U871 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U872 ( .A(KEYINPUT34), .B(n788), .ZN(n794) );
  NAND2_X1 U873 ( .A1(G116), .A2(n900), .ZN(n790) );
  NAND2_X1 U874 ( .A1(G128), .A2(n901), .ZN(n789) );
  NAND2_X1 U875 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U876 ( .A(KEYINPUT35), .B(n791), .ZN(n792) );
  XNOR2_X1 U877 ( .A(KEYINPUT87), .B(n792), .ZN(n793) );
  NOR2_X1 U878 ( .A1(n794), .A2(n793), .ZN(n795) );
  XNOR2_X1 U879 ( .A(n795), .B(KEYINPUT36), .ZN(n796) );
  XNOR2_X1 U880 ( .A(n796), .B(KEYINPUT88), .ZN(n893) );
  XNOR2_X1 U881 ( .A(G2067), .B(KEYINPUT37), .ZN(n828) );
  NOR2_X1 U882 ( .A1(n893), .A2(n828), .ZN(n931) );
  NAND2_X1 U883 ( .A1(n830), .A2(n931), .ZN(n797) );
  XOR2_X1 U884 ( .A(KEYINPUT89), .B(n797), .Z(n826) );
  NAND2_X1 U885 ( .A1(G95), .A2(n896), .ZN(n799) );
  NAND2_X1 U886 ( .A1(G131), .A2(n897), .ZN(n798) );
  NAND2_X1 U887 ( .A1(n799), .A2(n798), .ZN(n800) );
  XOR2_X1 U888 ( .A(KEYINPUT90), .B(n800), .Z(n804) );
  NAND2_X1 U889 ( .A1(n901), .A2(G119), .ZN(n802) );
  NAND2_X1 U890 ( .A1(G107), .A2(n900), .ZN(n801) );
  AND2_X1 U891 ( .A1(n802), .A2(n801), .ZN(n803) );
  NAND2_X1 U892 ( .A1(n804), .A2(n803), .ZN(n892) );
  NAND2_X1 U893 ( .A1(n892), .A2(G1991), .ZN(n814) );
  NAND2_X1 U894 ( .A1(G117), .A2(n900), .ZN(n806) );
  NAND2_X1 U895 ( .A1(G129), .A2(n901), .ZN(n805) );
  NAND2_X1 U896 ( .A1(n806), .A2(n805), .ZN(n809) );
  NAND2_X1 U897 ( .A1(n896), .A2(G105), .ZN(n807) );
  XOR2_X1 U898 ( .A(KEYINPUT38), .B(n807), .Z(n808) );
  NOR2_X1 U899 ( .A1(n809), .A2(n808), .ZN(n810) );
  XOR2_X1 U900 ( .A(KEYINPUT91), .B(n810), .Z(n812) );
  NAND2_X1 U901 ( .A1(n897), .A2(G141), .ZN(n811) );
  NAND2_X1 U902 ( .A1(n812), .A2(n811), .ZN(n890) );
  NAND2_X1 U903 ( .A1(G1996), .A2(n890), .ZN(n813) );
  NAND2_X1 U904 ( .A1(n814), .A2(n813), .ZN(n933) );
  AND2_X1 U905 ( .A1(n933), .A2(n830), .ZN(n823) );
  XOR2_X1 U906 ( .A(KEYINPUT92), .B(n823), .Z(n815) );
  XNOR2_X1 U907 ( .A(n818), .B(KEYINPUT103), .ZN(n820) );
  XNOR2_X1 U908 ( .A(G1986), .B(G290), .ZN(n988) );
  NAND2_X1 U909 ( .A1(n988), .A2(n830), .ZN(n819) );
  NAND2_X1 U910 ( .A1(n820), .A2(n819), .ZN(n833) );
  NOR2_X1 U911 ( .A1(G1996), .A2(n890), .ZN(n943) );
  NOR2_X1 U912 ( .A1(G1991), .A2(n892), .ZN(n939) );
  NOR2_X1 U913 ( .A1(G1986), .A2(G290), .ZN(n821) );
  NOR2_X1 U914 ( .A1(n939), .A2(n821), .ZN(n822) );
  NOR2_X1 U915 ( .A1(n823), .A2(n822), .ZN(n824) );
  NOR2_X1 U916 ( .A1(n943), .A2(n824), .ZN(n825) );
  XNOR2_X1 U917 ( .A(n825), .B(KEYINPUT39), .ZN(n827) );
  NAND2_X1 U918 ( .A1(n827), .A2(n826), .ZN(n829) );
  NAND2_X1 U919 ( .A1(n893), .A2(n828), .ZN(n930) );
  NAND2_X1 U920 ( .A1(n829), .A2(n930), .ZN(n831) );
  NAND2_X1 U921 ( .A1(n831), .A2(n830), .ZN(n832) );
  NAND2_X1 U922 ( .A1(n833), .A2(n832), .ZN(n834) );
  XNOR2_X1 U923 ( .A(KEYINPUT40), .B(n834), .ZN(G329) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n835), .ZN(G217) );
  AND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n836) );
  NAND2_X1 U926 ( .A1(G661), .A2(n836), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n837) );
  NAND2_X1 U928 ( .A1(n838), .A2(n837), .ZN(G188) );
  XNOR2_X1 U929 ( .A(G96), .B(KEYINPUT107), .ZN(G221) );
  INV_X1 U931 ( .A(G120), .ZN(G236) );
  INV_X1 U932 ( .A(G69), .ZN(G235) );
  NOR2_X1 U933 ( .A1(n840), .A2(n839), .ZN(G325) );
  INV_X1 U934 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U935 ( .A(G2443), .B(G2451), .ZN(n850) );
  XOR2_X1 U936 ( .A(G2446), .B(G2454), .Z(n842) );
  XNOR2_X1 U937 ( .A(KEYINPUT104), .B(G2435), .ZN(n841) );
  XNOR2_X1 U938 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U939 ( .A(KEYINPUT105), .B(G2438), .Z(n844) );
  XNOR2_X1 U940 ( .A(G1341), .B(G1348), .ZN(n843) );
  XNOR2_X1 U941 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U942 ( .A(n846), .B(n845), .Z(n848) );
  XNOR2_X1 U943 ( .A(G2427), .B(G2430), .ZN(n847) );
  XNOR2_X1 U944 ( .A(n848), .B(n847), .ZN(n849) );
  XNOR2_X1 U945 ( .A(n850), .B(n849), .ZN(n851) );
  NAND2_X1 U946 ( .A1(n851), .A2(G14), .ZN(n852) );
  XOR2_X1 U947 ( .A(KEYINPUT106), .B(n852), .Z(G401) );
  XOR2_X1 U948 ( .A(G1971), .B(G1956), .Z(n854) );
  XNOR2_X1 U949 ( .A(G1996), .B(G1991), .ZN(n853) );
  XNOR2_X1 U950 ( .A(n854), .B(n853), .ZN(n864) );
  XOR2_X1 U951 ( .A(KEYINPUT109), .B(KEYINPUT41), .Z(n856) );
  XNOR2_X1 U952 ( .A(G1961), .B(G2474), .ZN(n855) );
  XNOR2_X1 U953 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U954 ( .A(G1976), .B(G1981), .Z(n858) );
  XNOR2_X1 U955 ( .A(G1986), .B(G1966), .ZN(n857) );
  XNOR2_X1 U956 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U957 ( .A(n860), .B(n859), .Z(n862) );
  XNOR2_X1 U958 ( .A(KEYINPUT111), .B(KEYINPUT110), .ZN(n861) );
  XNOR2_X1 U959 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U960 ( .A(n864), .B(n863), .Z(G229) );
  XOR2_X1 U961 ( .A(G2100), .B(KEYINPUT43), .Z(n866) );
  XNOR2_X1 U962 ( .A(G2067), .B(G2678), .ZN(n865) );
  XNOR2_X1 U963 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U964 ( .A(n867), .B(KEYINPUT108), .Z(n869) );
  XNOR2_X1 U965 ( .A(G2072), .B(G2090), .ZN(n868) );
  XNOR2_X1 U966 ( .A(n869), .B(n868), .ZN(n873) );
  XOR2_X1 U967 ( .A(KEYINPUT42), .B(G2096), .Z(n871) );
  XNOR2_X1 U968 ( .A(G2078), .B(G2084), .ZN(n870) );
  XNOR2_X1 U969 ( .A(n871), .B(n870), .ZN(n872) );
  XNOR2_X1 U970 ( .A(n873), .B(n872), .ZN(G227) );
  NAND2_X1 U971 ( .A1(G124), .A2(n901), .ZN(n874) );
  XNOR2_X1 U972 ( .A(n874), .B(KEYINPUT44), .ZN(n876) );
  NAND2_X1 U973 ( .A1(G136), .A2(n897), .ZN(n875) );
  NAND2_X1 U974 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U975 ( .A(KEYINPUT112), .B(n877), .Z(n879) );
  NAND2_X1 U976 ( .A1(n896), .A2(G100), .ZN(n878) );
  NAND2_X1 U977 ( .A1(n879), .A2(n878), .ZN(n882) );
  NAND2_X1 U978 ( .A1(G112), .A2(n900), .ZN(n880) );
  XNOR2_X1 U979 ( .A(KEYINPUT113), .B(n880), .ZN(n881) );
  NOR2_X1 U980 ( .A1(n882), .A2(n881), .ZN(G162) );
  NAND2_X1 U981 ( .A1(G118), .A2(n900), .ZN(n884) );
  NAND2_X1 U982 ( .A1(G130), .A2(n901), .ZN(n883) );
  NAND2_X1 U983 ( .A1(n884), .A2(n883), .ZN(n889) );
  NAND2_X1 U984 ( .A1(G106), .A2(n896), .ZN(n886) );
  NAND2_X1 U985 ( .A1(G142), .A2(n897), .ZN(n885) );
  NAND2_X1 U986 ( .A1(n886), .A2(n885), .ZN(n887) );
  XOR2_X1 U987 ( .A(n887), .B(KEYINPUT45), .Z(n888) );
  NOR2_X1 U988 ( .A1(n889), .A2(n888), .ZN(n891) );
  XNOR2_X1 U989 ( .A(n891), .B(n890), .ZN(n916) );
  XNOR2_X1 U990 ( .A(n892), .B(G162), .ZN(n895) );
  XNOR2_X1 U991 ( .A(G164), .B(n893), .ZN(n894) );
  XNOR2_X1 U992 ( .A(n895), .B(n894), .ZN(n909) );
  NAND2_X1 U993 ( .A1(G103), .A2(n896), .ZN(n899) );
  NAND2_X1 U994 ( .A1(G139), .A2(n897), .ZN(n898) );
  NAND2_X1 U995 ( .A1(n899), .A2(n898), .ZN(n906) );
  NAND2_X1 U996 ( .A1(G115), .A2(n900), .ZN(n903) );
  NAND2_X1 U997 ( .A1(G127), .A2(n901), .ZN(n902) );
  NAND2_X1 U998 ( .A1(n903), .A2(n902), .ZN(n904) );
  XOR2_X1 U999 ( .A(KEYINPUT47), .B(n904), .Z(n905) );
  NOR2_X1 U1000 ( .A1(n906), .A2(n905), .ZN(n946) );
  XNOR2_X1 U1001 ( .A(G160), .B(n946), .ZN(n907) );
  XNOR2_X1 U1002 ( .A(n907), .B(n935), .ZN(n908) );
  XOR2_X1 U1003 ( .A(n909), .B(n908), .Z(n914) );
  XOR2_X1 U1004 ( .A(KEYINPUT114), .B(KEYINPUT46), .Z(n911) );
  XNOR2_X1 U1005 ( .A(KEYINPUT115), .B(KEYINPUT116), .ZN(n910) );
  XNOR2_X1 U1006 ( .A(n911), .B(n910), .ZN(n912) );
  XNOR2_X1 U1007 ( .A(KEYINPUT48), .B(n912), .ZN(n913) );
  XNOR2_X1 U1008 ( .A(n914), .B(n913), .ZN(n915) );
  XOR2_X1 U1009 ( .A(n916), .B(n915), .Z(n917) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n917), .ZN(G395) );
  XNOR2_X1 U1011 ( .A(G286), .B(n918), .ZN(n920) );
  XNOR2_X1 U1012 ( .A(n982), .B(G171), .ZN(n919) );
  XNOR2_X1 U1013 ( .A(n920), .B(n919), .ZN(n921) );
  XNOR2_X1 U1014 ( .A(n921), .B(n999), .ZN(n922) );
  NOR2_X1 U1015 ( .A1(G37), .A2(n922), .ZN(G397) );
  NOR2_X1 U1016 ( .A1(G229), .A2(G227), .ZN(n923) );
  XOR2_X1 U1017 ( .A(KEYINPUT49), .B(n923), .Z(n924) );
  NAND2_X1 U1018 ( .A1(G319), .A2(n924), .ZN(n925) );
  NOR2_X1 U1019 ( .A1(G401), .A2(n925), .ZN(n926) );
  XOR2_X1 U1020 ( .A(KEYINPUT117), .B(n926), .Z(n929) );
  NOR2_X1 U1021 ( .A1(G395), .A2(G397), .ZN(n927) );
  XNOR2_X1 U1022 ( .A(KEYINPUT118), .B(n927), .ZN(n928) );
  NAND2_X1 U1023 ( .A1(n929), .A2(n928), .ZN(G225) );
  INV_X1 U1024 ( .A(G225), .ZN(G308) );
  INV_X1 U1025 ( .A(G108), .ZN(G238) );
  INV_X1 U1026 ( .A(n930), .ZN(n932) );
  NOR2_X1 U1027 ( .A1(n932), .A2(n931), .ZN(n941) );
  INV_X1 U1028 ( .A(n933), .ZN(n937) );
  XOR2_X1 U1029 ( .A(G2084), .B(G160), .Z(n934) );
  NOR2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1031 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1032 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1033 ( .A1(n941), .A2(n940), .ZN(n953) );
  XOR2_X1 U1034 ( .A(G2090), .B(G162), .Z(n942) );
  NOR2_X1 U1035 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1036 ( .A(KEYINPUT119), .B(n944), .Z(n945) );
  XOR2_X1 U1037 ( .A(KEYINPUT51), .B(n945), .Z(n951) );
  XOR2_X1 U1038 ( .A(G2072), .B(n946), .Z(n948) );
  XOR2_X1 U1039 ( .A(G164), .B(G2078), .Z(n947) );
  NOR2_X1 U1040 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1041 ( .A(KEYINPUT50), .B(n949), .ZN(n950) );
  NAND2_X1 U1042 ( .A1(n951), .A2(n950), .ZN(n952) );
  NOR2_X1 U1043 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1044 ( .A(KEYINPUT52), .B(n954), .ZN(n955) );
  INV_X1 U1045 ( .A(KEYINPUT55), .ZN(n977) );
  NAND2_X1 U1046 ( .A1(n955), .A2(n977), .ZN(n956) );
  NAND2_X1 U1047 ( .A1(n956), .A2(G29), .ZN(n1038) );
  XNOR2_X1 U1048 ( .A(G2090), .B(G35), .ZN(n971) );
  XNOR2_X1 U1049 ( .A(G2067), .B(G26), .ZN(n958) );
  XNOR2_X1 U1050 ( .A(G1991), .B(G25), .ZN(n957) );
  NOR2_X1 U1051 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1052 ( .A1(G28), .A2(n959), .ZN(n968) );
  XNOR2_X1 U1053 ( .A(n960), .B(G32), .ZN(n963) );
  XNOR2_X1 U1054 ( .A(G27), .B(n961), .ZN(n962) );
  NOR2_X1 U1055 ( .A1(n963), .A2(n962), .ZN(n966) );
  XOR2_X1 U1056 ( .A(G2072), .B(KEYINPUT120), .Z(n964) );
  XNOR2_X1 U1057 ( .A(G33), .B(n964), .ZN(n965) );
  NAND2_X1 U1058 ( .A1(n966), .A2(n965), .ZN(n967) );
  NOR2_X1 U1059 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1060 ( .A(KEYINPUT53), .B(n969), .ZN(n970) );
  NOR2_X1 U1061 ( .A1(n971), .A2(n970), .ZN(n972) );
  XOR2_X1 U1062 ( .A(KEYINPUT121), .B(n972), .Z(n975) );
  XOR2_X1 U1063 ( .A(KEYINPUT54), .B(G34), .Z(n973) );
  XNOR2_X1 U1064 ( .A(G2084), .B(n973), .ZN(n974) );
  NAND2_X1 U1065 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1066 ( .A(n977), .B(n976), .ZN(n979) );
  INV_X1 U1067 ( .A(G29), .ZN(n978) );
  NAND2_X1 U1068 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1069 ( .A1(G11), .A2(n980), .ZN(n1036) );
  XNOR2_X1 U1070 ( .A(G16), .B(KEYINPUT56), .ZN(n1005) );
  XNOR2_X1 U1071 ( .A(n981), .B(G1956), .ZN(n986) );
  XNOR2_X1 U1072 ( .A(n982), .B(G1341), .ZN(n984) );
  XNOR2_X1 U1073 ( .A(G301), .B(G1961), .ZN(n983) );
  NOR2_X1 U1074 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1075 ( .A1(n986), .A2(n985), .ZN(n987) );
  NOR2_X1 U1076 ( .A1(n988), .A2(n987), .ZN(n1003) );
  XOR2_X1 U1077 ( .A(G168), .B(G1966), .Z(n989) );
  NOR2_X1 U1078 ( .A1(n990), .A2(n989), .ZN(n991) );
  XOR2_X1 U1079 ( .A(KEYINPUT57), .B(n991), .Z(n998) );
  NAND2_X1 U1080 ( .A1(n993), .A2(n992), .ZN(n995) );
  AND2_X1 U1081 ( .A1(G303), .A2(G1971), .ZN(n994) );
  NOR2_X1 U1082 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1083 ( .A(n996), .B(KEYINPUT122), .ZN(n997) );
  NAND2_X1 U1084 ( .A1(n998), .A2(n997), .ZN(n1001) );
  XNOR2_X1 U1085 ( .A(G1348), .B(n999), .ZN(n1000) );
  NOR2_X1 U1086 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1087 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1088 ( .A1(n1005), .A2(n1004), .ZN(n1034) );
  INV_X1 U1089 ( .A(G16), .ZN(n1032) );
  XNOR2_X1 U1090 ( .A(KEYINPUT127), .B(KEYINPUT61), .ZN(n1030) );
  XNOR2_X1 U1091 ( .A(KEYINPUT125), .B(G1966), .ZN(n1006) );
  XNOR2_X1 U1092 ( .A(n1006), .B(G21), .ZN(n1028) );
  XOR2_X1 U1093 ( .A(G1961), .B(G5), .Z(n1014) );
  XNOR2_X1 U1094 ( .A(G1971), .B(G22), .ZN(n1008) );
  XNOR2_X1 U1095 ( .A(G1976), .B(G23), .ZN(n1007) );
  NOR2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1097 ( .A(KEYINPUT126), .B(n1009), .Z(n1011) );
  XNOR2_X1 U1098 ( .A(G1986), .B(G24), .ZN(n1010) );
  NOR2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1100 ( .A(KEYINPUT58), .B(n1012), .ZN(n1013) );
  NAND2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1026) );
  XNOR2_X1 U1102 ( .A(G1341), .B(G19), .ZN(n1016) );
  XNOR2_X1 U1103 ( .A(G6), .B(G1981), .ZN(n1015) );
  NOR2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1023) );
  XOR2_X1 U1105 ( .A(KEYINPUT124), .B(G4), .Z(n1018) );
  XNOR2_X1 U1106 ( .A(G1348), .B(KEYINPUT59), .ZN(n1017) );
  XNOR2_X1 U1107 ( .A(n1018), .B(n1017), .ZN(n1019) );
  XOR2_X1 U1108 ( .A(KEYINPUT123), .B(n1019), .Z(n1021) );
  XNOR2_X1 U1109 ( .A(G1956), .B(G20), .ZN(n1020) );
  NOR2_X1 U1110 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1111 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1112 ( .A(KEYINPUT60), .B(n1024), .ZN(n1025) );
  NOR2_X1 U1113 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1114 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1115 ( .A(n1030), .B(n1029), .ZN(n1031) );
  NAND2_X1 U1116 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NAND2_X1 U1117 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NOR2_X1 U1118 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  NAND2_X1 U1119 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  XOR2_X1 U1120 ( .A(KEYINPUT62), .B(n1039), .Z(G311) );
  INV_X1 U1121 ( .A(G311), .ZN(G150) );
endmodule

