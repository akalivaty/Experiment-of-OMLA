//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 0 1 0 1 0 0 0 0 1 0 0 0 0 0 1 0 0 0 0 0 0 1 0 0 1 0 1 0 0 0 0 1 0 0 1 0 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:35 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n817, new_n818, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT81), .ZN(new_n189));
  INV_X1    g003(.A(G469), .ZN(new_n190));
  INV_X1    g004(.A(G902), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G953), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G227), .ZN(new_n194));
  XNOR2_X1  g008(.A(new_n194), .B(KEYINPUT82), .ZN(new_n195));
  XNOR2_X1  g009(.A(G110), .B(G140), .ZN(new_n196));
  XNOR2_X1  g010(.A(new_n195), .B(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G104), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT3), .B1(new_n198), .B2(G107), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT3), .ZN(new_n200));
  INV_X1    g014(.A(G107), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(new_n201), .A3(G104), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n198), .A2(G107), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n199), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G101), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT83), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G101), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n199), .A2(new_n202), .A3(new_n208), .A4(new_n203), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n204), .A2(KEYINPUT83), .A3(G101), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n207), .A2(KEYINPUT4), .A3(new_n209), .A4(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT0), .B(G128), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  OR2_X1    g027(.A1(KEYINPUT64), .A2(G146), .ZN(new_n214));
  NAND2_X1  g028(.A1(KEYINPUT64), .A2(G146), .ZN(new_n215));
  AOI21_X1  g029(.A(G143), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G146), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G143), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n213), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT4), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n204), .A2(new_n221), .A3(G101), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT65), .B1(new_n217), .B2(G143), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT65), .ZN(new_n224));
  INV_X1    g038(.A(G143), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n224), .A2(new_n225), .A3(G146), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n214), .A2(G143), .A3(new_n215), .ZN(new_n228));
  AND2_X1   g042(.A1(KEYINPUT0), .A2(G128), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  AND3_X1   g044(.A1(new_n220), .A2(new_n222), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n211), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n198), .A2(G107), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n201), .A2(G104), .ZN(new_n234));
  OAI21_X1  g048(.A(G101), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  AND2_X1   g049(.A1(new_n209), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G128), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n237), .A2(KEYINPUT1), .ZN(new_n238));
  AND3_X1   g052(.A1(new_n227), .A2(new_n228), .A3(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n237), .B1(new_n218), .B2(KEYINPUT1), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n240), .B1(new_n228), .B2(new_n227), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n236), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT10), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n227), .A2(new_n228), .A3(new_n238), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n237), .B1(new_n228), .B2(KEYINPUT1), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n214), .A2(new_n215), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n219), .B1(new_n247), .B2(new_n225), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n245), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  AND3_X1   g063(.A1(new_n209), .A2(new_n235), .A3(KEYINPUT10), .ZN(new_n250));
  AND3_X1   g064(.A1(new_n249), .A2(KEYINPUT84), .A3(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(KEYINPUT84), .B1(new_n249), .B2(new_n250), .ZN(new_n252));
  OAI211_X1 g066(.A(new_n232), .B(new_n244), .C1(new_n251), .C2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT11), .ZN(new_n254));
  INV_X1    g068(.A(G134), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  OR2_X1    g070(.A1(KEYINPUT68), .A2(G137), .ZN(new_n257));
  NAND2_X1  g071(.A1(KEYINPUT68), .A2(G137), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n255), .A2(G137), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT67), .ZN(new_n261));
  INV_X1    g075(.A(G137), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G134), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n261), .B1(new_n263), .B2(new_n254), .ZN(new_n264));
  AOI211_X1 g078(.A(KEYINPUT67), .B(KEYINPUT11), .C1(new_n262), .C2(G134), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n259), .B(new_n260), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G131), .ZN(new_n267));
  AOI21_X1  g081(.A(G131), .B1(new_n255), .B2(G137), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n259), .B(new_n268), .C1(new_n264), .C2(new_n265), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n253), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n254), .B1(new_n255), .B2(G137), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT67), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n263), .A2(new_n261), .A3(new_n254), .ZN(new_n274));
  AND2_X1   g088(.A1(KEYINPUT68), .A2(G137), .ZN(new_n275));
  NOR2_X1   g089(.A1(KEYINPUT68), .A2(G137), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AOI22_X1  g091(.A1(new_n273), .A2(new_n274), .B1(new_n277), .B2(new_n256), .ZN(new_n278));
  AOI22_X1  g092(.A1(G131), .A2(new_n266), .B1(new_n278), .B2(new_n268), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n249), .A2(new_n250), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT84), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n249), .A2(KEYINPUT84), .A3(new_n250), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n211), .A2(new_n231), .B1(new_n242), .B2(new_n243), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n279), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n197), .B1(new_n271), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n209), .A2(new_n235), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n288), .B(new_n245), .C1(new_n246), .C2(new_n248), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n242), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n270), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT12), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n290), .A2(KEYINPUT12), .A3(new_n270), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n284), .A2(new_n279), .A3(new_n285), .ZN(new_n296));
  INV_X1    g110(.A(new_n197), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(G902), .B1(new_n287), .B2(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n192), .B1(new_n299), .B2(new_n190), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n297), .B1(new_n253), .B2(new_n270), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n301), .A2(new_n286), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n297), .B1(new_n295), .B2(new_n296), .ZN(new_n303));
  OAI21_X1  g117(.A(KEYINPUT85), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AND3_X1   g118(.A1(new_n290), .A2(KEYINPUT12), .A3(new_n270), .ZN(new_n305));
  AOI21_X1  g119(.A(KEYINPUT12), .B1(new_n290), .B2(new_n270), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n197), .B1(new_n271), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT85), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n253), .A2(new_n270), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n310), .A2(new_n296), .A3(new_n297), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n308), .A2(new_n309), .A3(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n304), .A2(new_n312), .A3(G469), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n189), .B1(new_n300), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT20), .ZN(new_n315));
  NOR2_X1   g129(.A1(G475), .A2(G902), .ZN(new_n316));
  XOR2_X1   g130(.A(G113), .B(G122), .Z(new_n317));
  XOR2_X1   g131(.A(KEYINPUT91), .B(G104), .Z(new_n318));
  XOR2_X1   g132(.A(new_n317), .B(new_n318), .Z(new_n319));
  NAND2_X1  g133(.A1(KEYINPUT18), .A2(G131), .ZN(new_n320));
  INV_X1    g134(.A(G237), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(new_n193), .A3(G214), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT88), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n322), .A2(new_n323), .A3(new_n225), .ZN(new_n324));
  NOR2_X1   g138(.A1(G237), .A2(G953), .ZN(new_n325));
  OAI211_X1 g139(.A(new_n325), .B(G214), .C1(KEYINPUT88), .C2(G143), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n320), .B1(new_n327), .B2(KEYINPUT89), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT89), .ZN(new_n329));
  INV_X1    g143(.A(new_n320), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n324), .A2(new_n329), .A3(new_n326), .A4(new_n330), .ZN(new_n331));
  AND2_X1   g145(.A1(KEYINPUT64), .A2(G146), .ZN(new_n332));
  NOR2_X1   g146(.A1(KEYINPUT64), .A2(G146), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(G125), .B(G140), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OR2_X1    g150(.A1(new_n335), .A2(new_n217), .ZN(new_n337));
  AOI22_X1  g151(.A1(new_n328), .A2(new_n331), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n327), .A2(KEYINPUT17), .A3(G131), .ZN(new_n339));
  INV_X1    g153(.A(G140), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G125), .ZN(new_n341));
  INV_X1    g155(.A(G125), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G140), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n341), .A2(new_n343), .A3(KEYINPUT16), .ZN(new_n344));
  OR3_X1    g158(.A1(new_n342), .A2(KEYINPUT16), .A3(G140), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n344), .A2(new_n345), .A3(G146), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n344), .A2(new_n345), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n217), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n339), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(G131), .ZN(new_n350));
  AND3_X1   g164(.A1(new_n324), .A2(new_n350), .A3(new_n326), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n350), .B1(new_n324), .B2(new_n326), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT17), .ZN(new_n354));
  AOI22_X1  g168(.A1(new_n349), .A2(KEYINPUT92), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT92), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n339), .A2(new_n356), .A3(new_n346), .A4(new_n348), .ZN(new_n357));
  AOI211_X1 g171(.A(new_n319), .B(new_n338), .C1(new_n355), .C2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n319), .ZN(new_n359));
  OAI21_X1  g173(.A(KEYINPUT90), .B1(new_n351), .B2(new_n352), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n327), .A2(G131), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT90), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n324), .A2(new_n350), .A3(new_n326), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n335), .B(KEYINPUT19), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n334), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n360), .A2(new_n364), .A3(new_n346), .A4(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n328), .A2(new_n331), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n337), .A2(new_n336), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n359), .B1(new_n367), .B2(new_n370), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n315), .B(new_n316), .C1(new_n358), .C2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(KEYINPUT93), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n338), .B1(new_n355), .B2(new_n357), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n359), .ZN(new_n375));
  INV_X1    g189(.A(new_n371), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT93), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n377), .A2(new_n378), .A3(new_n315), .A4(new_n316), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n371), .B1(new_n374), .B2(new_n359), .ZN(new_n380));
  INV_X1    g194(.A(new_n316), .ZN(new_n381));
  OAI21_X1  g195(.A(KEYINPUT20), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n373), .A2(new_n379), .A3(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n374), .A2(new_n359), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n191), .B1(new_n384), .B2(new_n358), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G475), .ZN(new_n386));
  INV_X1    g200(.A(G478), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n387), .A2(KEYINPUT15), .ZN(new_n388));
  INV_X1    g202(.A(G217), .ZN(new_n389));
  NOR3_X1   g203(.A1(new_n187), .A2(new_n389), .A3(G953), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n225), .A2(G128), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n237), .A2(G143), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n392), .A2(new_n393), .A3(new_n255), .ZN(new_n394));
  INV_X1    g208(.A(G122), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G116), .ZN(new_n396));
  INV_X1    g210(.A(G116), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G122), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n399), .A2(G107), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n201), .B1(new_n396), .B2(new_n398), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n394), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n225), .A2(G128), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT13), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n392), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(KEYINPUT94), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT94), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n407), .B(new_n392), .C1(new_n403), .C2(new_n404), .ZN(new_n408));
  INV_X1    g222(.A(new_n392), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT13), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n406), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n402), .B1(new_n411), .B2(G134), .ZN(new_n412));
  OAI21_X1  g226(.A(G134), .B1(new_n409), .B2(new_n403), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n394), .ZN(new_n414));
  INV_X1    g228(.A(new_n400), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n397), .A2(KEYINPUT14), .A3(G122), .ZN(new_n416));
  OAI211_X1 g230(.A(G107), .B(new_n416), .C1(new_n399), .C2(KEYINPUT14), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n414), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n391), .B1(new_n412), .B2(new_n419), .ZN(new_n420));
  AOI22_X1  g234(.A1(new_n405), .A2(KEYINPUT94), .B1(KEYINPUT13), .B2(new_n409), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n255), .B1(new_n421), .B2(new_n408), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n418), .B(new_n390), .C1(new_n422), .C2(new_n402), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(KEYINPUT95), .B1(new_n424), .B2(new_n191), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT95), .ZN(new_n426));
  AOI211_X1 g240(.A(new_n426), .B(G902), .C1(new_n420), .C2(new_n423), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n388), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(G952), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n429), .A2(G953), .ZN(new_n430));
  INV_X1    g244(.A(G234), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n430), .B1(new_n431), .B2(new_n321), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  AOI211_X1 g247(.A(new_n191), .B(new_n193), .C1(G234), .C2(G237), .ZN(new_n434));
  XNOR2_X1  g248(.A(KEYINPUT21), .B(G898), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(G902), .B1(new_n420), .B2(new_n423), .ZN(new_n438));
  OAI22_X1  g252(.A1(new_n438), .A2(KEYINPUT95), .B1(KEYINPUT15), .B2(new_n387), .ZN(new_n439));
  AND3_X1   g253(.A1(new_n428), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n383), .A2(new_n386), .A3(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(G214), .B1(G237), .B2(G902), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(G210), .B1(G237), .B2(G902), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT69), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n446), .B1(new_n397), .B2(G119), .ZN(new_n447));
  INV_X1    g261(.A(G119), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(KEYINPUT69), .A3(G116), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n397), .A2(G119), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n447), .A2(new_n449), .A3(KEYINPUT5), .A4(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT86), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT5), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n452), .A2(new_n453), .A3(new_n448), .A4(G116), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n453), .A2(new_n448), .A3(G116), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(KEYINPUT86), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n451), .A2(G113), .A3(new_n454), .A4(new_n456), .ZN(new_n457));
  XOR2_X1   g271(.A(KEYINPUT2), .B(G113), .Z(new_n458));
  NAND4_X1  g272(.A1(new_n458), .A2(new_n447), .A3(new_n449), .A4(new_n450), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n236), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(G110), .B(G122), .ZN(new_n461));
  AND3_X1   g275(.A1(new_n204), .A2(KEYINPUT83), .A3(G101), .ZN(new_n462));
  AOI21_X1  g276(.A(KEYINPUT83), .B1(new_n204), .B2(G101), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n209), .A2(KEYINPUT4), .ZN(new_n464));
  NOR3_X1   g278(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n447), .A2(new_n449), .A3(new_n450), .ZN(new_n466));
  XNOR2_X1  g280(.A(KEYINPUT2), .B(G113), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n459), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n222), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n460), .B(new_n461), .C1(new_n465), .C2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n205), .ZN(new_n472));
  AOI22_X1  g286(.A1(new_n472), .A2(new_n221), .B1(new_n459), .B2(new_n468), .ZN(new_n473));
  AND2_X1   g287(.A1(new_n457), .A2(new_n459), .ZN(new_n474));
  AOI22_X1  g288(.A1(new_n211), .A2(new_n473), .B1(new_n474), .B2(new_n236), .ZN(new_n475));
  INV_X1    g289(.A(new_n461), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(KEYINPUT87), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n471), .B(KEYINPUT6), .C1(new_n475), .C2(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n460), .B1(new_n465), .B2(new_n470), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT6), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n479), .A2(KEYINPUT87), .A3(new_n480), .A4(new_n476), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n249), .A2(new_n342), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n193), .A2(G224), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n220), .A2(G125), .A3(new_n230), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n483), .B1(new_n482), .B2(new_n484), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AND3_X1   g301(.A1(new_n478), .A2(new_n481), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n482), .A2(new_n484), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n483), .A2(KEYINPUT7), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n461), .B(KEYINPUT8), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n236), .A2(new_n457), .A3(new_n459), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n236), .B1(new_n459), .B2(new_n457), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n482), .A2(new_n484), .A3(new_n490), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n492), .A2(new_n496), .A3(new_n471), .A4(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n191), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n445), .B1(new_n488), .B2(new_n499), .ZN(new_n500));
  AND2_X1   g314(.A1(new_n498), .A2(new_n191), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n478), .A2(new_n481), .A3(new_n487), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n501), .A2(new_n444), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n443), .B1(new_n500), .B2(new_n503), .ZN(new_n504));
  AND3_X1   g318(.A1(new_n314), .A2(new_n441), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n389), .B1(G234), .B2(new_n191), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT25), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n193), .A2(G221), .A3(G234), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n509), .B(KEYINPUT79), .ZN(new_n510));
  XNOR2_X1  g324(.A(KEYINPUT22), .B(G137), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n510), .B(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n346), .A2(new_n336), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  XOR2_X1   g328(.A(KEYINPUT24), .B(G110), .Z(new_n515));
  INV_X1    g329(.A(KEYINPUT74), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n448), .A2(G128), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n237), .A2(G119), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n237), .A2(G119), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n448), .A2(G128), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n520), .A2(new_n521), .A3(KEYINPUT74), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n515), .B1(new_n519), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n237), .A2(KEYINPUT23), .A3(G119), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n521), .B(new_n524), .C1(new_n517), .C2(KEYINPUT23), .ZN(new_n525));
  XOR2_X1   g339(.A(KEYINPUT76), .B(G110), .Z(new_n526));
  OAI22_X1  g340(.A1(new_n523), .A2(KEYINPUT77), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(KEYINPUT24), .B(G110), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n520), .A2(new_n521), .A3(KEYINPUT74), .ZN(new_n529));
  AOI21_X1  g343(.A(KEYINPUT74), .B1(new_n520), .B2(new_n521), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT77), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n514), .B1(new_n527), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n519), .A2(new_n522), .A3(new_n515), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT75), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT75), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n519), .A2(new_n537), .A3(new_n522), .A4(new_n515), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  AOI22_X1  g353(.A1(new_n348), .A2(new_n346), .B1(G110), .B2(new_n525), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n512), .B1(new_n534), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT78), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n539), .A2(new_n540), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n525), .A2(new_n526), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n545), .B1(new_n531), .B2(new_n532), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n523), .A2(KEYINPUT77), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n513), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n543), .B1(new_n544), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n534), .A2(KEYINPUT78), .A3(new_n541), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n542), .B1(new_n551), .B2(new_n512), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n508), .B1(new_n552), .B2(G902), .ZN(new_n553));
  AND3_X1   g367(.A1(new_n534), .A2(KEYINPUT78), .A3(new_n541), .ZN(new_n554));
  AOI21_X1  g368(.A(KEYINPUT78), .B1(new_n534), .B2(new_n541), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n512), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n542), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n558), .A2(KEYINPUT25), .A3(new_n191), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n507), .B1(new_n553), .B2(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n506), .A2(G902), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n325), .A2(G210), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n564), .B(KEYINPUT27), .ZN(new_n565));
  XNOR2_X1  g379(.A(KEYINPUT26), .B(G101), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n565), .B(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n220), .A2(new_n230), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(G134), .B1(new_n257), .B2(new_n258), .ZN(new_n571));
  INV_X1    g385(.A(new_n263), .ZN(new_n572));
  OAI21_X1  g386(.A(G131), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n269), .A2(new_n573), .ZN(new_n574));
  AOI22_X1  g388(.A1(new_n270), .A2(new_n570), .B1(new_n574), .B2(new_n249), .ZN(new_n575));
  INV_X1    g389(.A(new_n469), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n568), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT66), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n225), .B1(new_n332), .B2(new_n333), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n212), .B1(new_n580), .B2(new_n218), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n578), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n220), .A2(KEYINPUT66), .A3(new_n230), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n270), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n574), .A2(new_n249), .ZN(new_n585));
  AOI21_X1  g399(.A(KEYINPUT30), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NOR3_X1   g400(.A1(new_n332), .A2(new_n333), .A3(new_n225), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT1), .ZN(new_n588));
  OAI21_X1  g402(.A(G128), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n580), .A2(new_n218), .ZN(new_n590));
  AOI22_X1  g404(.A1(new_n334), .A2(G143), .B1(new_n223), .B2(new_n226), .ZN(new_n591));
  AOI22_X1  g405(.A1(new_n589), .A2(new_n590), .B1(new_n591), .B2(new_n238), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n269), .A2(new_n573), .ZN(new_n593));
  OAI21_X1  g407(.A(KEYINPUT30), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n569), .B1(new_n267), .B2(new_n269), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n469), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n577), .B1(new_n586), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(KEYINPUT31), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n582), .A2(new_n583), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n585), .B1(new_n599), .B2(new_n279), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n469), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT28), .ZN(new_n602));
  OAI22_X1  g416(.A1(new_n279), .A2(new_n569), .B1(new_n592), .B2(new_n593), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n602), .B1(new_n603), .B2(new_n469), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n350), .B1(new_n278), .B2(new_n260), .ZN(new_n605));
  INV_X1    g419(.A(new_n269), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n570), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n607), .A2(new_n585), .A3(KEYINPUT28), .A4(new_n576), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n601), .A2(new_n604), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n568), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT31), .ZN(new_n611));
  OAI211_X1 g425(.A(new_n577), .B(new_n611), .C1(new_n586), .C2(new_n596), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n598), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(G472), .A2(G902), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(KEYINPUT70), .B(KEYINPUT32), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT73), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT32), .ZN(new_n619));
  NOR3_X1   g433(.A1(new_n619), .A2(G472), .A3(G902), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n613), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n618), .B1(new_n613), .B2(new_n620), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n617), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT71), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n607), .A2(new_n585), .A3(new_n624), .A4(new_n576), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n592), .A2(new_n593), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n469), .B1(new_n626), .B2(new_n595), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n624), .B1(new_n575), .B2(new_n576), .ZN(new_n629));
  OAI21_X1  g443(.A(KEYINPUT28), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n604), .A2(KEYINPUT29), .A3(new_n567), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT72), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n630), .A2(new_n631), .A3(KEYINPUT72), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n575), .A2(new_n576), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n636), .B1(new_n586), .B2(new_n596), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n568), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT29), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n601), .A2(new_n604), .A3(new_n567), .A4(new_n608), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n634), .A2(new_n191), .A3(new_n635), .A4(new_n641), .ZN(new_n642));
  AND2_X1   g456(.A1(new_n642), .A2(G472), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n563), .B1(new_n623), .B2(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n644), .A2(KEYINPUT80), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT80), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n613), .A2(new_n620), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(KEYINPUT73), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n613), .A2(new_n618), .A3(new_n620), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n642), .A2(G472), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n650), .A2(new_n651), .A3(new_n617), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n646), .B1(new_n652), .B2(new_n563), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n505), .B1(new_n645), .B2(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G101), .ZN(G3));
  NAND2_X1  g469(.A1(new_n613), .A2(new_n191), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(G472), .ZN(new_n657));
  AND2_X1   g471(.A1(new_n657), .A2(new_n615), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n658), .A2(new_n563), .A3(new_n314), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n444), .B1(new_n501), .B2(new_n502), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n443), .B1(new_n660), .B2(KEYINPUT96), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT96), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n500), .A2(new_n662), .A3(new_n503), .ZN(new_n663));
  AND2_X1   g477(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n383), .A2(new_n386), .ZN(new_n665));
  OR2_X1    g479(.A1(new_n438), .A2(G478), .ZN(new_n666));
  OR2_X1    g480(.A1(new_n666), .A2(KEYINPUT98), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(KEYINPUT98), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT33), .ZN(new_n670));
  INV_X1    g484(.A(new_n424), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n670), .B1(new_n671), .B2(KEYINPUT97), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT97), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n424), .A2(new_n673), .A3(KEYINPUT33), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n387), .A2(G902), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n669), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n664), .A2(new_n665), .A3(new_n437), .A4(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n659), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(KEYINPUT34), .B(G104), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G6));
  NAND2_X1  g496(.A1(new_n382), .A2(new_n372), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n386), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n428), .A2(new_n439), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n664), .A2(new_n437), .A3(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n659), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(KEYINPUT99), .ZN(new_n690));
  XOR2_X1   g504(.A(KEYINPUT35), .B(G107), .Z(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G9));
  NOR2_X1   g506(.A1(new_n512), .A2(KEYINPUT36), .ZN(new_n693));
  OR2_X1    g507(.A1(new_n551), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n551), .A2(new_n693), .ZN(new_n695));
  AND3_X1   g509(.A1(new_n694), .A2(new_n561), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g510(.A(KEYINPUT100), .B1(new_n560), .B2(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(KEYINPUT25), .B1(new_n558), .B2(new_n191), .ZN(new_n698));
  AOI211_X1 g512(.A(new_n508), .B(G902), .C1(new_n556), .C2(new_n557), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n506), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT100), .ZN(new_n701));
  INV_X1    g515(.A(new_n696), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n700), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  AND3_X1   g517(.A1(new_n658), .A2(new_n697), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n505), .ZN(new_n705));
  XOR2_X1   g519(.A(KEYINPUT37), .B(G110), .Z(new_n706));
  XOR2_X1   g520(.A(new_n706), .B(KEYINPUT101), .Z(new_n707));
  XNOR2_X1  g521(.A(new_n705), .B(new_n707), .ZN(G12));
  NOR2_X1   g522(.A1(new_n623), .A2(new_n643), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n697), .A2(new_n703), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AND2_X1   g525(.A1(new_n314), .A2(new_n664), .ZN(new_n712));
  INV_X1    g526(.A(G900), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n433), .B1(new_n434), .B2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n683), .A2(new_n685), .A3(new_n386), .A4(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n711), .A2(KEYINPUT102), .A3(new_n712), .A4(new_n717), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n697), .A2(new_n703), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n719), .A2(new_n712), .A3(new_n652), .A4(new_n717), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT102), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G128), .ZN(G30));
  NOR2_X1   g538(.A1(new_n560), .A2(new_n696), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n686), .B1(new_n383), .B2(new_n386), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n725), .A2(new_n442), .A3(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(KEYINPUT104), .ZN(new_n728));
  XOR2_X1   g542(.A(new_n714), .B(KEYINPUT39), .Z(new_n729));
  NAND2_X1  g543(.A1(new_n314), .A2(new_n729), .ZN(new_n730));
  OR2_X1    g544(.A1(new_n730), .A2(KEYINPUT40), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(KEYINPUT40), .ZN(new_n732));
  AOI22_X1  g546(.A1(new_n648), .A2(new_n649), .B1(new_n616), .B2(new_n615), .ZN(new_n733));
  OR3_X1    g547(.A1(new_n628), .A2(new_n629), .A3(new_n567), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n637), .A2(new_n567), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n734), .A2(new_n735), .A3(KEYINPUT103), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n191), .ZN(new_n737));
  AOI21_X1  g551(.A(KEYINPUT103), .B1(new_n734), .B2(new_n735), .ZN(new_n738));
  OAI21_X1  g552(.A(G472), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n733), .A2(new_n739), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n500), .A2(KEYINPUT38), .A3(new_n503), .ZN(new_n741));
  AOI21_X1  g555(.A(KEYINPUT38), .B1(new_n500), .B2(new_n503), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AND2_X1   g557(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n728), .A2(new_n731), .A3(new_n732), .A4(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G143), .ZN(G45));
  NAND3_X1  g560(.A1(new_n665), .A2(new_n678), .A3(new_n715), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n719), .A2(new_n712), .A3(new_n652), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G146), .ZN(G48));
  INV_X1    g564(.A(KEYINPUT106), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n301), .A2(new_n307), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n297), .B1(new_n310), .B2(new_n296), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n191), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(G469), .ZN(new_n755));
  INV_X1    g569(.A(new_n189), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n190), .B(new_n191), .C1(new_n752), .C2(new_n753), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n755), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(KEYINPUT105), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT105), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n755), .A2(new_n760), .A3(new_n756), .A4(new_n757), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n652), .A2(new_n563), .A3(new_n759), .A4(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n751), .B1(new_n762), .B2(new_n679), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n560), .A2(new_n562), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n764), .B1(new_n733), .B2(new_n651), .ZN(new_n765));
  INV_X1    g579(.A(new_n679), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n759), .A2(new_n761), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n765), .A2(new_n766), .A3(new_n768), .A4(KEYINPUT106), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n763), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(KEYINPUT41), .B(G113), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n770), .B(new_n771), .ZN(G15));
  NOR3_X1   g586(.A1(new_n644), .A2(new_n767), .A3(new_n688), .ZN(new_n773));
  XNOR2_X1  g587(.A(KEYINPUT107), .B(G116), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n773), .B(new_n774), .ZN(G18));
  AND3_X1   g589(.A1(new_n755), .A2(new_n756), .A3(new_n757), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n664), .A2(new_n776), .A3(new_n441), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n709), .A2(new_n777), .A3(new_n710), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(new_n448), .ZN(G21));
  NAND2_X1  g593(.A1(new_n598), .A2(new_n612), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n567), .B1(new_n630), .B2(new_n604), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  AOI22_X1  g596(.A1(new_n782), .A2(new_n614), .B1(new_n656), .B2(G472), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n783), .A2(new_n664), .A3(new_n563), .A4(new_n726), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n759), .A2(new_n437), .A3(new_n761), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT108), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  OAI21_X1  g602(.A(KEYINPUT108), .B1(new_n784), .B2(new_n785), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G122), .ZN(G24));
  NAND2_X1  g605(.A1(new_n782), .A2(new_n614), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n657), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n725), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n664), .A2(new_n776), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n794), .A2(new_n748), .A3(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G125), .ZN(G27));
  INV_X1    g611(.A(KEYINPUT42), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n500), .A2(new_n442), .A3(new_n503), .ZN(new_n799));
  INV_X1    g613(.A(new_n192), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n308), .A2(G469), .A3(new_n311), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n757), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n799), .A2(new_n802), .A3(new_n756), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n803), .B(new_n563), .C1(new_n623), .C2(new_n643), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n798), .B1(new_n804), .B2(new_n747), .ZN(new_n805));
  INV_X1    g619(.A(new_n647), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT32), .B1(new_n613), .B2(new_n614), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT109), .ZN(new_n808));
  OR3_X1    g622(.A1(new_n806), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n808), .B1(new_n806), .B2(new_n807), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n809), .A2(new_n810), .A3(new_n651), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n799), .A2(new_n802), .A3(new_n756), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n747), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n811), .A2(new_n813), .A3(KEYINPUT42), .A4(new_n563), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n805), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(G131), .ZN(G33));
  XOR2_X1   g630(.A(new_n716), .B(KEYINPUT110), .Z(new_n817));
  NAND3_X1  g631(.A1(new_n765), .A2(new_n803), .A3(new_n817), .ZN(new_n818));
  XOR2_X1   g632(.A(KEYINPUT111), .B(G134), .Z(new_n819));
  XNOR2_X1  g633(.A(new_n818), .B(new_n819), .ZN(G36));
  OR3_X1    g634(.A1(new_n658), .A2(KEYINPUT113), .A3(new_n725), .ZN(new_n821));
  OAI21_X1  g635(.A(KEYINPUT113), .B1(new_n658), .B2(new_n725), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AOI22_X1  g637(.A1(new_n667), .A2(new_n668), .B1(new_n675), .B2(new_n676), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n665), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(KEYINPUT43), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT43), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n827), .B1(new_n665), .B2(new_n824), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n823), .A2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n799), .B1(new_n831), .B2(KEYINPUT44), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n823), .A2(KEYINPUT44), .A3(new_n829), .ZN(new_n833));
  AOI21_X1  g647(.A(KEYINPUT45), .B1(new_n304), .B2(new_n312), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n308), .A2(KEYINPUT45), .A3(new_n311), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(G469), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n800), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT46), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n839), .A2(KEYINPUT112), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n757), .B1(new_n837), .B2(new_n838), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT112), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n842), .B1(new_n837), .B2(new_n838), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n840), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n845), .A2(new_n756), .A3(new_n729), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n832), .A2(new_n833), .A3(new_n846), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(new_n262), .ZN(G39));
  NAND4_X1  g662(.A1(new_n709), .A2(new_n764), .A3(new_n748), .A4(new_n799), .ZN(new_n849));
  XOR2_X1   g663(.A(new_n849), .B(KEYINPUT114), .Z(new_n850));
  NAND3_X1  g664(.A1(new_n845), .A2(KEYINPUT47), .A3(new_n756), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT47), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n852), .B1(new_n844), .B2(new_n189), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n850), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n854), .B(new_n340), .ZN(G42));
  NOR3_X1   g669(.A1(new_n764), .A2(new_n189), .A3(new_n443), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT49), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n755), .A2(new_n757), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n856), .B(new_n825), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  XOR2_X1   g673(.A(new_n859), .B(KEYINPUT115), .Z(new_n860));
  INV_X1    g674(.A(new_n740), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n743), .B1(new_n857), .B2(new_n858), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n429), .A2(new_n193), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT54), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n802), .A2(new_n756), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n725), .A2(new_n715), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n861), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n868), .A2(new_n664), .A3(new_n726), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n749), .A2(new_n796), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n723), .A2(new_n869), .A3(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT52), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n870), .B1(new_n722), .B2(new_n718), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n875), .A2(KEYINPUT52), .A3(new_n869), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(KEYINPUT117), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT53), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n773), .A2(new_n778), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n770), .A2(new_n790), .A3(new_n815), .A4(new_n880), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n684), .A2(new_n685), .A3(new_n714), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n314), .A2(new_n882), .A3(new_n799), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n883), .A2(new_n719), .A3(new_n652), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n794), .A2(new_n813), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n818), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n504), .A2(new_n437), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n659), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n665), .A2(new_n678), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(KEYINPUT116), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT116), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n665), .A2(new_n678), .A3(new_n891), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n890), .B(new_n892), .C1(new_n665), .C2(new_n686), .ZN(new_n893));
  AOI22_X1  g707(.A1(new_n888), .A2(new_n893), .B1(new_n505), .B2(new_n704), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n886), .A2(new_n654), .A3(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n881), .A2(new_n895), .ZN(new_n896));
  AND4_X1   g710(.A1(KEYINPUT52), .A2(new_n723), .A3(new_n869), .A4(new_n871), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT52), .B1(new_n875), .B2(new_n869), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n878), .A2(new_n879), .A3(new_n899), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n877), .B(new_n896), .C1(KEYINPUT117), .C2(KEYINPUT53), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n865), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n886), .A2(KEYINPUT53), .A3(new_n654), .A4(new_n894), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n903), .B1(KEYINPUT118), .B2(new_n881), .ZN(new_n904));
  OR2_X1    g718(.A1(new_n881), .A2(KEYINPUT118), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n877), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(KEYINPUT53), .B1(new_n877), .B2(new_n896), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n906), .A2(new_n907), .A3(KEYINPUT54), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n432), .B1(new_n826), .B2(new_n828), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n776), .A2(new_n799), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n909), .A2(new_n563), .A3(new_n811), .A4(new_n910), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT48), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n861), .A2(new_n563), .A3(new_n433), .A4(new_n910), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n430), .B1(new_n913), .B2(new_n889), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n793), .A2(new_n764), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n909), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n914), .B1(new_n795), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n858), .A2(new_n189), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n851), .A2(new_n853), .A3(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n919), .A2(new_n799), .A3(new_n916), .ZN(new_n920));
  OR3_X1    g734(.A1(new_n913), .A2(new_n665), .A3(new_n678), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n743), .A2(new_n442), .A3(new_n758), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n909), .A2(new_n915), .A3(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT50), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n909), .A2(KEYINPUT50), .A3(new_n915), .A4(new_n922), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n909), .A2(new_n794), .A3(new_n910), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT119), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n909), .A2(KEYINPUT119), .A3(new_n794), .A4(new_n910), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n921), .A2(new_n927), .A3(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT51), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n920), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n934), .B1(new_n920), .B2(new_n933), .ZN(new_n936));
  OAI211_X1 g750(.A(new_n912), .B(new_n917), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n902), .A2(new_n908), .A3(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT120), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n864), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NOR4_X1   g754(.A1(new_n902), .A2(new_n908), .A3(new_n937), .A4(KEYINPUT120), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n863), .B1(new_n940), .B2(new_n941), .ZN(G75));
  INV_X1    g756(.A(KEYINPUT121), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n193), .A2(G952), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n899), .A2(new_n879), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n877), .A2(new_n904), .A3(new_n905), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n191), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(KEYINPUT56), .B1(new_n948), .B2(G210), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n478), .A2(new_n481), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(new_n487), .Z(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT55), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n945), .B1(new_n949), .B2(new_n953), .ZN(new_n954));
  OAI211_X1 g768(.A(G210), .B(G902), .C1(new_n906), .C2(new_n907), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT56), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n957), .A2(new_n952), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n943), .B1(new_n954), .B2(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n944), .B1(new_n957), .B2(new_n952), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n949), .A2(new_n953), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n960), .A2(KEYINPUT121), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n959), .A2(new_n962), .ZN(G51));
  NAND2_X1  g777(.A1(new_n287), .A2(new_n298), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT122), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n946), .A2(new_n947), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(KEYINPUT54), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n946), .A2(new_n865), .A3(new_n947), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n192), .B(KEYINPUT57), .Z(new_n970));
  OAI21_X1  g784(.A(new_n965), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n948), .ZN(new_n972));
  OR3_X1    g786(.A1(new_n972), .A2(new_n834), .A3(new_n836), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n944), .B1(new_n971), .B2(new_n973), .ZN(G54));
  NAND2_X1  g788(.A1(KEYINPUT58), .A2(G475), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n972), .A2(new_n380), .A3(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n975), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n377), .B1(new_n948), .B2(new_n977), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n976), .A2(new_n944), .A3(new_n978), .ZN(G60));
  NAND2_X1  g793(.A1(G478), .A2(G902), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT59), .Z(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n675), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n945), .B1(new_n969), .B2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(new_n675), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n982), .B1(new_n902), .B2(new_n908), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n984), .B1(new_n985), .B2(new_n986), .ZN(G63));
  NAND2_X1  g801(.A1(G217), .A2(G902), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(KEYINPUT60), .ZN(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n966), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(new_n552), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n989), .B1(new_n946), .B2(new_n947), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n694), .A2(new_n695), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n944), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n992), .A2(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT123), .ZN(new_n997));
  INV_X1    g811(.A(new_n994), .ZN(new_n998));
  OAI211_X1 g812(.A(new_n997), .B(new_n945), .C1(new_n991), .C2(new_n998), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n996), .A2(KEYINPUT61), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT61), .ZN(new_n1001));
  OAI211_X1 g815(.A(new_n992), .B(new_n995), .C1(new_n997), .C2(new_n1001), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n1000), .A2(new_n1002), .ZN(G66));
  INV_X1    g817(.A(G224), .ZN(new_n1004));
  OAI21_X1  g818(.A(G953), .B1(new_n435), .B2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n770), .A2(new_n790), .A3(new_n880), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n894), .A2(new_n654), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1005), .B1(new_n1008), .B2(G953), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n950), .B1(G898), .B2(new_n193), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1009), .B(new_n1010), .ZN(G69));
  NOR2_X1   g825(.A1(new_n594), .A2(new_n595), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n586), .A2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n1013), .B(new_n365), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n875), .A2(new_n745), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n1015), .A2(KEYINPUT62), .ZN(new_n1016));
  OR2_X1    g830(.A1(new_n645), .A2(new_n653), .ZN(new_n1017));
  AND4_X1   g831(.A1(new_n1017), .A2(new_n314), .A3(new_n729), .A4(new_n799), .ZN(new_n1018));
  XNOR2_X1  g832(.A(new_n893), .B(KEYINPUT124), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1016), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n847), .A2(new_n854), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1015), .A2(KEYINPUT62), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1014), .B1(new_n1023), .B2(new_n193), .ZN(new_n1024));
  NAND2_X1  g838(.A1(G900), .A2(G953), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1014), .A2(new_n1025), .ZN(new_n1026));
  AND2_X1   g840(.A1(new_n815), .A2(new_n818), .ZN(new_n1027));
  NAND4_X1  g841(.A1(new_n811), .A2(new_n563), .A3(new_n664), .A4(new_n726), .ZN(new_n1028));
  OAI211_X1 g842(.A(new_n1027), .B(new_n875), .C1(new_n846), .C2(new_n1028), .ZN(new_n1029));
  NOR3_X1   g843(.A1(new_n847), .A2(new_n854), .A3(new_n1029), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n1026), .B1(new_n1030), .B2(new_n193), .ZN(new_n1031));
  NOR2_X1   g845(.A1(new_n1024), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n193), .B1(G227), .B2(G900), .ZN(new_n1033));
  XNOR2_X1  g847(.A(new_n1033), .B(KEYINPUT125), .ZN(new_n1034));
  XOR2_X1   g848(.A(new_n1032), .B(new_n1034), .Z(G72));
  XNOR2_X1  g849(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1036));
  NAND2_X1  g850(.A1(G472), .A2(G902), .ZN(new_n1037));
  XNOR2_X1  g851(.A(new_n1036), .B(new_n1037), .ZN(new_n1038));
  INV_X1    g852(.A(new_n1038), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n1039), .B1(new_n1030), .B2(new_n1008), .ZN(new_n1040));
  OR2_X1    g854(.A1(new_n637), .A2(new_n567), .ZN(new_n1041));
  OAI21_X1  g855(.A(new_n945), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g856(.A(KEYINPUT127), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  OAI211_X1 g858(.A(KEYINPUT127), .B(new_n945), .C1(new_n1040), .C2(new_n1041), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g860(.A(new_n1008), .ZN(new_n1047));
  OAI21_X1  g861(.A(new_n1038), .B1(new_n1023), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g862(.A(new_n735), .ZN(new_n1049));
  NAND2_X1  g863(.A1(new_n900), .A2(new_n901), .ZN(new_n1050));
  AND3_X1   g864(.A1(new_n1041), .A2(new_n735), .A3(new_n1038), .ZN(new_n1051));
  AOI22_X1  g865(.A1(new_n1048), .A2(new_n1049), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  AND2_X1   g866(.A1(new_n1046), .A2(new_n1052), .ZN(G57));
endmodule


