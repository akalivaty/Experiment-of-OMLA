//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 0 0 1 1 1 0 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 1 1 0 0 1 1 1 1 1 1 0 1 1 0 0 0 0 0 1 0 0 0 0 0 1 1 1 0 1 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:38 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n718, new_n719, new_n720,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT81), .ZN(new_n188));
  INV_X1    g002(.A(G128), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G119), .ZN(new_n190));
  INV_X1    g004(.A(G119), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G128), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT24), .B(G110), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n189), .A2(KEYINPUT23), .A3(G119), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT78), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT78), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n198), .A2(new_n189), .A3(KEYINPUT23), .A4(G119), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT23), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n190), .A2(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n200), .A2(new_n202), .A3(new_n192), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT80), .B(G110), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n195), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G140), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G125), .ZN(new_n207));
  INV_X1    g021(.A(G125), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G140), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n207), .A2(new_n209), .A3(KEYINPUT16), .ZN(new_n210));
  OR3_X1    g024(.A1(new_n208), .A2(KEYINPUT16), .A3(G140), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(new_n211), .A3(G146), .ZN(new_n212));
  AND2_X1   g026(.A1(new_n207), .A2(new_n209), .ZN(new_n213));
  INV_X1    g027(.A(G146), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AND2_X1   g029(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n205), .A2(new_n216), .ZN(new_n217));
  AND3_X1   g031(.A1(new_n210), .A2(G146), .A3(new_n211), .ZN(new_n218));
  AOI21_X1  g032(.A(G146), .B1(new_n210), .B2(new_n211), .ZN(new_n219));
  OAI22_X1  g033(.A1(new_n218), .A2(new_n219), .B1(new_n193), .B2(new_n194), .ZN(new_n220));
  INV_X1    g034(.A(G110), .ZN(new_n221));
  AOI22_X1  g035(.A1(new_n197), .A2(new_n199), .B1(new_n191), .B2(G128), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n221), .B1(new_n222), .B2(new_n202), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT79), .ZN(new_n224));
  NOR3_X1   g038(.A1(new_n220), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n193), .A2(new_n194), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n210), .A2(new_n211), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(new_n214), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n226), .B1(new_n228), .B2(new_n212), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n203), .A2(G110), .ZN(new_n230));
  AOI21_X1  g044(.A(KEYINPUT79), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n188), .B(new_n217), .C1(new_n225), .C2(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT22), .B(G137), .ZN(new_n233));
  INV_X1    g047(.A(G953), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(G221), .A3(G234), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n233), .B(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n232), .A2(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n224), .B1(new_n220), .B2(new_n223), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n229), .A2(KEYINPUT79), .A3(new_n230), .ZN(new_n240));
  AOI22_X1  g054(.A1(new_n239), .A2(new_n240), .B1(new_n205), .B2(new_n216), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n241), .A2(new_n188), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n238), .A2(new_n242), .ZN(new_n243));
  NOR3_X1   g057(.A1(new_n241), .A2(new_n188), .A3(new_n237), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n187), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT25), .ZN(new_n246));
  NAND2_X1  g060(.A1(G217), .A2(G902), .ZN(new_n247));
  INV_X1    g061(.A(G217), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n247), .B1(new_n248), .B2(G234), .ZN(new_n249));
  XNOR2_X1  g063(.A(new_n249), .B(KEYINPUT77), .ZN(new_n250));
  INV_X1    g064(.A(new_n244), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n217), .B1(new_n225), .B2(new_n231), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT81), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n253), .A2(new_n232), .A3(new_n237), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT25), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n255), .A2(new_n256), .A3(new_n187), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n246), .A2(new_n250), .A3(new_n257), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n250), .A2(G902), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  AND3_X1   g074(.A1(new_n258), .A2(KEYINPUT82), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(KEYINPUT82), .B1(new_n258), .B2(new_n260), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT11), .ZN(new_n265));
  INV_X1    g079(.A(G134), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n265), .B1(new_n266), .B2(G137), .ZN(new_n267));
  INV_X1    g081(.A(G137), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n268), .A2(KEYINPUT11), .A3(G134), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n266), .A2(G137), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n267), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G131), .ZN(new_n272));
  INV_X1    g086(.A(G131), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n267), .A2(new_n269), .A3(new_n273), .A4(new_n270), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT65), .ZN(new_n276));
  INV_X1    g090(.A(G143), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n276), .B1(new_n277), .B2(G146), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n214), .A2(KEYINPUT65), .A3(G143), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n277), .A2(G146), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  AND2_X1   g095(.A1(KEYINPUT0), .A2(G128), .ZN(new_n282));
  NOR2_X1   g096(.A1(KEYINPUT0), .A2(G128), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n214), .A2(G143), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n286), .A2(new_n280), .A3(new_n282), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT66), .ZN(new_n288));
  XNOR2_X1  g102(.A(G143), .B(G146), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT66), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n289), .A2(new_n290), .A3(new_n282), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n285), .A2(new_n288), .A3(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(KEYINPUT67), .B1(new_n275), .B2(new_n292), .ZN(new_n293));
  AND2_X1   g107(.A1(new_n288), .A2(new_n291), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n272), .A2(new_n274), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT67), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n294), .A2(new_n295), .A3(new_n296), .A4(new_n285), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n293), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT1), .ZN(new_n299));
  AND3_X1   g113(.A1(new_n286), .A2(new_n280), .A3(G128), .ZN(new_n300));
  OAI21_X1  g114(.A(KEYINPUT1), .B1(new_n277), .B2(G146), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G128), .ZN(new_n302));
  AOI22_X1  g116(.A1(new_n299), .A2(new_n300), .B1(new_n281), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT68), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n266), .A2(G137), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n268), .A2(G134), .ZN(new_n306));
  OAI21_X1  g120(.A(G131), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n274), .A2(new_n307), .ZN(new_n308));
  NOR3_X1   g122(.A1(new_n303), .A2(new_n304), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n281), .A2(new_n302), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n289), .A2(new_n299), .A3(G128), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AND2_X1   g126(.A1(new_n274), .A2(new_n307), .ZN(new_n313));
  AOI21_X1  g127(.A(KEYINPUT68), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n309), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n264), .B1(new_n298), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G113), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT2), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT2), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G113), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G116), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(KEYINPUT69), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT69), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G116), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n191), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n191), .A2(G116), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n322), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT70), .ZN(new_n331));
  XNOR2_X1  g145(.A(KEYINPUT69), .B(G116), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n321), .B(new_n328), .C1(new_n332), .C2(new_n191), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n330), .A2(new_n331), .A3(new_n333), .ZN(new_n334));
  OAI211_X1 g148(.A(KEYINPUT70), .B(new_n322), .C1(new_n327), .C2(new_n329), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n294), .A2(new_n295), .A3(new_n285), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n312), .A2(new_n313), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n338), .A2(KEYINPUT30), .A3(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n316), .A2(new_n337), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT31), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n336), .A2(new_n338), .A3(new_n339), .ZN(new_n343));
  NOR2_X1   g157(.A1(G237), .A2(G953), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(G210), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n345), .B(G101), .ZN(new_n346));
  XNOR2_X1  g160(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n346), .B(new_n347), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n341), .A2(new_n342), .A3(new_n343), .A4(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT71), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n343), .ZN(new_n352));
  INV_X1    g166(.A(new_n340), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n293), .B(new_n297), .C1(new_n314), .C2(new_n309), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n353), .B1(new_n354), .B2(new_n264), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n352), .B1(new_n355), .B2(new_n337), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n356), .A2(KEYINPUT71), .A3(new_n342), .A4(new_n348), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n351), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT28), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n343), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT74), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n354), .A2(new_n361), .A3(new_n337), .ZN(new_n362));
  XNOR2_X1  g176(.A(KEYINPUT73), .B(KEYINPUT28), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n343), .A2(KEYINPUT74), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n365), .B1(new_n337), .B2(new_n354), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n360), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  XOR2_X1   g181(.A(new_n348), .B(KEYINPUT72), .Z(new_n368));
  NAND3_X1  g182(.A1(new_n341), .A2(new_n343), .A3(new_n348), .ZN(new_n369));
  AOI22_X1  g183(.A1(new_n367), .A2(new_n368), .B1(new_n369), .B2(KEYINPUT31), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n358), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G472), .ZN(new_n372));
  AND4_X1   g186(.A1(KEYINPUT32), .A2(new_n371), .A3(new_n372), .A4(new_n187), .ZN(new_n373));
  AOI21_X1  g187(.A(G902), .B1(new_n358), .B2(new_n370), .ZN(new_n374));
  AOI21_X1  g188(.A(KEYINPUT32), .B1(new_n374), .B2(new_n372), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n368), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n360), .B(new_n377), .C1(new_n364), .C2(new_n366), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(KEYINPUT75), .ZN(new_n379));
  AND2_X1   g193(.A1(new_n354), .A2(new_n337), .ZN(new_n380));
  OAI211_X1 g194(.A(new_n363), .B(new_n362), .C1(new_n380), .C2(new_n365), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT75), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n381), .A2(new_n382), .A3(new_n360), .A4(new_n377), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n341), .A2(new_n343), .ZN(new_n384));
  INV_X1    g198(.A(new_n348), .ZN(new_n385));
  AOI21_X1  g199(.A(KEYINPUT29), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n379), .A2(new_n383), .A3(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT76), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n360), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n336), .B1(new_n338), .B2(new_n339), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n352), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n390), .B1(new_n393), .B2(KEYINPUT28), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n394), .A2(KEYINPUT29), .ZN(new_n395));
  AOI21_X1  g209(.A(G902), .B1(new_n395), .B2(new_n348), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n379), .A2(new_n383), .A3(new_n386), .A4(KEYINPUT76), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n389), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G472), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n263), .B1(new_n376), .B2(new_n399), .ZN(new_n400));
  AND2_X1   g214(.A1(new_n234), .A2(G952), .ZN(new_n401));
  NAND2_X1  g215(.A1(G234), .A2(G237), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  XOR2_X1   g218(.A(KEYINPUT21), .B(G898), .Z(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n402), .A2(G902), .A3(G953), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n404), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(G214), .B1(G237), .B2(G902), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n411), .B(KEYINPUT84), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n288), .A2(new_n291), .ZN(new_n414));
  XNOR2_X1  g228(.A(KEYINPUT0), .B(G128), .ZN(new_n415));
  AOI21_X1  g229(.A(KEYINPUT65), .B1(new_n214), .B2(G143), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n214), .A2(G143), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n415), .B1(new_n418), .B2(new_n279), .ZN(new_n419));
  OAI21_X1  g233(.A(G125), .B1(new_n414), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n310), .A2(new_n208), .A3(new_n311), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n234), .A2(G224), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT7), .ZN(new_n425));
  NOR3_X1   g239(.A1(new_n421), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(G104), .ZN(new_n427));
  OAI21_X1  g241(.A(KEYINPUT3), .B1(new_n427), .B2(G107), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT3), .ZN(new_n429));
  INV_X1    g243(.A(G107), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n429), .A2(new_n430), .A3(G104), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n427), .A2(G107), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n428), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(G101), .ZN(new_n434));
  INV_X1    g248(.A(G101), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n428), .A2(new_n431), .A3(new_n435), .A4(new_n432), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n434), .A2(KEYINPUT4), .A3(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT4), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n433), .A2(new_n438), .A3(G101), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n336), .A2(new_n440), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n427), .A2(G107), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n430), .A2(G104), .ZN(new_n443));
  OAI21_X1  g257(.A(G101), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  AND2_X1   g258(.A1(new_n436), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n333), .ZN(new_n446));
  OAI211_X1 g260(.A(KEYINPUT5), .B(new_n328), .C1(new_n332), .C2(new_n191), .ZN(new_n447));
  OR2_X1    g261(.A1(new_n328), .A2(KEYINPUT5), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n447), .A2(G113), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(KEYINPUT85), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT85), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n447), .A2(new_n451), .A3(G113), .A4(new_n448), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n446), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n441), .A2(new_n453), .ZN(new_n454));
  XOR2_X1   g268(.A(G110), .B(G122), .Z(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n426), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n422), .A2(KEYINPUT88), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT88), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n310), .A2(new_n459), .A3(new_n208), .A4(new_n311), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n458), .A2(new_n420), .A3(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT89), .ZN(new_n462));
  AND3_X1   g276(.A1(new_n461), .A2(new_n462), .A3(new_n425), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n462), .B1(new_n461), .B2(new_n425), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  XOR2_X1   g279(.A(new_n455), .B(KEYINPUT8), .Z(new_n466));
  NAND2_X1  g280(.A1(new_n450), .A2(new_n452), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n445), .B1(new_n467), .B2(new_n333), .ZN(new_n468));
  INV_X1    g282(.A(new_n449), .ZN(new_n469));
  OAI21_X1  g283(.A(KEYINPUT87), .B1(new_n469), .B2(new_n446), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT87), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n449), .A2(new_n471), .A3(new_n333), .A4(new_n445), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n466), .B1(new_n468), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n457), .A2(new_n465), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n187), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT90), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT6), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n479), .B1(new_n454), .B2(new_n456), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n480), .B1(new_n456), .B2(new_n454), .ZN(new_n481));
  INV_X1    g295(.A(new_n454), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n482), .A2(new_n479), .A3(new_n455), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n421), .A2(new_n423), .ZN(new_n484));
  XOR2_X1   g298(.A(new_n424), .B(KEYINPUT86), .Z(new_n485));
  XOR2_X1   g299(.A(new_n484), .B(new_n485), .Z(new_n486));
  NAND3_X1  g300(.A1(new_n481), .A2(new_n483), .A3(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n475), .A2(KEYINPUT90), .A3(new_n187), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n478), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(G210), .B1(G237), .B2(G902), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n478), .A2(new_n490), .A3(new_n487), .A4(new_n488), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n413), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(G128), .B(G143), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n495), .B(new_n266), .ZN(new_n496));
  OR2_X1    g310(.A1(KEYINPUT93), .A2(G122), .ZN(new_n497));
  NAND2_X1  g311(.A1(KEYINPUT93), .A2(G122), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n323), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(G122), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n500), .B1(new_n324), .B2(new_n326), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n430), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT96), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT14), .ZN(new_n505));
  OAI21_X1  g319(.A(KEYINPUT95), .B1(new_n501), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT95), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n507), .B(KEYINPUT14), .C1(new_n332), .C2(new_n500), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n499), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n504), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AOI211_X1 g325(.A(KEYINPUT96), .B(new_n499), .C1(new_n506), .C2(new_n508), .ZN(new_n512));
  NOR3_X1   g326(.A1(new_n332), .A2(KEYINPUT14), .A3(new_n500), .ZN(new_n513));
  NOR3_X1   g327(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n496), .B(new_n503), .C1(new_n514), .C2(new_n430), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n502), .B(G107), .ZN(new_n516));
  NOR3_X1   g330(.A1(new_n189), .A2(KEYINPUT13), .A3(G143), .ZN(new_n517));
  AOI211_X1 g331(.A(new_n266), .B(new_n517), .C1(KEYINPUT13), .C2(new_n495), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n495), .A2(new_n266), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n519), .B(KEYINPUT94), .ZN(new_n520));
  OR3_X1    g334(.A1(new_n516), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n515), .A2(new_n521), .ZN(new_n522));
  XOR2_X1   g336(.A(KEYINPUT9), .B(G234), .Z(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NOR3_X1   g338(.A1(new_n524), .A2(new_n248), .A3(G953), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n515), .A2(new_n521), .A3(new_n525), .ZN(new_n528));
  AOI21_X1  g342(.A(G902), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(G478), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n529), .B1(KEYINPUT15), .B2(new_n530), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n515), .A2(new_n521), .A3(new_n525), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n525), .B1(new_n515), .B2(new_n521), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n187), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT15), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(new_n535), .A3(G478), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n531), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n218), .A2(new_n219), .ZN(new_n538));
  AND3_X1   g352(.A1(new_n344), .A2(G143), .A3(G214), .ZN(new_n539));
  AOI21_X1  g353(.A(G143), .B1(new_n344), .B2(G214), .ZN(new_n540));
  OAI211_X1 g354(.A(KEYINPUT17), .B(G131), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n539), .A2(new_n540), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(new_n273), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n538), .B(new_n541), .C1(new_n543), .C2(KEYINPUT17), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT91), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n546), .A2(KEYINPUT18), .A3(G131), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n213), .B(new_n214), .ZN(new_n548));
  NAND2_X1  g362(.A1(KEYINPUT18), .A2(G131), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n549), .B1(new_n542), .B2(new_n545), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n547), .B(new_n548), .C1(new_n550), .C2(new_n546), .ZN(new_n551));
  XNOR2_X1  g365(.A(G113), .B(G122), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n552), .B(new_n427), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n544), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  XOR2_X1   g368(.A(new_n213), .B(KEYINPUT19), .Z(new_n555));
  OAI211_X1 g369(.A(new_n543), .B(new_n212), .C1(G146), .C2(new_n555), .ZN(new_n556));
  AND2_X1   g370(.A1(new_n556), .A2(new_n551), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n554), .B1(new_n557), .B2(new_n553), .ZN(new_n558));
  INV_X1    g372(.A(G475), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n558), .A2(new_n559), .A3(new_n187), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT20), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT20), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n558), .A2(new_n562), .A3(new_n559), .A4(new_n187), .ZN(new_n563));
  INV_X1    g377(.A(new_n554), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n553), .B1(new_n544), .B2(new_n551), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n187), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(KEYINPUT92), .B(G475), .ZN(new_n567));
  AOI22_X1  g381(.A1(new_n561), .A2(new_n563), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n537), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(G469), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT10), .ZN(new_n572));
  INV_X1    g386(.A(new_n311), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n289), .B1(G128), .B2(new_n301), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n436), .A2(new_n444), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n572), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n437), .A2(new_n294), .A3(new_n285), .A4(new_n439), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n312), .A2(new_n445), .A3(KEYINPUT10), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n577), .A2(new_n578), .A3(new_n275), .A4(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(G110), .B(G140), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n234), .A2(G227), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n581), .B(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(KEYINPUT83), .B1(new_n312), .B2(new_n445), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n445), .B1(new_n573), .B2(new_n574), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT83), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n303), .A2(new_n587), .A3(new_n576), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n585), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n295), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT12), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n589), .A2(KEYINPUT12), .A3(new_n295), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n584), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n295), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n583), .B1(new_n596), .B2(new_n580), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n571), .B(new_n187), .C1(new_n594), .C2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n596), .A2(new_n580), .A3(new_n583), .ZN(new_n599));
  INV_X1    g413(.A(new_n580), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n600), .B1(new_n592), .B2(new_n593), .ZN(new_n601));
  OAI211_X1 g415(.A(G469), .B(new_n599), .C1(new_n601), .C2(new_n583), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n571), .A2(new_n187), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n598), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  OAI21_X1  g419(.A(G221), .B1(new_n524), .B2(G902), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AND3_X1   g421(.A1(new_n494), .A2(new_n570), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n400), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(G101), .ZN(G3));
  INV_X1    g424(.A(new_n263), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n374), .B(G472), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n611), .A2(new_n607), .A3(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT99), .ZN(new_n615));
  OAI21_X1  g429(.A(KEYINPUT97), .B1(new_n532), .B2(new_n533), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT33), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OAI211_X1 g432(.A(KEYINPUT97), .B(KEYINPUT33), .C1(new_n532), .C2(new_n533), .ZN(new_n619));
  AOI211_X1 g433(.A(new_n530), .B(G902), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n529), .A2(KEYINPUT98), .A3(G478), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT98), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n622), .B1(new_n534), .B2(new_n530), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n569), .B1(new_n620), .B2(new_n624), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n475), .A2(KEYINPUT90), .A3(new_n187), .ZN(new_n626));
  AOI21_X1  g440(.A(KEYINPUT90), .B1(new_n475), .B2(new_n187), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n490), .B1(new_n628), .B2(new_n487), .ZN(new_n629));
  INV_X1    g443(.A(new_n493), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n410), .B(new_n411), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n615), .B1(new_n625), .B2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n411), .ZN(new_n633));
  AOI211_X1 g447(.A(new_n409), .B(new_n633), .C1(new_n492), .C2(new_n493), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n527), .A2(new_n528), .ZN(new_n635));
  AOI21_X1  g449(.A(KEYINPUT33), .B1(new_n635), .B2(KEYINPUT97), .ZN(new_n636));
  INV_X1    g450(.A(new_n619), .ZN(new_n637));
  OAI211_X1 g451(.A(G478), .B(new_n187), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  OAI21_X1  g452(.A(KEYINPUT98), .B1(new_n529), .B2(G478), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n534), .A2(new_n622), .A3(new_n530), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n568), .B1(new_n638), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n634), .A2(KEYINPUT99), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n632), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n614), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT34), .B(G104), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G6));
  AOI21_X1  g461(.A(new_n633), .B1(new_n492), .B2(new_n493), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT100), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n563), .A2(new_n649), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n650), .A2(new_n561), .ZN(new_n651));
  OR2_X1    g465(.A1(new_n563), .A2(new_n649), .ZN(new_n652));
  AOI22_X1  g466(.A1(new_n651), .A2(new_n652), .B1(new_n566), .B2(new_n567), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n648), .A2(new_n653), .A3(new_n410), .A4(new_n537), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(KEYINPUT101), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT101), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n634), .A2(new_n656), .A3(new_n537), .A4(new_n653), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n614), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT35), .B(G107), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G9));
  NOR2_X1   g475(.A1(new_n237), .A2(KEYINPUT36), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n252), .B(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n259), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n258), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n608), .A2(new_n612), .A3(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT37), .B(G110), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT102), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n666), .B(new_n668), .ZN(G12));
  NAND3_X1  g483(.A1(new_n371), .A2(new_n372), .A3(new_n187), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT32), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n374), .A2(KEYINPUT32), .A3(new_n372), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n399), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n492), .A2(new_n493), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n675), .A2(new_n411), .A3(new_n665), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n403), .B(KEYINPUT104), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  XOR2_X1   g493(.A(KEYINPUT103), .B(G900), .Z(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n408), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  AND3_X1   g496(.A1(new_n653), .A2(new_n537), .A3(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n674), .A2(new_n677), .A3(new_n607), .A4(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G128), .ZN(G30));
  XNOR2_X1  g499(.A(new_n675), .B(KEYINPUT38), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT105), .B(KEYINPUT39), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n682), .B(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n607), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(KEYINPUT40), .ZN(new_n690));
  INV_X1    g504(.A(new_n369), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n691), .B1(new_n368), .B2(new_n393), .ZN(new_n692));
  OAI21_X1  g506(.A(G472), .B1(new_n692), .B2(G902), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n672), .A2(new_n673), .A3(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n686), .A2(new_n690), .A3(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n665), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n696), .B1(new_n689), .B2(KEYINPUT40), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n568), .B1(new_n531), .B2(new_n536), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NOR4_X1   g513(.A1(new_n695), .A2(new_n633), .A3(new_n697), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(new_n277), .ZN(G45));
  INV_X1    g515(.A(new_n682), .ZN(new_n702));
  AOI211_X1 g516(.A(new_n568), .B(new_n702), .C1(new_n638), .C2(new_n641), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n674), .A2(new_n677), .A3(new_n703), .A4(new_n607), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G146), .ZN(G48));
  OR2_X1    g519(.A1(new_n594), .A2(new_n597), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n571), .B1(new_n706), .B2(new_n187), .ZN(new_n707));
  INV_X1    g521(.A(new_n598), .ZN(new_n708));
  OR2_X1    g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(new_n606), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AND3_X1   g525(.A1(new_n674), .A2(new_n611), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n644), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT41), .B(G113), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G15));
  NAND2_X1  g529(.A1(new_n712), .A2(new_n658), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G116), .ZN(G18));
  AOI21_X1  g531(.A(new_n676), .B1(new_n376), .B2(new_n399), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n537), .A2(new_n569), .A3(new_n409), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n718), .A2(new_n711), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G119), .ZN(G21));
  NAND2_X1  g535(.A1(new_n371), .A2(new_n187), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(G472), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n369), .A2(KEYINPUT31), .ZN(new_n724));
  OAI211_X1 g538(.A(new_n358), .B(new_n724), .C1(new_n377), .C2(new_n394), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n725), .A2(new_n372), .A3(new_n187), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n258), .A2(new_n260), .ZN(new_n728));
  NOR4_X1   g542(.A1(new_n727), .A2(new_n728), .A3(new_n710), .A4(new_n709), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n631), .A2(new_n699), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G122), .ZN(G24));
  NOR2_X1   g546(.A1(new_n727), .A2(new_n696), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n733), .A2(new_n703), .A3(new_n648), .A4(new_n711), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G125), .ZN(G27));
  INV_X1    g549(.A(KEYINPUT42), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n569), .B(new_n682), .C1(new_n620), .C2(new_n624), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n629), .A2(new_n630), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT107), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n605), .A2(KEYINPUT106), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT106), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n598), .A2(new_n602), .A3(new_n741), .A4(new_n604), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n740), .A2(new_n606), .A3(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n738), .A2(new_n739), .A3(new_n411), .A4(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n492), .A2(new_n493), .A3(new_n411), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n740), .A2(new_n606), .A3(new_n742), .ZN(new_n746));
  OAI21_X1  g560(.A(KEYINPUT107), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n737), .B1(new_n744), .B2(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n728), .B1(new_n376), .B2(new_n399), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n736), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n744), .A2(new_n747), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n737), .A2(KEYINPUT42), .ZN(new_n752));
  AND3_X1   g566(.A1(new_n400), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G131), .ZN(G33));
  NAND3_X1  g569(.A1(new_n400), .A2(new_n751), .A3(new_n683), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT108), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n400), .A2(new_n751), .A3(KEYINPUT108), .A4(new_n683), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G134), .ZN(G36));
  NOR2_X1   g575(.A1(new_n612), .A2(new_n696), .ZN(new_n762));
  XOR2_X1   g576(.A(new_n762), .B(KEYINPUT110), .Z(new_n763));
  NAND2_X1  g577(.A1(new_n638), .A2(new_n641), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(new_n568), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(KEYINPUT43), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT43), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n764), .A2(new_n767), .A3(new_n568), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n763), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT44), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n745), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n599), .B1(new_n601), .B2(new_n583), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(KEYINPUT45), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(G469), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(KEYINPUT109), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT109), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n775), .A2(new_n778), .A3(G469), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n603), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n708), .B1(new_n780), .B2(KEYINPUT46), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT46), .ZN(new_n782));
  INV_X1    g596(.A(new_n779), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n778), .B1(new_n775), .B2(G469), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n782), .B1(new_n785), .B2(new_n603), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n710), .B1(new_n781), .B2(new_n786), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n787), .A2(new_n688), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n763), .A2(KEYINPUT44), .A3(new_n769), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n772), .A2(new_n773), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G137), .ZN(G39));
  NAND2_X1  g605(.A1(new_n777), .A2(new_n779), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n792), .A2(KEYINPUT46), .A3(new_n604), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(new_n598), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n780), .A2(KEYINPUT46), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n606), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(KEYINPUT47), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT47), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n787), .A2(new_n798), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n674), .A2(new_n611), .A3(new_n745), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n797), .A2(new_n799), .A3(new_n703), .A4(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G140), .ZN(G42));
  NOR2_X1   g616(.A1(new_n709), .A2(KEYINPUT49), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n686), .A2(new_n765), .A3(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n694), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n709), .A2(KEYINPUT49), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n258), .A2(new_n260), .A3(new_n412), .A4(new_n606), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(KEYINPUT111), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n804), .A2(new_n805), .A3(new_n806), .A4(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT116), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n709), .A2(new_n606), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n811), .B1(new_n797), .B2(new_n799), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n766), .A2(new_n678), .A3(new_n768), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n727), .A2(new_n728), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n813), .A2(new_n814), .A3(new_n773), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n810), .B1(new_n812), .B2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n811), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n787), .A2(new_n798), .ZN(new_n818));
  AOI211_X1 g632(.A(KEYINPUT47), .B(new_n710), .C1(new_n781), .C2(new_n786), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n817), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n815), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n820), .A2(KEYINPUT116), .A3(new_n821), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n745), .A2(new_n710), .A3(new_n709), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n766), .A2(new_n678), .A3(new_n768), .A4(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n733), .ZN(new_n825));
  OR3_X1    g639(.A1(new_n824), .A2(KEYINPUT117), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(KEYINPUT117), .B1(new_n824), .B2(new_n825), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n686), .A2(new_n411), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n813), .A2(new_n729), .A3(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT50), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n813), .A2(KEYINPUT50), .A3(new_n729), .A4(new_n829), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n805), .A2(new_n611), .A3(new_n404), .A4(new_n823), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n764), .A2(new_n569), .ZN(new_n836));
  AOI22_X1  g650(.A1(new_n832), .A2(new_n833), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n816), .A2(new_n822), .A3(new_n828), .A4(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT118), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT51), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n812), .A2(KEYINPUT119), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT119), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n820), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n842), .A2(new_n844), .A3(new_n821), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n832), .A2(new_n833), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n835), .A2(new_n836), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n846), .A2(new_n828), .A3(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n845), .A2(KEYINPUT51), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(new_n401), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n839), .B1(new_n838), .B2(new_n840), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n841), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n625), .A2(new_n631), .A3(new_n615), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT99), .B1(new_n634), .B2(new_n642), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n674), .A2(new_n611), .A3(new_n711), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n720), .B(new_n731), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n856), .B1(new_n657), .B2(new_n655), .ZN(new_n858));
  OAI21_X1  g672(.A(KEYINPUT112), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AOI22_X1  g673(.A1(new_n712), .A2(new_n644), .B1(new_n730), .B2(new_n729), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT112), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n860), .A2(new_n861), .A3(new_n716), .A4(new_n720), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n537), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n653), .A2(new_n682), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n674), .A2(new_n864), .A3(new_n607), .A4(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n866), .A2(new_n745), .ZN(new_n867));
  AOI211_X1 g681(.A(new_n727), .B(new_n737), .C1(new_n744), .C2(new_n747), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n665), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n869), .A2(new_n760), .A3(new_n754), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT52), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT114), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n694), .A2(new_n743), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n648), .A2(new_n696), .A3(new_n682), .A4(new_n698), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n675), .A2(new_n411), .A3(new_n698), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n696), .A2(new_n682), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n878), .A2(KEYINPUT114), .A3(new_n694), .A4(new_n743), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n734), .A2(new_n684), .A3(new_n704), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n871), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n875), .A2(new_n879), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n718), .B(new_n607), .C1(new_n683), .C2(new_n703), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n883), .A2(KEYINPUT52), .A3(new_n734), .A4(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n642), .A2(new_n494), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(KEYINPUT113), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n864), .A2(new_n569), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(new_n494), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT113), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n642), .A2(new_n891), .A3(new_n494), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n888), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n609), .B(new_n666), .C1(new_n893), .C2(new_n613), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n863), .A2(new_n870), .A3(new_n886), .A4(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT53), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT115), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n885), .A2(new_n899), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n734), .A2(new_n684), .A3(new_n704), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n901), .A2(KEYINPUT115), .A3(KEYINPUT52), .A4(new_n883), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n900), .A2(new_n882), .A3(new_n902), .ZN(new_n903));
  NOR4_X1   g717(.A1(new_n894), .A2(new_n857), .A3(new_n897), .A4(new_n858), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n903), .A2(new_n904), .A3(new_n870), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n898), .A2(new_n905), .ZN(new_n906));
  OR2_X1    g720(.A1(new_n906), .A2(KEYINPUT54), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n813), .A2(new_n648), .A3(new_n729), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n896), .A2(KEYINPUT53), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n894), .B1(new_n859), .B2(new_n862), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n910), .A2(new_n903), .A3(new_n897), .A4(new_n870), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(KEYINPUT54), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n852), .A2(new_n907), .A3(new_n908), .A4(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n834), .A2(new_n625), .ZN(new_n915));
  INV_X1    g729(.A(new_n749), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n824), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT48), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n914), .A2(new_n915), .A3(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(G952), .A2(G953), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n809), .B1(new_n919), .B2(new_n920), .ZN(G75));
  NOR2_X1   g735(.A1(new_n234), .A2(G952), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n903), .A2(new_n904), .ZN(new_n924));
  AOI22_X1  g738(.A1(new_n924), .A2(new_n870), .B1(new_n896), .B2(new_n897), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n925), .A2(new_n187), .ZN(new_n926));
  AOI21_X1  g740(.A(KEYINPUT56), .B1(new_n926), .B2(G210), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n481), .A2(new_n483), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(new_n486), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT55), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n923), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT120), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n932), .B1(new_n925), .B2(new_n187), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n906), .A2(KEYINPUT120), .A3(G902), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n491), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT56), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n930), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n931), .B1(new_n936), .B2(new_n938), .ZN(G51));
  AOI21_X1  g753(.A(KEYINPUT121), .B1(new_n935), .B2(new_n785), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT121), .ZN(new_n941));
  AOI211_X1 g755(.A(new_n941), .B(new_n792), .C1(new_n933), .C2(new_n934), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n906), .B(KEYINPUT54), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n604), .A2(KEYINPUT57), .ZN(new_n945));
  OR2_X1    g759(.A1(new_n604), .A2(KEYINPUT57), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n706), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n922), .B1(new_n943), .B2(new_n948), .ZN(G54));
  NAND2_X1  g763(.A1(KEYINPUT58), .A2(G475), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(KEYINPUT122), .Z(new_n951));
  AND3_X1   g765(.A1(new_n935), .A2(new_n558), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n558), .B1(new_n935), .B2(new_n951), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n952), .A2(new_n953), .A3(new_n922), .ZN(G60));
  NAND2_X1  g768(.A1(new_n618), .A2(new_n619), .ZN(new_n955));
  NAND2_X1  g769(.A1(G478), .A2(G902), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT59), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n944), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n907), .A2(new_n913), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n955), .B1(new_n959), .B2(new_n957), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n958), .A2(new_n960), .A3(new_n922), .ZN(G63));
  XOR2_X1   g775(.A(new_n247), .B(KEYINPUT60), .Z(new_n962));
  NAND3_X1  g776(.A1(new_n906), .A2(new_n663), .A3(new_n962), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n906), .A2(new_n962), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n923), .B(new_n963), .C1(new_n964), .C2(new_n255), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT61), .Z(G66));
  INV_X1    g780(.A(G224), .ZN(new_n967));
  OAI21_X1  g781(.A(G953), .B1(new_n406), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n968), .B1(new_n910), .B2(G953), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n928), .B1(G898), .B2(new_n234), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(G69));
  NAND3_X1  g785(.A1(new_n772), .A2(new_n773), .A3(new_n789), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n972), .B1(new_n916), .B2(new_n876), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n881), .B1(new_n973), .B2(new_n788), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n801), .A2(new_n754), .A3(new_n760), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n974), .A2(new_n234), .A3(new_n975), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n355), .B(new_n555), .ZN(new_n977));
  XOR2_X1   g791(.A(KEYINPUT123), .B(KEYINPUT124), .Z(new_n978));
  XNOR2_X1  g792(.A(new_n977), .B(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(G900), .A2(G953), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n976), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT126), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n700), .A2(new_n881), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT62), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n400), .B1(new_n642), .B2(new_n889), .ZN(new_n985));
  OR3_X1    g799(.A1(new_n985), .A2(new_n689), .A3(new_n745), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n984), .A2(new_n790), .A3(new_n801), .A4(new_n986), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n987), .A2(new_n234), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n979), .B(KEYINPUT125), .Z(new_n989));
  OAI211_X1 g803(.A(new_n981), .B(new_n982), .C1(new_n988), .C2(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n234), .B1(G227), .B2(G900), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n990), .B(new_n991), .ZN(G72));
  NAND2_X1  g806(.A1(G472), .A2(G902), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(KEYINPUT63), .Z(new_n994));
  INV_X1    g808(.A(new_n910), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n994), .B1(new_n987), .B2(new_n995), .ZN(new_n996));
  OR2_X1    g810(.A1(new_n996), .A2(KEYINPUT127), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(KEYINPUT127), .ZN(new_n998));
  NAND4_X1  g812(.A1(new_n997), .A2(new_n384), .A3(new_n348), .A4(new_n998), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n974), .A2(new_n910), .A3(new_n975), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n348), .B1(new_n1000), .B2(new_n994), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n922), .B1(new_n1001), .B2(new_n356), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n356), .A2(new_n348), .ZN(new_n1003));
  OAI211_X1 g817(.A(new_n912), .B(new_n994), .C1(new_n691), .C2(new_n1003), .ZN(new_n1004));
  AND3_X1   g818(.A1(new_n999), .A2(new_n1002), .A3(new_n1004), .ZN(G57));
endmodule


