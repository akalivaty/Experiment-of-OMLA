

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763;

  XNOR2_X1 U382 ( .A(n453), .B(n452), .ZN(n491) );
  BUF_X1 U383 ( .A(G953), .Z(n749) );
  INV_X1 U384 ( .A(G953), .ZN(n377) );
  XNOR2_X2 U385 ( .A(n536), .B(n535), .ZN(n543) );
  XNOR2_X2 U386 ( .A(G119), .B(G116), .ZN(n410) );
  XNOR2_X1 U387 ( .A(n575), .B(KEYINPUT40), .ZN(n588) );
  INV_X1 U388 ( .A(n604), .ZN(n373) );
  XNOR2_X1 U389 ( .A(n363), .B(KEYINPUT89), .ZN(n362) );
  INV_X1 U390 ( .A(n749), .ZN(n368) );
  XNOR2_X1 U391 ( .A(G146), .B(G125), .ZN(n435) );
  INV_X1 U392 ( .A(G953), .ZN(n383) );
  NAND2_X1 U393 ( .A1(n369), .A2(n368), .ZN(n367) );
  XNOR2_X1 U394 ( .A(n370), .B(KEYINPUT121), .ZN(n369) );
  NOR2_X1 U395 ( .A1(n655), .A2(n618), .ZN(n617) );
  NAND2_X1 U396 ( .A1(n373), .A2(n372), .ZN(n386) );
  XNOR2_X1 U397 ( .A(n577), .B(n576), .ZN(n698) );
  AND2_X1 U398 ( .A1(n372), .A2(n391), .ZN(n371) );
  INV_X1 U399 ( .A(n680), .ZN(n372) );
  OR2_X1 U400 ( .A1(n666), .A2(n667), .ZN(n662) );
  XNOR2_X1 U401 ( .A(n457), .B(n456), .ZN(n709) );
  XNOR2_X1 U402 ( .A(n495), .B(n494), .ZN(n634) );
  XNOR2_X1 U403 ( .A(n364), .B(KEYINPUT25), .ZN(n500) );
  NAND2_X1 U404 ( .A1(n497), .A2(G217), .ZN(n364) );
  XNOR2_X1 U405 ( .A(n362), .B(n435), .ZN(n361) );
  XOR2_X1 U406 ( .A(n418), .B(KEYINPUT90), .Z(n378) );
  XNOR2_X1 U407 ( .A(n643), .B(G146), .ZN(n485) );
  XNOR2_X1 U408 ( .A(n471), .B(n470), .ZN(n643) );
  XNOR2_X1 U409 ( .A(n459), .B(n365), .ZN(n497) );
  NAND2_X1 U410 ( .A1(n383), .A2(G224), .ZN(n363) );
  XNOR2_X1 U411 ( .A(G902), .B(KEYINPUT15), .ZN(n618) );
  XNOR2_X1 U412 ( .A(KEYINPUT20), .B(KEYINPUT92), .ZN(n365) );
  XNOR2_X2 U413 ( .A(G143), .B(G128), .ZN(n450) );
  XNOR2_X1 U414 ( .A(KEYINPUT73), .B(KEYINPUT22), .ZN(n466) );
  XNOR2_X1 U415 ( .A(n361), .B(n360), .ZN(n409) );
  NAND2_X1 U416 ( .A1(n359), .A2(n427), .ZN(n428) );
  AND2_X1 U417 ( .A1(n359), .A2(n599), .ZN(n738) );
  XNOR2_X2 U418 ( .A(n590), .B(KEYINPUT19), .ZN(n359) );
  XNOR2_X1 U419 ( .A(n382), .B(n405), .ZN(n360) );
  XNOR2_X1 U420 ( .A(n367), .B(n366), .ZN(G75) );
  INV_X1 U421 ( .A(KEYINPUT53), .ZN(n366) );
  NAND2_X1 U422 ( .A1(n701), .A2(n404), .ZN(n370) );
  NAND2_X1 U423 ( .A1(n373), .A2(n371), .ZN(n388) );
  XNOR2_X1 U424 ( .A(n588), .B(G131), .ZN(G33) );
  BUF_X1 U425 ( .A(n641), .Z(n374) );
  BUF_X1 U426 ( .A(n506), .Z(n375) );
  BUF_X1 U427 ( .A(n655), .Z(n376) );
  NAND2_X2 U428 ( .A1(n402), .A2(n401), .ZN(n590) );
  OR2_X1 U429 ( .A1(n655), .A2(n623), .ZN(n658) );
  XNOR2_X2 U430 ( .A(n450), .B(n449), .ZN(n471) );
  OR2_X1 U431 ( .A1(n558), .A2(n557), .ZN(n560) );
  XNOR2_X1 U432 ( .A(n601), .B(n573), .ZN(n680) );
  XNOR2_X1 U433 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n405) );
  XOR2_X1 U434 ( .A(KEYINPUT82), .B(KEYINPUT39), .Z(n391) );
  INV_X1 U435 ( .A(n679), .ZN(n401) );
  XNOR2_X1 U436 ( .A(G113), .B(KEYINPUT70), .ZN(n411) );
  NOR2_X1 U437 ( .A1(G237), .A2(n749), .ZN(n438) );
  XNOR2_X1 U438 ( .A(n544), .B(KEYINPUT45), .ZN(n545) );
  XNOR2_X1 U439 ( .A(KEYINPUT88), .B(G110), .ZN(n406) );
  XNOR2_X1 U440 ( .A(G128), .B(G110), .ZN(n488) );
  XNOR2_X1 U441 ( .A(G140), .B(KEYINPUT10), .ZN(n436) );
  XNOR2_X1 U442 ( .A(G116), .B(G107), .ZN(n447) );
  XNOR2_X1 U443 ( .A(n498), .B(KEYINPUT105), .ZN(n499) );
  AND2_X1 U444 ( .A1(n464), .A2(n463), .ZN(n465) );
  INV_X1 U445 ( .A(KEYINPUT6), .ZN(n390) );
  NAND2_X1 U446 ( .A1(n630), .A2(n749), .ZN(n725) );
  XNOR2_X1 U447 ( .A(n513), .B(KEYINPUT35), .ZN(n641) );
  NAND2_X1 U448 ( .A1(n384), .A2(n558), .ZN(n379) );
  XOR2_X1 U449 ( .A(KEYINPUT66), .B(KEYINPUT0), .Z(n380) );
  XNOR2_X1 U450 ( .A(n381), .B(KEYINPUT78), .ZN(n620) );
  NAND2_X1 U451 ( .A1(n617), .A2(n616), .ZN(n381) );
  XNOR2_X1 U452 ( .A(G143), .B(G128), .ZN(n382) );
  NAND2_X1 U453 ( .A1(n690), .A2(n509), .ZN(n399) );
  XNOR2_X1 U454 ( .A(n467), .B(n466), .ZN(n384) );
  XNOR2_X1 U455 ( .A(n467), .B(n466), .ZN(n504) );
  NAND2_X1 U456 ( .A1(n504), .A2(n394), .ZN(n400) );
  XNOR2_X1 U457 ( .A(n385), .B(KEYINPUT30), .ZN(n568) );
  NOR2_X1 U458 ( .A1(n669), .A2(n679), .ZN(n385) );
  NAND2_X1 U459 ( .A1(n386), .A2(n387), .ZN(n389) );
  NAND2_X1 U460 ( .A1(n388), .A2(n389), .ZN(n574) );
  INV_X1 U461 ( .A(n391), .ZN(n387) );
  XNOR2_X1 U462 ( .A(n669), .B(n390), .ZN(n558) );
  XNOR2_X2 U463 ( .A(n392), .B(n393), .ZN(n669) );
  NOR2_X1 U464 ( .A1(n704), .A2(G902), .ZN(n392) );
  XOR2_X1 U465 ( .A(n478), .B(KEYINPUT72), .Z(n393) );
  XNOR2_X2 U466 ( .A(n581), .B(KEYINPUT1), .ZN(n595) );
  AND2_X1 U467 ( .A1(n558), .A2(n499), .ZN(n394) );
  NAND2_X1 U468 ( .A1(n508), .A2(n465), .ZN(n467) );
  XNOR2_X1 U469 ( .A(n395), .B(n485), .ZN(n704) );
  XNOR2_X1 U470 ( .A(n396), .B(n475), .ZN(n395) );
  XNOR2_X1 U471 ( .A(n477), .B(n476), .ZN(n396) );
  NAND2_X1 U472 ( .A1(n397), .A2(n512), .ZN(n513) );
  XNOR2_X1 U473 ( .A(n399), .B(n398), .ZN(n397) );
  INV_X1 U474 ( .A(KEYINPUT34), .ZN(n398) );
  XNOR2_X2 U475 ( .A(n510), .B(KEYINPUT33), .ZN(n690) );
  INV_X1 U476 ( .A(n375), .ZN(n702) );
  XNOR2_X2 U477 ( .A(n400), .B(KEYINPUT32), .ZN(n506) );
  INV_X1 U478 ( .A(n563), .ZN(n402) );
  XNOR2_X1 U479 ( .A(n416), .B(n378), .ZN(n563) );
  XOR2_X1 U480 ( .A(n619), .B(KEYINPUT65), .Z(n403) );
  AND2_X1 U481 ( .A1(n700), .A2(n699), .ZN(n404) );
  INV_X1 U482 ( .A(n703), .ZN(n505) );
  NOR2_X1 U483 ( .A1(n612), .A2(n611), .ZN(n613) );
  INV_X1 U484 ( .A(KEYINPUT79), .ZN(n660) );
  XNOR2_X1 U485 ( .A(G107), .B(G104), .ZN(n407) );
  XNOR2_X1 U486 ( .A(n407), .B(n406), .ZN(n754) );
  XNOR2_X2 U487 ( .A(KEYINPUT4), .B(G101), .ZN(n473) );
  XNOR2_X1 U488 ( .A(n473), .B(KEYINPUT71), .ZN(n408) );
  XNOR2_X1 U489 ( .A(n754), .B(n408), .ZN(n482) );
  XNOR2_X1 U490 ( .A(n409), .B(n482), .ZN(n414) );
  XNOR2_X1 U491 ( .A(n410), .B(KEYINPUT3), .ZN(n412) );
  XNOR2_X1 U492 ( .A(n412), .B(n411), .ZN(n477) );
  XNOR2_X1 U493 ( .A(KEYINPUT16), .B(G122), .ZN(n413) );
  XNOR2_X1 U494 ( .A(n477), .B(n413), .ZN(n757) );
  XNOR2_X1 U495 ( .A(n414), .B(n757), .ZN(n625) );
  INV_X1 U496 ( .A(n618), .ZN(n415) );
  NOR2_X1 U497 ( .A1(n625), .A2(n415), .ZN(n416) );
  INV_X1 U498 ( .A(G902), .ZN(n496) );
  INV_X1 U499 ( .A(G237), .ZN(n417) );
  NAND2_X1 U500 ( .A1(n496), .A2(n417), .ZN(n419) );
  NAND2_X1 U501 ( .A1(n419), .A2(G210), .ZN(n418) );
  NAND2_X1 U502 ( .A1(n419), .A2(G214), .ZN(n420) );
  XNOR2_X1 U503 ( .A(n420), .B(KEYINPUT91), .ZN(n679) );
  NAND2_X1 U504 ( .A1(G237), .A2(G234), .ZN(n421) );
  XNOR2_X1 U505 ( .A(n421), .B(KEYINPUT14), .ZN(n551) );
  AND2_X1 U506 ( .A1(n749), .A2(G902), .ZN(n423) );
  INV_X1 U507 ( .A(G898), .ZN(n422) );
  NAND2_X1 U508 ( .A1(n423), .A2(n422), .ZN(n425) );
  NAND2_X1 U509 ( .A1(n368), .A2(G952), .ZN(n424) );
  NAND2_X1 U510 ( .A1(n425), .A2(n424), .ZN(n426) );
  AND2_X1 U511 ( .A1(n551), .A2(n426), .ZN(n427) );
  XNOR2_X2 U512 ( .A(n428), .B(n380), .ZN(n508) );
  XOR2_X1 U513 ( .A(G113), .B(G104), .Z(n430) );
  XNOR2_X1 U514 ( .A(G143), .B(G122), .ZN(n429) );
  XNOR2_X1 U515 ( .A(n430), .B(n429), .ZN(n434) );
  XOR2_X1 U516 ( .A(KEYINPUT12), .B(KEYINPUT100), .Z(n432) );
  XNOR2_X1 U517 ( .A(KEYINPUT11), .B(KEYINPUT98), .ZN(n431) );
  XNOR2_X1 U518 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U519 ( .A(n434), .B(n433), .ZN(n437) );
  XNOR2_X1 U520 ( .A(n436), .B(n435), .ZN(n645) );
  XNOR2_X1 U521 ( .A(n437), .B(n645), .ZN(n442) );
  XNOR2_X2 U522 ( .A(KEYINPUT69), .B(G131), .ZN(n469) );
  XNOR2_X1 U523 ( .A(n469), .B(KEYINPUT99), .ZN(n440) );
  XNOR2_X1 U524 ( .A(KEYINPUT74), .B(n438), .ZN(n474) );
  NAND2_X1 U525 ( .A1(n474), .A2(G214), .ZN(n439) );
  XNOR2_X1 U526 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U527 ( .A(n442), .B(n441), .ZN(n713) );
  NAND2_X1 U528 ( .A1(n713), .A2(n496), .ZN(n446) );
  XOR2_X1 U529 ( .A(KEYINPUT13), .B(KEYINPUT102), .Z(n444) );
  XNOR2_X1 U530 ( .A(KEYINPUT101), .B(G475), .ZN(n443) );
  XOR2_X1 U531 ( .A(n444), .B(n443), .Z(n445) );
  XNOR2_X1 U532 ( .A(n446), .B(n445), .ZN(n529) );
  XOR2_X1 U533 ( .A(KEYINPUT9), .B(G122), .Z(n448) );
  XNOR2_X1 U534 ( .A(n448), .B(n447), .ZN(n451) );
  INV_X1 U535 ( .A(G134), .ZN(n449) );
  XNOR2_X1 U536 ( .A(n451), .B(n471), .ZN(n457) );
  NAND2_X1 U537 ( .A1(n377), .A2(G234), .ZN(n453) );
  INV_X1 U538 ( .A(KEYINPUT8), .ZN(n452) );
  NAND2_X1 U539 ( .A1(n491), .A2(G217), .ZN(n455) );
  XNOR2_X1 U540 ( .A(KEYINPUT103), .B(KEYINPUT7), .ZN(n454) );
  XNOR2_X1 U541 ( .A(n455), .B(n454), .ZN(n456) );
  NAND2_X1 U542 ( .A1(n709), .A2(n496), .ZN(n458) );
  XNOR2_X1 U543 ( .A(n458), .B(G478), .ZN(n525) );
  OR2_X1 U544 ( .A1(n529), .A2(n525), .ZN(n683) );
  INV_X1 U545 ( .A(n683), .ZN(n464) );
  NAND2_X1 U546 ( .A1(n618), .A2(G234), .ZN(n459) );
  NAND2_X1 U547 ( .A1(n497), .A2(G221), .ZN(n462) );
  INV_X1 U548 ( .A(KEYINPUT93), .ZN(n460) );
  XNOR2_X1 U549 ( .A(n460), .B(KEYINPUT21), .ZN(n461) );
  XNOR2_X1 U550 ( .A(n462), .B(n461), .ZN(n667) );
  INV_X1 U551 ( .A(n667), .ZN(n463) );
  INV_X1 U552 ( .A(G137), .ZN(n468) );
  XNOR2_X1 U553 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U554 ( .A(KEYINPUT94), .B(KEYINPUT5), .ZN(n472) );
  XNOR2_X1 U555 ( .A(n473), .B(n472), .ZN(n476) );
  AND2_X1 U556 ( .A1(n474), .A2(G210), .ZN(n475) );
  XNOR2_X1 U557 ( .A(G472), .B(KEYINPUT95), .ZN(n478) );
  NAND2_X1 U558 ( .A1(n377), .A2(G227), .ZN(n479) );
  XNOR2_X1 U559 ( .A(n479), .B(G140), .ZN(n481) );
  XNOR2_X1 U560 ( .A(KEYINPUT75), .B(KEYINPUT76), .ZN(n480) );
  XNOR2_X1 U561 ( .A(n481), .B(n480), .ZN(n483) );
  XNOR2_X1 U562 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U563 ( .A(n485), .B(n484), .ZN(n722) );
  OR2_X2 U564 ( .A1(n722), .A2(G902), .ZN(n487) );
  INV_X1 U565 ( .A(G469), .ZN(n486) );
  XNOR2_X2 U566 ( .A(n487), .B(n486), .ZN(n581) );
  XOR2_X1 U567 ( .A(G137), .B(G119), .Z(n489) );
  XOR2_X1 U568 ( .A(n489), .B(n488), .Z(n490) );
  XNOR2_X1 U569 ( .A(n490), .B(n645), .ZN(n495) );
  XOR2_X1 U570 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n493) );
  NAND2_X1 U571 ( .A1(G221), .A2(n491), .ZN(n492) );
  XNOR2_X1 U572 ( .A(n493), .B(n492), .ZN(n494) );
  NAND2_X1 U573 ( .A1(n634), .A2(n496), .ZN(n501) );
  XOR2_X1 U574 ( .A(n501), .B(n500), .Z(n554) );
  OR2_X1 U575 ( .A1(n595), .A2(n554), .ZN(n498) );
  XNOR2_X1 U576 ( .A(n501), .B(n500), .ZN(n666) );
  AND2_X1 U577 ( .A1(n669), .A2(n666), .ZN(n502) );
  AND2_X1 U578 ( .A1(n595), .A2(n502), .ZN(n503) );
  AND2_X1 U579 ( .A1(n384), .A2(n503), .ZN(n703) );
  NAND2_X1 U580 ( .A1(n506), .A2(n505), .ZN(n507) );
  XNOR2_X1 U581 ( .A(n507), .B(KEYINPUT86), .ZN(n537) );
  BUF_X1 U582 ( .A(n508), .Z(n509) );
  OR2_X2 U583 ( .A1(n595), .A2(n662), .ZN(n517) );
  OR2_X2 U584 ( .A1(n517), .A2(n558), .ZN(n510) );
  NAND2_X1 U585 ( .A1(n529), .A2(n525), .ZN(n511) );
  XNOR2_X1 U586 ( .A(n511), .B(KEYINPUT106), .ZN(n602) );
  INV_X1 U587 ( .A(n602), .ZN(n512) );
  OR2_X2 U588 ( .A1(n537), .A2(n641), .ZN(n514) );
  NAND2_X1 U589 ( .A1(n514), .A2(KEYINPUT44), .ZN(n534) );
  XNOR2_X1 U590 ( .A(n379), .B(KEYINPUT83), .ZN(n516) );
  AND2_X1 U591 ( .A1(n595), .A2(n554), .ZN(n515) );
  NAND2_X1 U592 ( .A1(n516), .A2(n515), .ZN(n642) );
  INV_X1 U593 ( .A(n509), .ZN(n522) );
  OR2_X1 U594 ( .A1(n517), .A2(n669), .ZN(n674) );
  OR2_X1 U595 ( .A1(n522), .A2(n674), .ZN(n519) );
  XOR2_X1 U596 ( .A(KEYINPUT97), .B(KEYINPUT31), .Z(n518) );
  XNOR2_X1 U597 ( .A(n519), .B(n518), .ZN(n743) );
  OR2_X1 U598 ( .A1(n581), .A2(n662), .ZN(n570) );
  INV_X1 U599 ( .A(n570), .ZN(n520) );
  NAND2_X1 U600 ( .A1(n520), .A2(n669), .ZN(n521) );
  OR2_X1 U601 ( .A1(n522), .A2(n521), .ZN(n524) );
  INV_X1 U602 ( .A(KEYINPUT96), .ZN(n523) );
  XNOR2_X1 U603 ( .A(n524), .B(n523), .ZN(n731) );
  OR2_X1 U604 ( .A1(n743), .A2(n731), .ZN(n531) );
  INV_X1 U605 ( .A(n525), .ZN(n528) );
  OR2_X1 U606 ( .A1(n529), .A2(n528), .ZN(n527) );
  INV_X1 U607 ( .A(KEYINPUT104), .ZN(n526) );
  XNOR2_X1 U608 ( .A(n527), .B(n526), .ZN(n744) );
  AND2_X1 U609 ( .A1(n529), .A2(n528), .ZN(n740) );
  OR2_X1 U610 ( .A1(n744), .A2(n740), .ZN(n685) );
  INV_X1 U611 ( .A(KEYINPUT77), .ZN(n530) );
  XNOR2_X1 U612 ( .A(n685), .B(n530), .ZN(n598) );
  NAND2_X1 U613 ( .A1(n531), .A2(n598), .ZN(n532) );
  AND2_X1 U614 ( .A1(n642), .A2(n532), .ZN(n533) );
  NAND2_X1 U615 ( .A1(n534), .A2(n533), .ZN(n536) );
  INV_X1 U616 ( .A(KEYINPUT84), .ZN(n535) );
  BUF_X1 U617 ( .A(n537), .Z(n538) );
  XNOR2_X1 U618 ( .A(n538), .B(KEYINPUT85), .ZN(n541) );
  OR2_X1 U619 ( .A1(n641), .A2(KEYINPUT44), .ZN(n539) );
  XNOR2_X1 U620 ( .A(n539), .B(KEYINPUT67), .ZN(n540) );
  NAND2_X1 U621 ( .A1(n541), .A2(n540), .ZN(n542) );
  NAND2_X1 U622 ( .A1(n543), .A2(n542), .ZN(n546) );
  INV_X1 U623 ( .A(KEYINPUT64), .ZN(n544) );
  XNOR2_X2 U624 ( .A(n546), .B(n545), .ZN(n655) );
  NAND2_X1 U625 ( .A1(G902), .A2(n551), .ZN(n547) );
  NOR2_X1 U626 ( .A1(G900), .A2(n547), .ZN(n548) );
  NAND2_X1 U627 ( .A1(n749), .A2(n548), .ZN(n550) );
  INV_X1 U628 ( .A(KEYINPUT107), .ZN(n549) );
  XNOR2_X1 U629 ( .A(n550), .B(n549), .ZN(n553) );
  AND2_X1 U630 ( .A1(n551), .A2(G952), .ZN(n696) );
  NAND2_X1 U631 ( .A1(n696), .A2(n368), .ZN(n552) );
  NAND2_X1 U632 ( .A1(n553), .A2(n552), .ZN(n567) );
  NOR2_X1 U633 ( .A1(n667), .A2(n554), .ZN(n555) );
  NAND2_X1 U634 ( .A1(n567), .A2(n555), .ZN(n578) );
  INV_X1 U635 ( .A(n578), .ZN(n556) );
  NAND2_X1 U636 ( .A1(n740), .A2(n556), .ZN(n557) );
  INV_X1 U637 ( .A(KEYINPUT108), .ZN(n559) );
  XNOR2_X1 U638 ( .A(n560), .B(n559), .ZN(n592) );
  NAND2_X1 U639 ( .A1(n595), .A2(n592), .ZN(n561) );
  NOR2_X1 U640 ( .A1(n679), .A2(n561), .ZN(n562) );
  XNOR2_X1 U641 ( .A(n562), .B(KEYINPUT43), .ZN(n565) );
  BUF_X1 U642 ( .A(n563), .Z(n601) );
  INV_X1 U643 ( .A(n601), .ZN(n564) );
  NOR2_X1 U644 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U645 ( .A(n566), .B(KEYINPUT109), .ZN(n763) );
  AND2_X1 U646 ( .A1(n568), .A2(n567), .ZN(n572) );
  INV_X1 U647 ( .A(KEYINPUT110), .ZN(n569) );
  XNOR2_X1 U648 ( .A(n570), .B(n569), .ZN(n571) );
  NAND2_X1 U649 ( .A1(n572), .A2(n571), .ZN(n604) );
  INV_X1 U650 ( .A(KEYINPUT38), .ZN(n573) );
  NAND2_X1 U651 ( .A1(n574), .A2(n744), .ZN(n640) );
  AND2_X1 U652 ( .A1(n763), .A2(n640), .ZN(n615) );
  NAND2_X1 U653 ( .A1(n574), .A2(n740), .ZN(n575) );
  OR2_X1 U654 ( .A1(n680), .A2(n679), .ZN(n687) );
  OR2_X1 U655 ( .A1(n687), .A2(n683), .ZN(n577) );
  XOR2_X1 U656 ( .A(KEYINPUT111), .B(KEYINPUT41), .Z(n576) );
  OR2_X1 U657 ( .A1(n669), .A2(n578), .ZN(n580) );
  INV_X1 U658 ( .A(KEYINPUT28), .ZN(n579) );
  XNOR2_X1 U659 ( .A(n580), .B(n579), .ZN(n583) );
  INV_X1 U660 ( .A(n581), .ZN(n582) );
  AND2_X1 U661 ( .A1(n583), .A2(n582), .ZN(n599) );
  NAND2_X1 U662 ( .A1(n698), .A2(n599), .ZN(n586) );
  INV_X1 U663 ( .A(KEYINPUT112), .ZN(n584) );
  XNOR2_X1 U664 ( .A(n584), .B(KEYINPUT42), .ZN(n585) );
  XNOR2_X1 U665 ( .A(n586), .B(n585), .ZN(n762) );
  INV_X1 U666 ( .A(n762), .ZN(n587) );
  NAND2_X1 U667 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U668 ( .A(n589), .B(KEYINPUT46), .ZN(n612) );
  INV_X1 U669 ( .A(n590), .ZN(n591) );
  NAND2_X1 U670 ( .A1(n592), .A2(n591), .ZN(n594) );
  XNOR2_X1 U671 ( .A(KEYINPUT36), .B(KEYINPUT87), .ZN(n593) );
  XNOR2_X1 U672 ( .A(n594), .B(n593), .ZN(n596) );
  INV_X1 U673 ( .A(n595), .ZN(n663) );
  AND2_X1 U674 ( .A1(n596), .A2(n663), .ZN(n746) );
  XNOR2_X1 U675 ( .A(n746), .B(KEYINPUT81), .ZN(n610) );
  XOR2_X1 U676 ( .A(KEYINPUT47), .B(KEYINPUT68), .Z(n597) );
  AND2_X1 U677 ( .A1(n598), .A2(n597), .ZN(n600) );
  NAND2_X1 U678 ( .A1(n600), .A2(n738), .ZN(n605) );
  OR2_X1 U679 ( .A1(n602), .A2(n601), .ZN(n603) );
  OR2_X1 U680 ( .A1(n604), .A2(n603), .ZN(n639) );
  NAND2_X1 U681 ( .A1(n605), .A2(n639), .ZN(n608) );
  NAND2_X1 U682 ( .A1(n738), .A2(n685), .ZN(n606) );
  AND2_X1 U683 ( .A1(n606), .A2(KEYINPUT47), .ZN(n607) );
  NOR2_X1 U684 ( .A1(n608), .A2(n607), .ZN(n609) );
  NAND2_X1 U685 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U686 ( .A(n613), .B(KEYINPUT48), .ZN(n614) );
  NAND2_X1 U687 ( .A1(n615), .A2(n614), .ZN(n622) );
  XNOR2_X2 U688 ( .A(n622), .B(KEYINPUT80), .ZN(n656) );
  INV_X1 U689 ( .A(n656), .ZN(n616) );
  INV_X1 U690 ( .A(KEYINPUT2), .ZN(n621) );
  OR2_X1 U691 ( .A1(n618), .A2(n621), .ZN(n619) );
  NAND2_X1 U692 ( .A1(n620), .A2(n403), .ZN(n624) );
  OR2_X1 U693 ( .A1(n622), .A2(n621), .ZN(n623) );
  AND2_X2 U694 ( .A1(n624), .A2(n658), .ZN(n719) );
  NAND2_X1 U695 ( .A1(n719), .A2(G210), .ZN(n629) );
  BUF_X1 U696 ( .A(n625), .Z(n626) );
  XNOR2_X1 U697 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n627) );
  XNOR2_X1 U698 ( .A(n626), .B(n627), .ZN(n628) );
  XNOR2_X1 U699 ( .A(n629), .B(n628), .ZN(n631) );
  INV_X1 U700 ( .A(G952), .ZN(n630) );
  NAND2_X1 U701 ( .A1(n631), .A2(n725), .ZN(n633) );
  INV_X1 U702 ( .A(KEYINPUT56), .ZN(n632) );
  XNOR2_X1 U703 ( .A(n633), .B(n632), .ZN(G51) );
  NAND2_X1 U704 ( .A1(n719), .A2(G217), .ZN(n635) );
  XNOR2_X1 U705 ( .A(n635), .B(n634), .ZN(n636) );
  NAND2_X1 U706 ( .A1(n636), .A2(n725), .ZN(n638) );
  INV_X1 U707 ( .A(KEYINPUT124), .ZN(n637) );
  XNOR2_X1 U708 ( .A(n638), .B(n637), .ZN(G66) );
  XNOR2_X1 U709 ( .A(n639), .B(G143), .ZN(G45) );
  XNOR2_X1 U710 ( .A(n640), .B(G134), .ZN(G36) );
  XOR2_X1 U711 ( .A(n374), .B(G122), .Z(G24) );
  XNOR2_X1 U712 ( .A(n642), .B(G101), .ZN(G3) );
  XOR2_X1 U713 ( .A(KEYINPUT4), .B(KEYINPUT125), .Z(n644) );
  XNOR2_X1 U714 ( .A(n645), .B(n644), .ZN(n646) );
  XNOR2_X1 U715 ( .A(n643), .B(n646), .ZN(n648) );
  XNOR2_X1 U716 ( .A(n656), .B(n648), .ZN(n647) );
  NAND2_X1 U717 ( .A1(n647), .A2(n368), .ZN(n654) );
  XNOR2_X1 U718 ( .A(n648), .B(G227), .ZN(n649) );
  XNOR2_X1 U719 ( .A(n649), .B(KEYINPUT126), .ZN(n650) );
  NAND2_X1 U720 ( .A1(n650), .A2(G900), .ZN(n651) );
  XOR2_X1 U721 ( .A(KEYINPUT127), .B(n651), .Z(n652) );
  NAND2_X1 U722 ( .A1(n749), .A2(n652), .ZN(n653) );
  NAND2_X1 U723 ( .A1(n654), .A2(n653), .ZN(G72) );
  NOR2_X1 U724 ( .A1(n656), .A2(n655), .ZN(n657) );
  OR2_X1 U725 ( .A1(n657), .A2(KEYINPUT2), .ZN(n659) );
  NAND2_X1 U726 ( .A1(n659), .A2(n658), .ZN(n661) );
  XNOR2_X1 U727 ( .A(n661), .B(n660), .ZN(n701) );
  INV_X1 U728 ( .A(n662), .ZN(n664) );
  NOR2_X1 U729 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U730 ( .A(n665), .B(KEYINPUT50), .ZN(n672) );
  AND2_X1 U731 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U732 ( .A(n668), .B(KEYINPUT49), .ZN(n670) );
  NAND2_X1 U733 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U734 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U735 ( .A(n673), .B(KEYINPUT117), .ZN(n675) );
  AND2_X1 U736 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U737 ( .A(KEYINPUT51), .B(n676), .ZN(n677) );
  NAND2_X1 U738 ( .A1(n677), .A2(n698), .ZN(n678) );
  XOR2_X1 U739 ( .A(KEYINPUT118), .B(n678), .Z(n694) );
  AND2_X1 U740 ( .A1(n680), .A2(n679), .ZN(n681) );
  XOR2_X1 U741 ( .A(KEYINPUT119), .B(n681), .Z(n682) );
  NOR2_X1 U742 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U743 ( .A(n684), .B(KEYINPUT120), .ZN(n689) );
  INV_X1 U744 ( .A(n685), .ZN(n686) );
  NOR2_X1 U745 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U746 ( .A1(n689), .A2(n688), .ZN(n692) );
  INV_X1 U747 ( .A(n690), .ZN(n691) );
  NOR2_X1 U748 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U749 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U750 ( .A(KEYINPUT52), .B(n695), .Z(n697) );
  NAND2_X1 U751 ( .A1(n697), .A2(n696), .ZN(n700) );
  NAND2_X1 U752 ( .A1(n690), .A2(n698), .ZN(n699) );
  XOR2_X1 U753 ( .A(n702), .B(G119), .Z(G21) );
  XOR2_X1 U754 ( .A(G110), .B(n703), .Z(G12) );
  NAND2_X1 U755 ( .A1(n719), .A2(G472), .ZN(n706) );
  XOR2_X1 U756 ( .A(KEYINPUT62), .B(n704), .Z(n705) );
  XNOR2_X1 U757 ( .A(n706), .B(n705), .ZN(n707) );
  NAND2_X1 U758 ( .A1(n707), .A2(n725), .ZN(n708) );
  XNOR2_X1 U759 ( .A(n708), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U760 ( .A1(n719), .A2(G478), .ZN(n710) );
  XNOR2_X1 U761 ( .A(n710), .B(n709), .ZN(n711) );
  NAND2_X1 U762 ( .A1(n711), .A2(n725), .ZN(n712) );
  XNOR2_X1 U763 ( .A(n712), .B(KEYINPUT123), .ZN(G63) );
  NAND2_X1 U764 ( .A1(n719), .A2(G475), .ZN(n715) );
  XOR2_X1 U765 ( .A(KEYINPUT59), .B(n713), .Z(n714) );
  XNOR2_X1 U766 ( .A(n715), .B(n714), .ZN(n716) );
  NAND2_X1 U767 ( .A1(n716), .A2(n725), .ZN(n718) );
  INV_X1 U768 ( .A(KEYINPUT60), .ZN(n717) );
  XNOR2_X1 U769 ( .A(n718), .B(n717), .ZN(G60) );
  NAND2_X1 U770 ( .A1(n719), .A2(G469), .ZN(n724) );
  XOR2_X1 U771 ( .A(KEYINPUT122), .B(KEYINPUT57), .Z(n720) );
  XNOR2_X1 U772 ( .A(n720), .B(KEYINPUT58), .ZN(n721) );
  XNOR2_X1 U773 ( .A(n722), .B(n721), .ZN(n723) );
  XNOR2_X1 U774 ( .A(n724), .B(n723), .ZN(n727) );
  INV_X1 U775 ( .A(n725), .ZN(n726) );
  NOR2_X1 U776 ( .A1(n727), .A2(n726), .ZN(G54) );
  XOR2_X1 U777 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n729) );
  NAND2_X1 U778 ( .A1(n740), .A2(n731), .ZN(n728) );
  XNOR2_X1 U779 ( .A(n729), .B(n728), .ZN(n730) );
  XNOR2_X1 U780 ( .A(G104), .B(n730), .ZN(G6) );
  XOR2_X1 U781 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n733) );
  NAND2_X1 U782 ( .A1(n731), .A2(n744), .ZN(n732) );
  XNOR2_X1 U783 ( .A(n733), .B(n732), .ZN(n734) );
  XNOR2_X1 U784 ( .A(G107), .B(n734), .ZN(G9) );
  XOR2_X1 U785 ( .A(KEYINPUT29), .B(KEYINPUT115), .Z(n736) );
  NAND2_X1 U786 ( .A1(n738), .A2(n744), .ZN(n735) );
  XNOR2_X1 U787 ( .A(n736), .B(n735), .ZN(n737) );
  XOR2_X1 U788 ( .A(G128), .B(n737), .Z(G30) );
  NAND2_X1 U789 ( .A1(n738), .A2(n740), .ZN(n739) );
  XNOR2_X1 U790 ( .A(n739), .B(G146), .ZN(G48) );
  NAND2_X1 U791 ( .A1(n743), .A2(n740), .ZN(n741) );
  XNOR2_X1 U792 ( .A(n741), .B(KEYINPUT116), .ZN(n742) );
  XNOR2_X1 U793 ( .A(G113), .B(n742), .ZN(G15) );
  NAND2_X1 U794 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U795 ( .A(n745), .B(G116), .ZN(G18) );
  XNOR2_X1 U796 ( .A(G125), .B(n746), .ZN(n747) );
  XNOR2_X1 U797 ( .A(n747), .B(KEYINPUT37), .ZN(G27) );
  INV_X1 U798 ( .A(n376), .ZN(n748) );
  NAND2_X1 U799 ( .A1(n748), .A2(n368), .ZN(n753) );
  NAND2_X1 U800 ( .A1(n749), .A2(G224), .ZN(n750) );
  XNOR2_X1 U801 ( .A(KEYINPUT61), .B(n750), .ZN(n751) );
  NAND2_X1 U802 ( .A1(n751), .A2(G898), .ZN(n752) );
  NAND2_X1 U803 ( .A1(n753), .A2(n752), .ZN(n761) );
  BUF_X1 U804 ( .A(n754), .Z(n755) );
  XNOR2_X1 U805 ( .A(n755), .B(G101), .ZN(n756) );
  XNOR2_X1 U806 ( .A(n757), .B(n756), .ZN(n759) );
  NOR2_X1 U807 ( .A1(n368), .A2(G898), .ZN(n758) );
  NOR2_X1 U808 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U809 ( .A(n761), .B(n760), .ZN(G69) );
  XOR2_X1 U810 ( .A(G137), .B(n762), .Z(G39) );
  XNOR2_X1 U811 ( .A(G140), .B(n763), .ZN(G42) );
endmodule

