//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 1 0 0 1 1 1 1 1 0 1 0 0 1 0 1 0 0 1 0 0 0 0 0 1 1 1 1 1 0 0 0 1 1 0 1 0 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:50 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n546, new_n548, new_n549, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n628, new_n629, new_n632,
    new_n634, new_n635, new_n636, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1178,
    new_n1179, new_n1180, new_n1181;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT64), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT65), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AND3_X1   g035(.A1(KEYINPUT66), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n461));
  AOI21_X1  g036(.A(KEYINPUT3), .B1(KEYINPUT66), .B2(G2104), .ZN(new_n462));
  OAI211_X1 g037(.A(G137), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G101), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n460), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(G125), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n460), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n466), .A2(new_n471), .ZN(G160));
  NAND2_X1  g047(.A1(KEYINPUT66), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g050(.A1(KEYINPUT66), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n477), .A2(new_n460), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  AOI22_X1  g056(.A1(G124), .A2(new_n479), .B1(new_n481), .B2(G136), .ZN(new_n482));
  INV_X1    g057(.A(G2104), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n460), .A2(G100), .ZN(new_n484));
  NAND2_X1  g059(.A1(G112), .A2(G2105), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT67), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n482), .A2(new_n487), .ZN(G162));
  NAND2_X1  g063(.A1(KEYINPUT4), .A2(G138), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n489), .B1(new_n475), .B2(new_n476), .ZN(new_n490));
  AND2_X1   g065(.A1(G102), .A2(G2104), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n460), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G126), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n493), .B1(new_n475), .B2(new_n476), .ZN(new_n494));
  NAND2_X1  g069(.A1(G114), .A2(G2104), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(G2105), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  OAI211_X1 g072(.A(G138), .B(new_n460), .C1(new_n467), .C2(new_n468), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n492), .A2(new_n497), .A3(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  OR2_X1    g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n505), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  OR2_X1    g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G50), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  AND2_X1   g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  AND2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  OAI22_X1  g093(.A1(new_n515), .A2(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n513), .B1(new_n514), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n508), .A2(new_n520), .ZN(G166));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  INV_X1    g098(.A(new_n512), .ZN(new_n524));
  XOR2_X1   g099(.A(KEYINPUT68), .B(G51), .Z(new_n525));
  OAI21_X1  g100(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n516), .A2(new_n515), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n510), .A2(new_n511), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G89), .ZN(new_n529));
  NAND2_X1  g104(.A1(G63), .A2(G651), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n527), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n526), .A2(new_n531), .ZN(G168));
  AOI22_X1  g107(.A1(new_n505), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n533), .A2(new_n507), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n512), .A2(G52), .ZN(new_n535));
  INV_X1    g110(.A(G90), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n536), .B2(new_n519), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n534), .A2(new_n537), .ZN(G171));
  AOI22_X1  g113(.A1(new_n505), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n539), .A2(new_n507), .ZN(new_n540));
  INV_X1    g115(.A(new_n519), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n541), .A2(G81), .B1(G43), .B2(new_n512), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(G153));
  AND3_X1   g120(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G36), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n546), .A2(new_n549), .ZN(G188));
  INV_X1    g125(.A(G65), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT70), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n505), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n527), .A2(KEYINPUT70), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n551), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  AND2_X1   g130(.A1(G78), .A2(G543), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT71), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n507), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g134(.A(KEYINPUT71), .B1(new_n555), .B2(new_n556), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  INV_X1    g137(.A(G53), .ZN(new_n563));
  OAI211_X1 g138(.A(KEYINPUT69), .B(new_n562), .C1(new_n524), .C2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n541), .A2(G91), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT69), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n563), .B1(new_n566), .B2(KEYINPUT9), .ZN(new_n567));
  OAI211_X1 g142(.A(new_n512), .B(new_n567), .C1(new_n566), .C2(KEYINPUT9), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n564), .A2(new_n565), .A3(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n561), .A2(new_n570), .ZN(G299));
  INV_X1    g146(.A(G171), .ZN(G301));
  INV_X1    g147(.A(G168), .ZN(G286));
  INV_X1    g148(.A(G166), .ZN(G303));
  INV_X1    g149(.A(KEYINPUT73), .ZN(new_n575));
  INV_X1    g150(.A(G74), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n503), .A2(new_n576), .A3(new_n504), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n575), .B1(new_n577), .B2(G651), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n575), .A3(G651), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT72), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n512), .A2(new_n582), .A3(G49), .ZN(new_n583));
  OAI211_X1 g158(.A(G49), .B(G543), .C1(new_n517), .C2(new_n518), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(KEYINPUT72), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n583), .A2(new_n585), .B1(new_n541), .B2(G87), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n581), .A2(new_n586), .ZN(G288));
  NAND3_X1  g162(.A1(new_n512), .A2(KEYINPUT75), .A3(G48), .ZN(new_n588));
  OAI211_X1 g163(.A(G48), .B(G543), .C1(new_n517), .C2(new_n518), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT75), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(G73), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G61), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n527), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n588), .A2(new_n591), .B1(new_n594), .B2(G651), .ZN(new_n595));
  INV_X1    g170(.A(G86), .ZN(new_n596));
  OAI21_X1  g171(.A(KEYINPUT74), .B1(new_n519), .B2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT74), .ZN(new_n598));
  NAND4_X1  g173(.A1(new_n505), .A2(new_n528), .A3(new_n598), .A4(G86), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  AND2_X1   g175(.A1(new_n595), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(G305));
  AOI22_X1  g177(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n603), .A2(new_n507), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT76), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n604), .B(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT77), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n541), .A2(G85), .B1(G47), .B2(new_n512), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n607), .B1(new_n606), .B2(new_n608), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(G290));
  INV_X1    g188(.A(G868), .ZN(new_n614));
  NOR2_X1   g189(.A1(G301), .A2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(G92), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n519), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT10), .ZN(new_n618));
  INV_X1    g193(.A(G66), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n619), .B1(new_n553), .B2(new_n554), .ZN(new_n620));
  AND2_X1   g195(.A1(G79), .A2(G543), .ZN(new_n621));
  OAI21_X1  g196(.A(G651), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n512), .A2(G54), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n618), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n615), .B1(new_n625), .B2(new_n614), .ZN(G284));
  AOI21_X1  g201(.A(new_n615), .B1(new_n625), .B2(new_n614), .ZN(G321));
  NOR2_X1   g202(.A1(G286), .A2(new_n614), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n569), .B1(new_n559), .B2(new_n560), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n628), .B1(new_n629), .B2(new_n614), .ZN(G280));
  XOR2_X1   g205(.A(G280), .B(KEYINPUT78), .Z(G297));
  INV_X1    g206(.A(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n625), .B1(new_n632), .B2(G860), .ZN(G148));
  NAND2_X1  g208(.A1(new_n544), .A2(new_n614), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n625), .A2(new_n632), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n634), .B1(new_n635), .B2(new_n614), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT79), .ZN(G323));
  XNOR2_X1  g212(.A(G323), .B(KEYINPUT11), .ZN(G282));
  MUX2_X1   g213(.A(G99), .B(G111), .S(G2105), .Z(new_n639));
  AOI22_X1  g214(.A1(new_n479), .A2(G123), .B1(G2104), .B2(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(G135), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n640), .B1(new_n641), .B2(new_n480), .ZN(new_n642));
  INV_X1    g217(.A(G2096), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n460), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT12), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT13), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n648), .A2(G2100), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n648), .A2(G2100), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n644), .A2(new_n649), .A3(new_n650), .ZN(G156));
  INV_X1    g226(.A(KEYINPUT14), .ZN(new_n652));
  XOR2_X1   g227(.A(KEYINPUT15), .B(G2435), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2438), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2427), .ZN(new_n655));
  INV_X1    g230(.A(G2430), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n652), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n657), .B1(new_n656), .B2(new_n655), .ZN(new_n658));
  XOR2_X1   g233(.A(G2451), .B(G2454), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT16), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT80), .ZN(new_n661));
  XOR2_X1   g236(.A(G2443), .B(G2446), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n658), .B(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G1341), .B(G1348), .Z(new_n665));
  NOR2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT81), .ZN(new_n667));
  INV_X1    g242(.A(G14), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n668), .B1(new_n664), .B2(new_n665), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(G401));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  XNOR2_X1  g247(.A(G2072), .B(G2078), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2067), .B(G2678), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(KEYINPUT82), .B(KEYINPUT18), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n672), .A2(KEYINPUT17), .A3(new_n673), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n672), .B1(KEYINPUT17), .B2(new_n673), .ZN(new_n679));
  INV_X1    g254(.A(new_n674), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n678), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n672), .A2(new_n674), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n673), .B1(new_n682), .B2(KEYINPUT17), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n677), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(new_n643), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G2100), .ZN(G227));
  XNOR2_X1  g261(.A(G1971), .B(G1976), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT83), .B(KEYINPUT19), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(G1956), .B(G2474), .Z(new_n690));
  XOR2_X1   g265(.A(G1961), .B(G1966), .Z(new_n691));
  AND2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT20), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n690), .A2(new_n691), .ZN(new_n695));
  NOR3_X1   g270(.A1(new_n689), .A2(new_n692), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n689), .B2(new_n695), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1991), .B(G1996), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1981), .B(G1986), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n700), .B(new_n703), .ZN(G229));
  NOR2_X1   g279(.A1(G16), .A2(G19), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(new_n544), .B2(G16), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(G1341), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT31), .B(G11), .Z(new_n708));
  INV_X1    g283(.A(G29), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n642), .A2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(G28), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n711), .A2(KEYINPUT30), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT91), .Z(new_n713));
  AOI21_X1  g288(.A(G29), .B1(new_n711), .B2(KEYINPUT30), .ZN(new_n714));
  AOI211_X1 g289(.A(new_n708), .B(new_n710), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G16), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G5), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G171), .B2(new_n716), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT24), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G34), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n709), .B1(new_n719), .B2(G34), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(KEYINPUT89), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(KEYINPUT89), .B2(new_n721), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(G160), .B2(G29), .ZN(new_n724));
  OAI221_X1 g299(.A(new_n715), .B1(G1961), .B2(new_n718), .C1(G2084), .C2(new_n724), .ZN(new_n725));
  AOI211_X1 g300(.A(new_n707), .B(new_n725), .C1(G2084), .C2(new_n724), .ZN(new_n726));
  NOR2_X1   g301(.A1(G4), .A2(G16), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(new_n625), .B2(G16), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(G1348), .ZN(new_n730));
  NOR2_X1   g305(.A1(G27), .A2(G29), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G164), .B2(G29), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n729), .A2(new_n730), .B1(G2078), .B2(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n732), .A2(G2078), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(new_n728), .B2(G1348), .ZN(new_n735));
  NOR2_X1   g310(.A1(G168), .A2(new_n716), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n716), .B2(G21), .ZN(new_n737));
  INV_X1    g312(.A(G1966), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n737), .A2(new_n738), .B1(G1961), .B2(new_n718), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(new_n738), .B2(new_n737), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n709), .A2(G26), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT28), .Z(new_n742));
  MUX2_X1   g317(.A(G104), .B(G116), .S(G2105), .Z(new_n743));
  AOI22_X1  g318(.A1(new_n479), .A2(G128), .B1(G2104), .B2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(G140), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n744), .B1(new_n745), .B2(new_n480), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n742), .B1(new_n746), .B2(G29), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT87), .B(G2067), .Z(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n740), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g325(.A1(new_n726), .A2(new_n733), .A3(new_n735), .A4(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(G29), .A2(G35), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G162), .B2(G29), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT92), .B(KEYINPUT29), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n755), .A2(G2090), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT93), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n481), .A2(G139), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT88), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n467), .A2(new_n468), .ZN(new_n760));
  AOI22_X1  g335(.A1(new_n760), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n761));
  INV_X1    g336(.A(new_n465), .ZN(new_n762));
  AOI21_X1  g337(.A(KEYINPUT25), .B1(new_n762), .B2(G103), .ZN(new_n763));
  AND3_X1   g338(.A1(new_n762), .A2(KEYINPUT25), .A3(G103), .ZN(new_n764));
  OAI221_X1 g339(.A(new_n759), .B1(new_n460), .B2(new_n761), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  MUX2_X1   g340(.A(G33), .B(new_n765), .S(G29), .Z(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(G2072), .Z(new_n767));
  NAND2_X1  g342(.A1(new_n716), .A2(G20), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT23), .Z(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G299), .B2(G16), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G1956), .ZN(new_n771));
  NAND3_X1  g346(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT26), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n772), .A2(new_n773), .ZN(new_n775));
  AOI22_X1  g350(.A1(new_n774), .A2(new_n775), .B1(G105), .B2(new_n762), .ZN(new_n776));
  INV_X1    g351(.A(G141), .ZN(new_n777));
  INV_X1    g352(.A(G129), .ZN(new_n778));
  OAI221_X1 g353(.A(new_n776), .B1(new_n480), .B2(new_n777), .C1(new_n778), .C2(new_n478), .ZN(new_n779));
  MUX2_X1   g354(.A(G32), .B(new_n779), .S(G29), .Z(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT90), .Z(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT27), .B(G1996), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  AOI22_X1  g358(.A1(new_n781), .A2(new_n782), .B1(new_n755), .B2(G2090), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n767), .A2(new_n771), .A3(new_n783), .A4(new_n784), .ZN(new_n785));
  NOR3_X1   g360(.A1(new_n751), .A2(new_n757), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n716), .A2(G23), .ZN(new_n787));
  INV_X1    g362(.A(G288), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(new_n788), .B2(new_n716), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT33), .B(G1976), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(G6), .A2(G16), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n601), .B2(G16), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT32), .B(G1981), .Z(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n716), .A2(G22), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT85), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(G303), .B2(G16), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G1971), .ZN(new_n799));
  AND3_X1   g374(.A1(new_n791), .A2(new_n795), .A3(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n801), .A2(KEYINPUT34), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n612), .A2(G16), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G16), .B2(G24), .ZN(new_n804));
  INV_X1    g379(.A(G1986), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n804), .A2(new_n805), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n481), .A2(G131), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n479), .A2(G119), .ZN(new_n809));
  MUX2_X1   g384(.A(G95), .B(G107), .S(G2105), .Z(new_n810));
  NAND2_X1  g385(.A1(new_n810), .A2(G2104), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n808), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  MUX2_X1   g387(.A(G25), .B(new_n812), .S(G29), .Z(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT35), .B(G1991), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT84), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n813), .B(new_n815), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(KEYINPUT86), .B2(KEYINPUT36), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n802), .A2(new_n806), .A3(new_n807), .A4(new_n817), .ZN(new_n818));
  AND2_X1   g393(.A1(new_n801), .A2(KEYINPUT34), .ZN(new_n819));
  NOR2_X1   g394(.A1(KEYINPUT86), .A2(KEYINPUT36), .ZN(new_n820));
  OR3_X1    g395(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n820), .B1(new_n818), .B2(new_n819), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n786), .A2(new_n821), .A3(new_n822), .ZN(G150));
  INV_X1    g398(.A(G150), .ZN(G311));
  INV_X1    g399(.A(G67), .ZN(new_n825));
  INV_X1    g400(.A(G80), .ZN(new_n826));
  OAI22_X1  g401(.A1(new_n527), .A2(new_n825), .B1(new_n826), .B2(new_n509), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n507), .B1(new_n827), .B2(KEYINPUT94), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(KEYINPUT94), .B2(new_n827), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n541), .A2(G93), .B1(G55), .B2(new_n512), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(G860), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT37), .Z(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n543), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n544), .A2(new_n829), .A3(new_n830), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT38), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n624), .A2(new_n632), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  AND2_X1   g414(.A1(new_n839), .A2(KEYINPUT39), .ZN(new_n840));
  INV_X1    g415(.A(G860), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(new_n839), .B2(KEYINPUT39), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n833), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(KEYINPUT95), .Z(G145));
  XNOR2_X1  g419(.A(new_n642), .B(G160), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(G162), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n812), .B(new_n646), .ZN(new_n847));
  MUX2_X1   g422(.A(G106), .B(G118), .S(G2105), .Z(new_n848));
  AOI22_X1  g423(.A1(new_n479), .A2(G130), .B1(G2104), .B2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(G142), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n849), .B1(new_n850), .B2(new_n480), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n847), .B(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n746), .B(new_n501), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n852), .A2(new_n854), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n765), .B(new_n779), .ZN(new_n857));
  AND3_X1   g432(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n857), .B1(new_n855), .B2(new_n856), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n846), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(KEYINPUT96), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT96), .ZN(new_n862));
  OAI211_X1 g437(.A(new_n862), .B(new_n846), .C1(new_n858), .C2(new_n859), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  NOR3_X1   g439(.A1(new_n858), .A2(new_n859), .A3(new_n846), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n865), .A2(G37), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g443(.A1(new_n831), .A2(G868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT41), .ZN(new_n870));
  AND3_X1   g445(.A1(new_n561), .A2(new_n570), .A3(new_n624), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n629), .A2(new_n624), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT98), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OR3_X1    g450(.A1(new_n629), .A2(KEYINPUT97), .A3(new_n624), .ZN(new_n876));
  OAI21_X1  g451(.A(KEYINPUT97), .B1(new_n629), .B2(new_n624), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n629), .A2(new_n624), .ZN(new_n878));
  NAND4_X1  g453(.A1(new_n876), .A2(new_n877), .A3(KEYINPUT41), .A4(new_n878), .ZN(new_n879));
  OAI211_X1 g454(.A(KEYINPUT98), .B(new_n870), .C1(new_n871), .C2(new_n872), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n875), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n836), .B(new_n635), .ZN(new_n882));
  OR2_X1    g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AND2_X1   g458(.A1(new_n877), .A2(new_n878), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(new_n876), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(new_n882), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT42), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n883), .A2(KEYINPUT42), .A3(new_n887), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n788), .B1(new_n610), .B2(new_n611), .ZN(new_n893));
  INV_X1    g468(.A(new_n611), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n894), .A2(G288), .A3(new_n609), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(G166), .B(KEYINPUT99), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(new_n601), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(KEYINPUT100), .B1(new_n896), .B2(new_n898), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n896), .A2(KEYINPUT100), .A3(new_n898), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n899), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(KEYINPUT101), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n892), .A2(new_n904), .ZN(new_n905));
  NAND4_X1  g480(.A1(new_n890), .A2(KEYINPUT101), .A3(new_n903), .A4(new_n891), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n869), .B1(new_n907), .B2(G868), .ZN(G295));
  AOI21_X1  g483(.A(new_n869), .B1(new_n907), .B2(G868), .ZN(G331));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n910));
  NAND2_X1  g485(.A1(G171), .A2(KEYINPUT102), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT102), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n912), .B1(new_n534), .B2(new_n537), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n911), .A2(G168), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(G301), .A2(G286), .A3(new_n912), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n914), .A2(new_n834), .A3(new_n835), .A4(new_n915), .ZN(new_n916));
  OR2_X1    g491(.A1(new_n916), .A2(KEYINPUT103), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(KEYINPUT103), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n914), .A2(new_n915), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(new_n836), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n917), .A2(new_n918), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n881), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n920), .A2(new_n916), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n923), .B1(new_n884), .B2(new_n876), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(KEYINPUT104), .B1(new_n922), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT104), .ZN(new_n927));
  AOI211_X1 g502(.A(new_n927), .B(new_n924), .C1(new_n881), .C2(new_n921), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n903), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT43), .ZN(new_n930));
  INV_X1    g505(.A(new_n902), .ZN(new_n931));
  OAI22_X1  g506(.A1(new_n931), .A2(new_n900), .B1(new_n898), .B2(new_n896), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n924), .B1(new_n881), .B2(new_n921), .ZN(new_n933));
  AOI21_X1  g508(.A(G37), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n929), .A2(new_n930), .A3(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT41), .B1(new_n871), .B2(new_n872), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(new_n923), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n886), .B1(new_n921), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n937), .A2(new_n870), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n903), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n934), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(KEYINPUT43), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n910), .B1(new_n935), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n929), .A2(KEYINPUT43), .A3(new_n934), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n941), .A2(new_n930), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT44), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n943), .A2(new_n946), .ZN(G397));
  XOR2_X1   g522(.A(new_n746), .B(G2067), .Z(new_n948));
  INV_X1    g523(.A(G1996), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n779), .B(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  OR2_X1    g526(.A1(new_n812), .A2(new_n815), .ZN(new_n952));
  OAI22_X1  g527(.A1(new_n951), .A2(new_n952), .B1(G2067), .B2(new_n746), .ZN(new_n953));
  INV_X1    g528(.A(G1384), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n501), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT45), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(G160), .A2(G40), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n953), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n948), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n959), .B1(new_n961), .B2(new_n779), .ZN(new_n962));
  NAND2_X1  g537(.A1(KEYINPUT124), .A2(KEYINPUT46), .ZN(new_n963));
  INV_X1    g538(.A(new_n959), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n949), .B1(KEYINPUT124), .B2(KEYINPUT46), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n963), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n959), .A2(KEYINPUT124), .A3(KEYINPUT46), .A4(new_n949), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n962), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  XNOR2_X1  g543(.A(KEYINPUT125), .B(KEYINPUT47), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n968), .B(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n612), .A2(new_n805), .A3(new_n959), .ZN(new_n971));
  XOR2_X1   g546(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n972));
  XNOR2_X1  g547(.A(new_n971), .B(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n812), .A2(new_n815), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n948), .A2(new_n950), .A3(new_n974), .A4(new_n952), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(new_n959), .ZN(new_n976));
  XOR2_X1   g551(.A(new_n976), .B(KEYINPUT126), .Z(new_n977));
  AOI211_X1 g552(.A(new_n960), .B(new_n970), .C1(new_n973), .C2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(G1981), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n595), .A2(new_n979), .A3(new_n600), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n541), .A2(G86), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n595), .A2(new_n981), .ZN(new_n982));
  OAI211_X1 g557(.A(KEYINPUT49), .B(new_n980), .C1(new_n982), .C2(new_n979), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT49), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n595), .A2(new_n979), .A3(new_n600), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n979), .B1(new_n595), .B2(new_n981), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n984), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G8), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n461), .A2(new_n462), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n495), .B1(new_n989), .B2(new_n493), .ZN(new_n990));
  AOI22_X1  g565(.A1(new_n990), .A2(G2105), .B1(new_n499), .B2(new_n498), .ZN(new_n991));
  AOI21_X1  g566(.A(G1384), .B1(new_n991), .B2(new_n492), .ZN(new_n992));
  INV_X1    g567(.A(G40), .ZN(new_n993));
  NOR3_X1   g568(.A1(new_n466), .A2(new_n471), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n988), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n983), .A2(new_n987), .A3(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G1976), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n996), .A2(new_n997), .A3(new_n788), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(new_n980), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT112), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT112), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n998), .A2(new_n1001), .A3(new_n980), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1000), .A2(new_n995), .A3(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g578(.A(KEYINPUT109), .B(G1976), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1004), .B1(new_n581), .B2(new_n586), .ZN(new_n1005));
  OAI21_X1  g580(.A(KEYINPUT110), .B1(new_n1005), .B2(KEYINPUT52), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1004), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n583), .A2(new_n585), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n541), .A2(G87), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n580), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1011), .A2(new_n578), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1007), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT110), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n581), .A2(new_n586), .A3(G1976), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1006), .A2(new_n1016), .A3(new_n995), .A4(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n994), .A2(new_n954), .A3(new_n501), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1019), .A2(new_n1017), .A3(G8), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT108), .ZN(new_n1021));
  AND3_X1   g596(.A1(new_n1020), .A2(new_n1021), .A3(KEYINPUT52), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1021), .B1(new_n1020), .B2(KEYINPUT52), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n996), .B(new_n1018), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g599(.A(new_n1024), .B(KEYINPUT111), .ZN(new_n1025));
  OAI211_X1 g600(.A(KEYINPUT55), .B(G8), .C1(new_n508), .C2(new_n520), .ZN(new_n1026));
  OR2_X1    g601(.A1(new_n1026), .A2(KEYINPUT106), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1026), .ZN(new_n1028));
  OAI21_X1  g603(.A(G8), .B1(new_n508), .B2(new_n520), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT106), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1027), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n958), .B1(new_n955), .B2(new_n956), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n501), .A2(KEYINPUT45), .A3(new_n954), .ZN(new_n1034));
  AOI21_X1  g609(.A(G1971), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT105), .B(KEYINPUT50), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n501), .A2(new_n954), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(new_n994), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT50), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1039), .B1(new_n501), .B2(new_n954), .ZN(new_n1040));
  NOR3_X1   g615(.A1(new_n1038), .A2(G2090), .A3(new_n1040), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1032), .B(G8), .C1(new_n1035), .C2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT107), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n501), .A2(KEYINPUT45), .A3(new_n954), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT45), .B1(new_n501), .B2(new_n954), .ZN(new_n1045));
  NOR3_X1   g620(.A1(new_n1044), .A2(new_n1045), .A3(new_n958), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n955), .A2(KEYINPUT50), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1047), .A2(new_n994), .A3(new_n1037), .ZN(new_n1048));
  OAI22_X1  g623(.A1(new_n1046), .A2(G1971), .B1(new_n1048), .B2(G2090), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT107), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1049), .A2(new_n1050), .A3(G8), .A4(new_n1032), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1043), .A2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1003), .B1(new_n1025), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1025), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1032), .B1(new_n1049), .B2(G8), .ZN(new_n1055));
  INV_X1    g630(.A(G2084), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1047), .A2(new_n1056), .A3(new_n994), .A4(new_n1037), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1057), .B1(new_n1046), .B2(G1966), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(G8), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT63), .ZN(new_n1060));
  NOR4_X1   g635(.A1(new_n1055), .A2(new_n1059), .A3(new_n1060), .A4(G286), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1054), .A2(new_n1061), .ZN(new_n1062));
  OAI211_X1 g637(.A(KEYINPUT113), .B(new_n994), .C1(new_n992), .C2(new_n1036), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT113), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1036), .B1(new_n501), .B2(new_n954), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1064), .B1(new_n1065), .B2(new_n958), .ZN(new_n1066));
  INV_X1    g641(.A(G2090), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n992), .A2(new_n1039), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1063), .A2(new_n1066), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1070));
  INV_X1    g645(.A(G1971), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1069), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(G8), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1032), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1024), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1059), .A2(G286), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1076), .A2(new_n1052), .A3(new_n1077), .ZN(new_n1078));
  XNOR2_X1  g653(.A(KEYINPUT114), .B(KEYINPUT63), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1053), .B1(new_n1062), .B2(new_n1080), .ZN(new_n1081));
  OAI211_X1 g656(.A(KEYINPUT51), .B(G8), .C1(new_n1058), .C2(G286), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT121), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n994), .B1(new_n992), .B2(KEYINPUT45), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n738), .B1(new_n1085), .B2(new_n1044), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n988), .B1(new_n1086), .B2(new_n1057), .ZN(new_n1087));
  NOR2_X1   g662(.A1(G168), .A2(new_n988), .ZN(new_n1088));
  OAI211_X1 g663(.A(KEYINPUT121), .B(KEYINPUT51), .C1(new_n1087), .C2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT51), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1088), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1059), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1084), .A2(new_n1089), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1087), .A2(G286), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1093), .A2(KEYINPUT62), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(KEYINPUT62), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1076), .A2(new_n1052), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT122), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1076), .A2(new_n1052), .A3(KEYINPUT122), .ZN(new_n1101));
  INV_X1    g676(.A(G2078), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n957), .A2(new_n1102), .A3(new_n1034), .A4(new_n994), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT53), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1033), .A2(KEYINPUT53), .A3(new_n1102), .A4(new_n1034), .ZN(new_n1106));
  INV_X1    g681(.A(G1961), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1048), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1105), .A2(new_n1106), .A3(new_n1108), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1100), .A2(G171), .A3(new_n1101), .A4(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1081), .B1(new_n1097), .B2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1063), .A2(new_n1066), .A3(new_n1068), .ZN(new_n1112));
  XNOR2_X1  g687(.A(KEYINPUT115), .B(G1956), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1113), .ZN(new_n1114));
  AND2_X1   g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT57), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n629), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  XOR2_X1   g694(.A(KEYINPUT56), .B(G2072), .Z(new_n1120));
  NOR2_X1   g695(.A1(new_n1070), .A2(new_n1120), .ZN(new_n1121));
  NOR3_X1   g696(.A1(new_n1115), .A2(new_n1119), .A3(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g697(.A(new_n1122), .B(KEYINPUT61), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1033), .A2(new_n949), .A3(new_n1034), .ZN(new_n1125));
  XOR2_X1   g700(.A(KEYINPUT58), .B(G1341), .Z(new_n1126));
  NAND2_X1  g701(.A1(new_n1019), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT118), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1019), .A2(KEYINPUT118), .A3(new_n1126), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1125), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(new_n544), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1124), .B1(new_n1132), .B2(KEYINPUT120), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1019), .A2(G2067), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1134), .B1(new_n1048), .B2(new_n730), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n624), .B1(new_n1135), .B2(KEYINPUT60), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1136), .B1(KEYINPUT60), .B2(new_n1135), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1119), .B1(new_n1115), .B2(new_n1121), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1133), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1132), .A2(KEYINPUT119), .ZN(new_n1140));
  NOR3_X1   g715(.A1(new_n1124), .A2(KEYINPUT119), .A3(KEYINPUT120), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1131), .A2(new_n544), .A3(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1135), .A2(KEYINPUT60), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1140), .B(new_n1142), .C1(new_n625), .C2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1139), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1121), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT116), .ZN(new_n1148));
  AND3_X1   g723(.A1(new_n1146), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1148), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT117), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1119), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(KEYINPUT117), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1153));
  OAI22_X1  g728(.A1(new_n1149), .A2(new_n1150), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1155), .A2(G1348), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n625), .B1(new_n1156), .B2(new_n1134), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1154), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1122), .ZN(new_n1159));
  AOI22_X1  g734(.A1(new_n1123), .A2(new_n1145), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1109), .A2(G171), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1105), .A2(new_n1108), .A3(G301), .A4(new_n1106), .ZN(new_n1163));
  AND3_X1   g738(.A1(new_n1162), .A2(KEYINPUT54), .A3(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(KEYINPUT54), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  AND4_X1   g741(.A1(new_n1100), .A2(new_n1161), .A3(new_n1101), .A4(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1160), .B1(new_n1167), .B2(KEYINPUT123), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1100), .A2(new_n1161), .A3(new_n1101), .A4(new_n1166), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT123), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1111), .B1(new_n1168), .B2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n975), .B1(new_n805), .B2(new_n612), .ZN(new_n1173));
  NAND2_X1  g748(.A1(G290), .A2(G1986), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n964), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n978), .B1(new_n1172), .B2(new_n1175), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g751(.A(G319), .ZN(new_n1178));
  NOR3_X1   g752(.A1(G229), .A2(G227), .A3(new_n1178), .ZN(new_n1179));
  NAND2_X1  g753(.A1(new_n670), .A2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g754(.A(new_n1180), .B1(new_n864), .B2(new_n866), .ZN(new_n1181));
  AND3_X1   g755(.A1(new_n1181), .A2(new_n945), .A3(new_n944), .ZN(G308));
  NAND3_X1  g756(.A1(new_n1181), .A2(new_n945), .A3(new_n944), .ZN(G225));
endmodule


