//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 0 0 0 1 1 1 0 1 1 1 0 0 1 0 0 1 1 1 0 1 0 0 0 0 0 0 0 0 1 0 1 1 0 0 1 1 0 0 0 0 1 0 0 1 1 0 0 1 0 0 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:00 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(G137), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n188), .A2(KEYINPUT11), .A3(G134), .ZN(new_n189));
  INV_X1    g003(.A(G134), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G137), .ZN(new_n191));
  AOI21_X1  g005(.A(KEYINPUT11), .B1(new_n188), .B2(G134), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT66), .ZN(new_n193));
  OAI211_X1 g007(.A(new_n189), .B(new_n191), .C1(new_n192), .C2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT11), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n195), .B1(new_n190), .B2(G137), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(KEYINPUT66), .ZN(new_n197));
  OAI21_X1  g011(.A(G131), .B1(new_n194), .B2(new_n197), .ZN(new_n198));
  AND2_X1   g012(.A1(new_n189), .A2(new_n191), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n192), .A2(new_n193), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n196), .A2(KEYINPUT66), .ZN(new_n201));
  INV_X1    g015(.A(G131), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n199), .A2(new_n200), .A3(new_n201), .A4(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n198), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT69), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT64), .B1(new_n207), .B2(G146), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT64), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(new_n210), .A3(G143), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n207), .A2(G146), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n208), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(KEYINPUT0), .A2(G128), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(KEYINPUT0), .A2(G128), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n213), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT65), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n213), .A2(KEYINPUT65), .A3(new_n217), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n207), .A2(G146), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(new_n212), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  AOI22_X1  g039(.A1(new_n220), .A2(new_n221), .B1(new_n215), .B2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n198), .A2(KEYINPUT69), .A3(new_n203), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n206), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT1), .ZN(new_n229));
  OAI21_X1  g043(.A(G128), .B1(new_n222), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n213), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT67), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT67), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n213), .A2(new_n230), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G128), .ZN(new_n236));
  NOR3_X1   g050(.A1(new_n224), .A2(KEYINPUT1), .A3(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n191), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n190), .A2(G137), .ZN(new_n241));
  OAI21_X1  g055(.A(G131), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n203), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n239), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G119), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G116), .ZN(new_n247));
  INV_X1    g061(.A(G116), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G119), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n250), .A2(KEYINPUT68), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT2), .B(G113), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n251), .B(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n228), .A2(new_n245), .A3(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT28), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n254), .ZN(new_n259));
  INV_X1    g073(.A(new_n204), .ZN(new_n260));
  AND3_X1   g074(.A1(new_n213), .A2(KEYINPUT65), .A3(new_n217), .ZN(new_n261));
  AOI21_X1  g075(.A(KEYINPUT65), .B1(new_n213), .B2(new_n217), .ZN(new_n262));
  OAI22_X1  g076(.A1(new_n261), .A2(new_n262), .B1(new_n214), .B2(new_n224), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n243), .B1(new_n235), .B2(new_n238), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n259), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n266), .B1(new_n255), .B2(new_n256), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n258), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G237), .ZN(new_n269));
  INV_X1    g083(.A(G953), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n269), .A2(new_n270), .A3(G210), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n271), .B(KEYINPUT27), .ZN(new_n272));
  XNOR2_X1  g086(.A(KEYINPUT26), .B(G101), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n272), .B(new_n273), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n274), .B(KEYINPUT70), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT29), .B1(new_n268), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n228), .A2(new_n245), .A3(KEYINPUT30), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT30), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n279), .B1(new_n264), .B2(new_n265), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n278), .A2(new_n280), .A3(new_n259), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n255), .ZN(new_n282));
  INV_X1    g096(.A(new_n274), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(G902), .B1(new_n277), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n228), .A2(new_n245), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n259), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n287), .A2(KEYINPUT73), .A3(new_n255), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT73), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n286), .A2(new_n289), .A3(new_n259), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n288), .A2(KEYINPUT28), .A3(new_n290), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n291), .A2(KEYINPUT29), .A3(new_n274), .A4(new_n257), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n187), .B1(new_n285), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT32), .ZN(new_n294));
  NOR2_X1   g108(.A1(G472), .A2(G902), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT71), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n297), .B(new_n275), .C1(new_n258), .C2(new_n267), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  AND3_X1   g113(.A1(new_n198), .A2(KEYINPUT69), .A3(new_n203), .ZN(new_n300));
  AOI21_X1  g114(.A(KEYINPUT69), .B1(new_n198), .B2(new_n203), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n265), .B1(new_n302), .B2(new_n226), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n303), .A2(KEYINPUT28), .A3(new_n254), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n304), .A2(new_n257), .A3(new_n266), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n297), .B1(new_n305), .B2(new_n275), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n299), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n281), .A2(new_n255), .A3(new_n274), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT31), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n281), .A2(KEYINPUT31), .A3(new_n255), .A4(new_n274), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n296), .B1(new_n307), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n294), .B1(new_n313), .B2(KEYINPUT72), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT71), .B1(new_n268), .B2(new_n276), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n312), .A2(new_n315), .A3(new_n298), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n295), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT72), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(new_n318), .A3(KEYINPUT32), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n293), .B1(new_n314), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G217), .ZN(new_n321));
  INV_X1    g135(.A(G902), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n321), .B1(G234), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(KEYINPUT22), .B(G137), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n270), .A2(G221), .A3(G234), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n325), .B(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G140), .ZN(new_n328));
  NOR2_X1   g142(.A1(KEYINPUT74), .A2(G125), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(KEYINPUT74), .A2(G125), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n328), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NOR2_X1   g146(.A1(G125), .A2(G140), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT16), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n330), .A2(new_n331), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT16), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n335), .A2(new_n336), .A3(new_n328), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n334), .A2(G146), .A3(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n331), .ZN(new_n339));
  OAI21_X1  g153(.A(G140), .B1(new_n339), .B2(new_n329), .ZN(new_n340));
  INV_X1    g154(.A(new_n333), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n336), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  AOI211_X1 g156(.A(KEYINPUT16), .B(G140), .C1(new_n330), .C2(new_n331), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n210), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n338), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT23), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n346), .B1(new_n246), .B2(G128), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n236), .A2(KEYINPUT23), .A3(G119), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n347), .B(new_n348), .C1(G119), .C2(new_n236), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(G110), .ZN(new_n350));
  XOR2_X1   g164(.A(KEYINPUT24), .B(G110), .Z(new_n351));
  XNOR2_X1  g165(.A(G119), .B(G128), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n345), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(KEYINPUT75), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT75), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n345), .A2(new_n358), .A3(new_n355), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  XNOR2_X1  g174(.A(G125), .B(G140), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n210), .ZN(new_n362));
  XOR2_X1   g176(.A(KEYINPUT76), .B(G110), .Z(new_n363));
  OAI22_X1  g177(.A1(new_n349), .A2(new_n363), .B1(new_n352), .B2(new_n351), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n338), .A2(new_n362), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(KEYINPUT77), .B1(new_n360), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n358), .B1(new_n345), .B2(new_n355), .ZN(new_n367));
  AOI211_X1 g181(.A(KEYINPUT75), .B(new_n354), .C1(new_n338), .C2(new_n344), .ZN(new_n368));
  OAI211_X1 g182(.A(KEYINPUT77), .B(new_n365), .C1(new_n367), .C2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n327), .B1(new_n366), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n327), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n371), .A2(new_n322), .A3(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT25), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n365), .B1(new_n367), .B2(new_n368), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT77), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n372), .B1(new_n379), .B2(new_n369), .ZN(new_n380));
  INV_X1    g194(.A(new_n373), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(KEYINPUT25), .A3(new_n322), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n324), .B1(new_n376), .B2(new_n383), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n323), .A2(G902), .ZN(new_n385));
  AND2_X1   g199(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n320), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(G214), .B1(G237), .B2(G902), .ZN(new_n390));
  XOR2_X1   g204(.A(new_n390), .B(KEYINPUT85), .Z(new_n391));
  NAND2_X1  g205(.A1(G234), .A2(G237), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(G952), .A3(new_n270), .ZN(new_n393));
  XNOR2_X1  g207(.A(KEYINPUT21), .B(G898), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n392), .A2(G902), .A3(G953), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n393), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(G210), .B1(G237), .B2(G902), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT6), .ZN(new_n401));
  INV_X1    g215(.A(G104), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(KEYINPUT81), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT81), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G104), .ZN(new_n405));
  AOI21_X1  g219(.A(G107), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(G107), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n407), .A2(G104), .ZN(new_n408));
  OAI21_X1  g222(.A(G101), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n250), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(KEYINPUT5), .ZN(new_n411));
  OAI21_X1  g225(.A(G113), .B1(new_n247), .B2(KEYINPUT5), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  AOI22_X1  g227(.A1(new_n411), .A2(new_n413), .B1(new_n410), .B2(new_n253), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT3), .ZN(new_n415));
  OAI21_X1  g229(.A(KEYINPUT82), .B1(new_n406), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT82), .ZN(new_n417));
  XNOR2_X1  g231(.A(KEYINPUT81), .B(G104), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n417), .B(KEYINPUT3), .C1(new_n418), .C2(G107), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  NOR3_X1   g234(.A1(new_n402), .A2(KEYINPUT3), .A3(G107), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(G101), .B1(new_n418), .B2(G107), .ZN(new_n423));
  AND4_X1   g237(.A1(KEYINPUT83), .A2(new_n420), .A3(new_n422), .A4(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n421), .B1(new_n416), .B2(new_n419), .ZN(new_n425));
  AOI21_X1  g239(.A(KEYINPUT83), .B1(new_n425), .B2(new_n423), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n409), .B(new_n414), .C1(new_n424), .C2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT86), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n420), .A2(new_n422), .A3(new_n423), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT83), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n425), .A2(KEYINPUT83), .A3(new_n423), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT86), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n433), .A2(new_n434), .A3(new_n409), .A4(new_n414), .ZN(new_n435));
  INV_X1    g249(.A(G101), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n418), .A2(G107), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n436), .B1(new_n425), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT4), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n433), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n254), .B1(new_n438), .B2(new_n439), .ZN(new_n442));
  AOI22_X1  g256(.A1(new_n428), .A2(new_n435), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(G110), .B(G122), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n401), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n441), .A2(new_n442), .ZN(new_n446));
  INV_X1    g260(.A(new_n409), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n447), .B1(new_n431), .B2(new_n432), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n434), .B1(new_n448), .B2(new_n414), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n427), .A2(KEYINPUT86), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n446), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n444), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n445), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n235), .A2(new_n238), .A3(new_n330), .A4(new_n331), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n263), .A2(new_n335), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n270), .A2(G224), .ZN(new_n458));
  XOR2_X1   g272(.A(new_n458), .B(KEYINPUT87), .Z(new_n459));
  XNOR2_X1  g273(.A(new_n457), .B(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n451), .A2(new_n401), .A3(new_n452), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n454), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n444), .B(new_n446), .C1(new_n449), .C2(new_n450), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT92), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n458), .A2(KEYINPUT7), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n464), .B1(new_n457), .B2(new_n465), .ZN(new_n466));
  OR3_X1    g280(.A1(new_n457), .A2(new_n464), .A3(new_n465), .ZN(new_n467));
  OR2_X1    g281(.A1(new_n455), .A2(KEYINPUT91), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n455), .A2(KEYINPUT91), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(new_n456), .A3(new_n469), .ZN(new_n470));
  AOI22_X1  g284(.A1(new_n466), .A2(new_n467), .B1(new_n470), .B2(new_n465), .ZN(new_n471));
  XOR2_X1   g285(.A(new_n444), .B(KEYINPUT8), .Z(new_n472));
  OAI21_X1  g286(.A(new_n409), .B1(new_n424), .B2(new_n426), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n472), .B1(new_n473), .B2(new_n414), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n413), .A2(KEYINPUT88), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT88), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n412), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n475), .A2(new_n411), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n410), .A2(new_n253), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n480), .B(KEYINPUT89), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n448), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n474), .A2(KEYINPUT90), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(KEYINPUT90), .B1(new_n474), .B2(new_n482), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n463), .B(new_n471), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n485), .A2(KEYINPUT93), .A3(new_n322), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n462), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(KEYINPUT93), .B1(new_n485), .B2(new_n322), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n400), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n485), .A2(new_n322), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT93), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n492), .A2(new_n399), .A3(new_n462), .A4(new_n486), .ZN(new_n493));
  AOI211_X1 g307(.A(new_n391), .B(new_n398), .C1(new_n489), .C2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(G469), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n270), .A2(G227), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n496), .B(KEYINPUT80), .ZN(new_n497));
  XNOR2_X1  g311(.A(G110), .B(G140), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n497), .B(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n263), .B1(new_n438), .B2(new_n439), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n237), .B1(new_n232), .B2(new_n234), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT10), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI22_X1  g318(.A1(new_n441), .A2(new_n501), .B1(new_n448), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n237), .B1(new_n224), .B2(new_n230), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n409), .B(new_n507), .C1(new_n424), .C2(new_n426), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n508), .A2(KEYINPUT84), .A3(new_n503), .ZN(new_n509));
  AOI21_X1  g323(.A(KEYINPUT84), .B1(new_n508), .B2(new_n503), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n505), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n302), .ZN(new_n512));
  INV_X1    g326(.A(new_n302), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n505), .B(new_n513), .C1(new_n509), .C2(new_n510), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n500), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  AND2_X1   g329(.A1(new_n204), .A2(KEYINPUT12), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n448), .A2(new_n239), .ZN(new_n517));
  INV_X1    g331(.A(new_n508), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n473), .A2(new_n502), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n513), .B1(new_n520), .B2(new_n508), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n519), .B1(new_n521), .B2(KEYINPUT12), .ZN(new_n522));
  AND3_X1   g336(.A1(new_n522), .A2(new_n514), .A3(new_n500), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n495), .B(new_n322), .C1(new_n515), .C2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(G469), .A2(G902), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n522), .A2(new_n514), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n499), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n512), .A2(new_n514), .A3(new_n500), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n527), .A2(G469), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n524), .A2(new_n525), .A3(new_n529), .ZN(new_n530));
  XOR2_X1   g344(.A(KEYINPUT9), .B(G234), .Z(new_n531));
  XNOR2_X1  g345(.A(new_n531), .B(KEYINPUT78), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(new_n322), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(G221), .ZN(new_n534));
  XOR2_X1   g348(.A(new_n534), .B(KEYINPUT79), .Z(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n530), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n236), .A2(G143), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n207), .A2(G128), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n540), .B(new_n190), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n248), .A2(KEYINPUT14), .A3(G122), .ZN(new_n542));
  XNOR2_X1  g356(.A(G116), .B(G122), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  OAI211_X1 g358(.A(G107), .B(new_n542), .C1(new_n544), .C2(KEYINPUT14), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n543), .A2(new_n407), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n541), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  OR2_X1    g361(.A1(new_n547), .A2(KEYINPUT96), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n543), .B(new_n407), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n540), .A2(new_n190), .ZN(new_n550));
  AND2_X1   g364(.A1(new_n538), .A2(KEYINPUT13), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n538), .A2(KEYINPUT13), .ZN(new_n552));
  NOR3_X1   g366(.A1(new_n551), .A2(new_n552), .A3(new_n539), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n549), .B(new_n550), .C1(new_n553), .C2(new_n190), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n547), .A2(KEYINPUT96), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n548), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n532), .A2(G217), .A3(new_n270), .ZN(new_n557));
  OR2_X1    g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n557), .ZN(new_n559));
  AOI21_X1  g373(.A(G902), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT97), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI211_X1 g376(.A(KEYINPUT97), .B(G902), .C1(new_n558), .C2(new_n559), .ZN(new_n563));
  INV_X1    g377(.A(G478), .ZN(new_n564));
  OAI22_X1  g378(.A1(new_n562), .A2(new_n563), .B1(KEYINPUT15), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n269), .A2(new_n270), .A3(G214), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(new_n207), .ZN(new_n567));
  NAND2_X1  g381(.A1(KEYINPUT18), .A2(G131), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n567), .B(new_n568), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n332), .A2(new_n333), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n362), .B1(new_n571), .B2(new_n210), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n567), .A2(KEYINPUT17), .A3(G131), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n567), .B(G131), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n574), .B1(new_n575), .B2(KEYINPUT17), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n573), .B1(new_n576), .B2(new_n345), .ZN(new_n577));
  XNOR2_X1  g391(.A(G113), .B(G122), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n578), .B(new_n402), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT19), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n361), .A2(new_n581), .ZN(new_n582));
  OR2_X1    g396(.A1(new_n582), .A2(KEYINPUT94), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(KEYINPUT94), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n583), .B(new_n584), .C1(new_n571), .C2(new_n581), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n338), .B(new_n575), .C1(new_n585), .C2(G146), .ZN(new_n586));
  INV_X1    g400(.A(new_n579), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n586), .A2(new_n587), .A3(new_n573), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n580), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(G475), .A2(G902), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  OR3_X1    g405(.A1(new_n589), .A2(KEYINPUT20), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(KEYINPUT20), .B1(new_n589), .B2(new_n591), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n560), .A2(new_n561), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT15), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n595), .A2(new_n596), .A3(G478), .ZN(new_n597));
  OR2_X1    g411(.A1(new_n579), .A2(KEYINPUT95), .ZN(new_n598));
  OR2_X1    g412(.A1(new_n577), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n577), .A2(new_n598), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n599), .A2(new_n322), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(G475), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n565), .A2(new_n594), .A3(new_n597), .A4(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n537), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n389), .A2(new_n494), .A3(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(G101), .ZN(G3));
  NAND3_X1  g420(.A1(new_n530), .A2(new_n387), .A3(new_n536), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n187), .B1(new_n316), .B2(new_n322), .ZN(new_n608));
  OAI21_X1  g422(.A(KEYINPUT98), .B1(new_n608), .B2(new_n313), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT98), .ZN(new_n610));
  AOI21_X1  g424(.A(G902), .B1(new_n307), .B2(new_n312), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n610), .B1(new_n611), .B2(new_n187), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n607), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g428(.A(new_n614), .B(KEYINPUT99), .Z(new_n615));
  NAND2_X1  g429(.A1(new_n489), .A2(new_n493), .ZN(new_n616));
  INV_X1    g430(.A(new_n391), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT100), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n616), .A2(KEYINPUT100), .A3(new_n617), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n560), .A2(new_n564), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n564), .A2(new_n322), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n558), .A2(new_n559), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT33), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n626), .B1(new_n629), .B2(G478), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n594), .A2(new_n602), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n632), .A2(new_n398), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n615), .A2(new_n622), .A3(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT34), .B(G104), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G6));
  NAND2_X1  g450(.A1(new_n565), .A2(new_n597), .ZN(new_n637));
  INV_X1    g451(.A(new_n631), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n639), .A2(new_n398), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n615), .A2(new_n622), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT35), .B(G107), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G9));
  NOR2_X1   g457(.A1(new_n374), .A2(new_n375), .ZN(new_n644));
  AOI21_X1  g458(.A(KEYINPUT25), .B1(new_n382), .B2(new_n322), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n323), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n372), .A2(KEYINPUT36), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n377), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n385), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n609), .A2(new_n612), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(KEYINPUT101), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT101), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n609), .A2(new_n650), .A3(new_n653), .A4(new_n612), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n652), .A2(new_n494), .A3(new_n604), .A4(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT37), .B(G110), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G12));
  INV_X1    g471(.A(new_n293), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n313), .A2(KEYINPUT72), .A3(new_n294), .ZN(new_n659));
  AOI21_X1  g473(.A(KEYINPUT32), .B1(new_n317), .B2(new_n318), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n514), .A2(new_n500), .ZN(new_n662));
  AOI22_X1  g476(.A1(new_n662), .A2(new_n512), .B1(new_n526), .B2(new_n499), .ZN(new_n663));
  OAI21_X1  g477(.A(G469), .B1(new_n663), .B2(G902), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n535), .B1(new_n664), .B2(new_n524), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n270), .A2(G900), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n392), .A2(G902), .ZN(new_n668));
  OR3_X1    g482(.A1(new_n667), .A2(KEYINPUT102), .A3(new_n668), .ZN(new_n669));
  OAI21_X1  g483(.A(KEYINPUT102), .B1(new_n667), .B2(new_n668), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n669), .A2(new_n393), .A3(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n639), .A2(new_n672), .ZN(new_n673));
  AND3_X1   g487(.A1(new_n661), .A2(new_n665), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g488(.A(KEYINPUT100), .B1(new_n616), .B2(new_n617), .ZN(new_n675));
  AOI211_X1 g489(.A(new_n619), .B(new_n391), .C1(new_n489), .C2(new_n493), .ZN(new_n676));
  OAI211_X1 g490(.A(new_n674), .B(new_n650), .C1(new_n675), .C2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G128), .ZN(G30));
  XNOR2_X1  g492(.A(new_n616), .B(KEYINPUT38), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n187), .A2(new_n322), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  AND3_X1   g495(.A1(new_n288), .A2(new_n275), .A3(new_n290), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n308), .A2(G472), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n681), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT103), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n686), .B1(new_n314), .B2(new_n319), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n637), .ZN(new_n689));
  NOR4_X1   g503(.A1(new_n650), .A2(new_n689), .A3(new_n391), .A4(new_n638), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n679), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  OR2_X1    g505(.A1(new_n691), .A2(KEYINPUT104), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(KEYINPUT104), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n671), .B(KEYINPUT39), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n665), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g509(.A(new_n695), .B(KEYINPUT40), .Z(new_n696));
  NAND3_X1  g510(.A1(new_n692), .A2(new_n693), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(KEYINPUT105), .B(G143), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G45));
  NAND3_X1  g513(.A1(new_n630), .A2(new_n631), .A3(new_n671), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n320), .A2(new_n537), .A3(new_n700), .ZN(new_n701));
  OAI211_X1 g515(.A(new_n701), .B(new_n650), .C1(new_n675), .C2(new_n676), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G146), .ZN(G48));
  OAI21_X1  g517(.A(new_n322), .B1(new_n515), .B2(new_n523), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(G469), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n705), .A2(new_n536), .A3(new_n524), .ZN(new_n706));
  NOR3_X1   g520(.A1(new_n320), .A2(new_n706), .A3(new_n388), .ZN(new_n707));
  OAI211_X1 g521(.A(new_n707), .B(new_n633), .C1(new_n675), .C2(new_n676), .ZN(new_n708));
  XNOR2_X1  g522(.A(KEYINPUT41), .B(G113), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G15));
  OAI211_X1 g524(.A(new_n707), .B(new_n640), .C1(new_n675), .C2(new_n676), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G116), .ZN(G18));
  INV_X1    g526(.A(new_n649), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n384), .A2(new_n713), .ZN(new_n714));
  NOR4_X1   g528(.A1(new_n320), .A2(new_n398), .A3(new_n603), .A4(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n706), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n717), .B1(new_n675), .B2(new_n676), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(KEYINPUT106), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT106), .ZN(new_n720));
  OAI211_X1 g534(.A(new_n720), .B(new_n717), .C1(new_n675), .C2(new_n676), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n716), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(new_n246), .ZN(G21));
  INV_X1    g537(.A(new_n312), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n276), .B1(new_n291), .B2(new_n257), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n295), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n316), .A2(new_n322), .ZN(new_n727));
  XOR2_X1   g541(.A(KEYINPUT107), .B(G472), .Z(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n387), .A2(new_n726), .A3(new_n729), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n730), .A2(new_n706), .A3(new_n398), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n689), .A2(new_n638), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n731), .B(new_n732), .C1(new_n675), .C2(new_n676), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G122), .ZN(G24));
  NAND2_X1  g548(.A1(new_n729), .A2(new_n726), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n700), .A2(new_n735), .A3(new_n714), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n720), .B1(new_n622), .B2(new_n717), .ZN(new_n737));
  INV_X1    g551(.A(new_n721), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G125), .ZN(G27));
  NAND3_X1  g554(.A1(new_n489), .A2(new_n617), .A3(new_n493), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n741), .A2(new_n537), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n700), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n658), .B1(KEYINPUT32), .B2(new_n313), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n317), .A2(new_n294), .ZN(new_n746));
  OAI211_X1 g560(.A(new_n744), .B(new_n387), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  OAI21_X1  g561(.A(KEYINPUT42), .B1(new_n743), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n700), .A2(KEYINPUT42), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n742), .A2(new_n661), .A3(new_n749), .A4(new_n387), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(new_n202), .ZN(G33));
  NAND4_X1  g566(.A1(new_n742), .A2(new_n661), .A3(new_n387), .A4(new_n673), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G134), .ZN(G36));
  OAI211_X1 g568(.A(new_n623), .B(new_n625), .C1(new_n628), .C2(new_n564), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT43), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT108), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n631), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n638), .A2(KEYINPUT108), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n757), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT109), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n761), .B(new_n762), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n756), .B1(new_n755), .B2(new_n631), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n765), .A2(KEYINPUT44), .A3(new_n613), .A4(new_n650), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(KEYINPUT110), .ZN(new_n767));
  OR2_X1    g581(.A1(new_n663), .A2(KEYINPUT45), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n663), .A2(KEYINPUT45), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n768), .A2(G469), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(KEYINPUT46), .B1(new_n770), .B2(new_n525), .ZN(new_n771));
  INV_X1    g585(.A(new_n524), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n770), .A2(KEYINPUT46), .A3(new_n525), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n535), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n775), .A2(new_n694), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n765), .A2(new_n613), .A3(new_n650), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT44), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n741), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n767), .A2(new_n776), .A3(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G137), .ZN(G39));
  XOR2_X1   g595(.A(new_n775), .B(KEYINPUT47), .Z(new_n782));
  AND3_X1   g596(.A1(new_n489), .A2(new_n617), .A3(new_n493), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n783), .A2(new_n320), .A3(new_n388), .A4(new_n744), .ZN(new_n784));
  OR2_X1    g598(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G140), .ZN(G42));
  INV_X1    g600(.A(new_n679), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n705), .A2(new_n524), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(KEYINPUT49), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n755), .A2(new_n391), .A3(new_n535), .ZN(new_n790));
  AND4_X1   g604(.A1(new_n387), .A2(new_n790), .A3(new_n759), .A4(new_n760), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n787), .A2(new_n687), .A3(new_n789), .A4(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n393), .B1(new_n763), .B2(new_n764), .ZN(new_n793));
  INV_X1    g607(.A(new_n730), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n795), .A2(new_n617), .A3(new_n706), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n787), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT50), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n796), .A2(KEYINPUT50), .A3(new_n787), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n741), .A2(new_n706), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n793), .A2(new_n802), .ZN(new_n803));
  XOR2_X1   g617(.A(new_n803), .B(KEYINPUT117), .Z(new_n804));
  NAND4_X1  g618(.A1(new_n804), .A2(new_n650), .A3(new_n726), .A4(new_n729), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n788), .A2(new_n535), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n782), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n795), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n807), .A2(new_n783), .A3(new_n808), .ZN(new_n809));
  OR3_X1    g623(.A1(new_n688), .A2(new_n388), .A3(new_n393), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n811), .A2(new_n638), .A3(new_n755), .A4(new_n802), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n801), .A2(new_n805), .A3(new_n809), .A4(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT51), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT118), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n815), .B(new_n816), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n387), .B1(new_n745), .B2(new_n746), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n804), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT48), .ZN(new_n821));
  OR3_X1    g635(.A1(new_n820), .A2(KEYINPUT120), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n820), .A2(new_n821), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(KEYINPUT119), .ZN(new_n824));
  OAI21_X1  g638(.A(KEYINPUT120), .B1(new_n820), .B2(new_n821), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT119), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n820), .A2(new_n826), .A3(new_n821), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n822), .A2(new_n824), .A3(new_n825), .A4(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(KEYINPUT116), .B(KEYINPUT51), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n813), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n795), .B1(new_n721), .B2(new_n719), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n811), .A2(new_n802), .ZN(new_n832));
  OAI211_X1 g646(.A(G952), .B(new_n270), .C1(new_n832), .C2(new_n632), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n828), .A2(new_n830), .A3(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n715), .B1(new_n737), .B2(new_n738), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n708), .A2(new_n711), .A3(new_n733), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n836), .A2(KEYINPUT115), .A3(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT115), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n708), .A2(new_n711), .A3(new_n733), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n839), .B1(new_n722), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n748), .A2(new_n750), .A3(new_n753), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n714), .A2(new_n603), .A3(new_n672), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n783), .A2(new_n661), .A3(new_n843), .A4(new_n665), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT112), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT112), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n742), .A2(new_n846), .A3(new_n661), .A4(new_n843), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n742), .A2(new_n736), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n845), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n639), .A2(KEYINPUT111), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT111), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n637), .A2(new_n638), .A3(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n850), .A2(new_n632), .A3(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n614), .A2(new_n494), .A3(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n655), .A2(new_n854), .A3(new_n605), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n842), .A2(new_n849), .A3(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n838), .A2(new_n841), .A3(KEYINPUT53), .A4(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n714), .A2(new_n671), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n687), .A2(new_n537), .A3(new_n859), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n860), .B(new_n732), .C1(new_n675), .C2(new_n676), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n677), .A2(new_n702), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(KEYINPUT113), .B1(new_n739), .B2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT52), .ZN(new_n864));
  INV_X1    g678(.A(new_n736), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n865), .B1(new_n719), .B2(new_n721), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n677), .A2(new_n702), .A3(new_n861), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n864), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n739), .A2(KEYINPUT52), .A3(new_n862), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n863), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n863), .A2(KEYINPUT52), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n858), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT54), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT114), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n869), .A2(new_n868), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n849), .A2(new_n855), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n748), .A2(new_n750), .A3(new_n753), .ZN(new_n878));
  AND4_X1   g692(.A1(new_n836), .A2(new_n877), .A3(new_n837), .A4(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT53), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n875), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI211_X1 g696(.A(KEYINPUT114), .B(KEYINPUT53), .C1(new_n876), .C2(new_n879), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n873), .B(new_n874), .C1(new_n882), .C2(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n870), .A2(new_n872), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n836), .A2(new_n877), .A3(new_n837), .A4(new_n878), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n886), .A2(KEYINPUT53), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n886), .B1(new_n868), .B2(new_n869), .ZN(new_n889));
  OAI22_X1  g703(.A1(new_n885), .A2(new_n888), .B1(new_n881), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n884), .B1(new_n890), .B2(new_n874), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n817), .A2(new_n835), .A3(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(G952), .A2(G953), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n792), .B1(new_n892), .B2(new_n893), .ZN(G75));
  AND2_X1   g708(.A1(new_n454), .A2(new_n461), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(new_n460), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT55), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT113), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n898), .B1(new_n866), .B2(new_n867), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT52), .B1(new_n739), .B2(new_n862), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n866), .A2(new_n867), .A3(new_n864), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n857), .B1(new_n902), .B2(new_n871), .ZN(new_n903));
  OAI21_X1  g717(.A(KEYINPUT114), .B1(new_n889), .B2(KEYINPUT53), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n880), .A2(new_n875), .A3(new_n881), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(G210), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n906), .A2(new_n907), .A3(new_n322), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n897), .B1(new_n908), .B2(KEYINPUT56), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n270), .A2(G952), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT121), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n913), .B1(new_n906), .B2(new_n322), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n873), .B1(new_n882), .B2(new_n883), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n915), .A2(KEYINPUT121), .A3(G902), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n914), .A2(new_n916), .A3(new_n400), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n897), .A2(KEYINPUT56), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n912), .B1(new_n917), .B2(new_n918), .ZN(G51));
  INV_X1    g733(.A(KEYINPUT122), .ZN(new_n920));
  INV_X1    g734(.A(new_n770), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n914), .A2(new_n916), .A3(new_n921), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n525), .B(KEYINPUT57), .Z(new_n923));
  INV_X1    g737(.A(new_n884), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n904), .A2(new_n905), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n874), .B1(new_n925), .B2(new_n873), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n923), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  OR2_X1    g741(.A1(new_n515), .A2(new_n523), .ZN(new_n928));
  AOI22_X1  g742(.A1(new_n920), .A2(new_n922), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  OR2_X1    g743(.A1(new_n922), .A2(new_n920), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n910), .B1(new_n929), .B2(new_n930), .ZN(G54));
  AND2_X1   g745(.A1(KEYINPUT58), .A2(G475), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n914), .A2(new_n916), .A3(new_n932), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n933), .A2(KEYINPUT123), .A3(new_n589), .ZN(new_n934));
  AOI21_X1  g748(.A(KEYINPUT123), .B1(new_n933), .B2(new_n589), .ZN(new_n935));
  INV_X1    g749(.A(new_n589), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n914), .A2(new_n916), .A3(new_n936), .A4(new_n932), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n911), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n934), .A2(new_n935), .A3(new_n938), .ZN(G60));
  XOR2_X1   g753(.A(new_n624), .B(KEYINPUT59), .Z(new_n940));
  AOI21_X1  g754(.A(new_n628), .B1(new_n891), .B2(new_n940), .ZN(new_n941));
  OR2_X1    g755(.A1(new_n924), .A2(new_n926), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n628), .A2(new_n940), .ZN(new_n943));
  AOI211_X1 g757(.A(new_n910), .B(new_n941), .C1(new_n942), .C2(new_n943), .ZN(G63));
  NAND2_X1  g758(.A1(G217), .A2(G902), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT60), .Z(new_n946));
  AOI21_X1  g760(.A(new_n382), .B1(new_n915), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n947), .A2(new_n910), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n915), .A2(new_n648), .A3(new_n946), .ZN(new_n949));
  XNOR2_X1  g763(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n950));
  AND3_X1   g764(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n950), .B1(new_n948), .B2(new_n949), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n951), .A2(new_n952), .ZN(G66));
  AOI21_X1  g767(.A(new_n270), .B1(new_n395), .B2(G224), .ZN(new_n954));
  INV_X1    g768(.A(new_n855), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n836), .A2(new_n837), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n954), .B1(new_n956), .B2(new_n270), .ZN(new_n957));
  INV_X1    g771(.A(G898), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n895), .B1(new_n958), .B2(G953), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n957), .B(new_n959), .ZN(G69));
  NAND2_X1  g774(.A1(new_n278), .A2(new_n280), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(new_n585), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n776), .A2(new_n622), .A3(new_n732), .A4(new_n819), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n780), .A2(new_n963), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n739), .A2(new_n677), .A3(new_n702), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n964), .A2(new_n785), .A3(new_n878), .A4(new_n965), .ZN(new_n966));
  AND2_X1   g780(.A1(new_n966), .A2(new_n270), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n962), .B1(new_n967), .B2(new_n666), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n742), .A2(new_n389), .A3(new_n694), .A4(new_n853), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n785), .A2(new_n780), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n965), .A2(new_n697), .ZN(new_n971));
  OR2_X1    g785(.A1(new_n971), .A2(KEYINPUT62), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(KEYINPUT62), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n970), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n974), .A2(new_n270), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n968), .B1(new_n962), .B2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(G227), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n666), .B1(new_n977), .B2(G953), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT125), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(new_n979), .ZN(new_n981));
  OAI211_X1 g795(.A(new_n968), .B(new_n981), .C1(new_n975), .C2(new_n962), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n980), .A2(new_n982), .ZN(G72));
  XNOR2_X1  g797(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n681), .B(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n986), .B1(new_n966), .B2(new_n956), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n987), .A2(new_n255), .A3(new_n281), .A4(new_n283), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n284), .A2(new_n308), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(new_n986), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n988), .B(new_n911), .C1(new_n890), .C2(new_n990), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n986), .B1(new_n974), .B2(new_n956), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n992), .B(KEYINPUT127), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n283), .B1(new_n281), .B2(new_n255), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n991), .B1(new_n993), .B2(new_n994), .ZN(G57));
endmodule


