

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783;

  BUF_X1 U381 ( .A(n739), .Z(n747) );
  AND2_X2 U382 ( .A1(n368), .A2(n513), .ZN(n739) );
  XNOR2_X1 U383 ( .A(n406), .B(n465), .ZN(n510) );
  XNOR2_X1 U384 ( .A(n501), .B(n500), .ZN(n595) );
  XNOR2_X1 U385 ( .A(n512), .B(n457), .ZN(n759) );
  INV_X1 U386 ( .A(G953), .ZN(n771) );
  NOR2_X2 U387 ( .A1(n603), .A2(n597), .ZN(n598) );
  NOR2_X2 U388 ( .A1(n754), .A2(n439), .ZN(n438) );
  NOR2_X2 U389 ( .A1(n560), .A2(n717), .ZN(n561) );
  XNOR2_X2 U390 ( .A(n578), .B(KEYINPUT32), .ZN(n783) );
  NOR2_X1 U391 ( .A1(n372), .A2(n371), .ZN(n370) );
  XNOR2_X1 U392 ( .A(n564), .B(n565), .ZN(n780) );
  AND2_X1 U393 ( .A1(n376), .A2(n397), .ZN(n684) );
  NOR2_X1 U394 ( .A1(n622), .A2(n621), .ZN(n628) );
  OR2_X1 U395 ( .A1(n697), .A2(n599), .ZN(n620) );
  NAND2_X1 U396 ( .A1(n448), .A2(n447), .ZN(n569) );
  NAND2_X2 U397 ( .A1(n424), .A2(n421), .ZN(n704) );
  XNOR2_X1 U398 ( .A(n392), .B(n651), .ZN(n653) );
  XNOR2_X1 U399 ( .A(n393), .B(G478), .ZN(n566) );
  XNOR2_X1 U400 ( .A(KEYINPUT23), .B(KEYINPUT95), .ZN(n486) );
  INV_X1 U401 ( .A(n700), .ZN(n402) );
  XNOR2_X1 U402 ( .A(n505), .B(n464), .ZN(n767) );
  NOR2_X1 U403 ( .A1(n587), .A2(n364), .ZN(n418) );
  XNOR2_X1 U404 ( .A(n411), .B(KEYINPUT109), .ZN(n636) );
  XOR2_X1 U405 ( .A(KEYINPUT79), .B(n593), .Z(n621) );
  NOR2_X1 U406 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U407 ( .A(n429), .B(KEYINPUT108), .ZN(n591) );
  NOR2_X1 U408 ( .A1(n590), .A2(n430), .ZN(n429) );
  XNOR2_X1 U409 ( .A(n559), .B(n558), .ZN(n717) );
  XNOR2_X1 U410 ( .A(n557), .B(KEYINPUT107), .ZN(n558) );
  NAND2_X1 U411 ( .A1(n616), .A2(n610), .ZN(n378) );
  INV_X1 U412 ( .A(KEYINPUT84), .ZN(n483) );
  NOR2_X1 U413 ( .A1(n684), .A2(n362), .ZN(n379) );
  XNOR2_X1 U414 ( .A(n596), .B(KEYINPUT70), .ZN(n603) );
  NOR2_X1 U415 ( .A1(G902), .A2(G237), .ZN(n514) );
  NOR2_X1 U416 ( .A1(G953), .A2(G237), .ZN(n533) );
  XOR2_X1 U417 ( .A(KEYINPUT97), .B(KEYINPUT11), .Z(n535) );
  XOR2_X1 U418 ( .A(KEYINPUT98), .B(KEYINPUT12), .Z(n532) );
  XNOR2_X1 U419 ( .A(G101), .B(G104), .ZN(n472) );
  XOR2_X1 U420 ( .A(G107), .B(G110), .Z(n473) );
  XOR2_X1 U421 ( .A(G137), .B(G140), .Z(n495) );
  XNOR2_X1 U422 ( .A(n767), .B(n419), .ZN(n477) );
  INV_X1 U423 ( .A(KEYINPUT4), .ZN(n420) );
  XNOR2_X1 U424 ( .A(n507), .B(n506), .ZN(n508) );
  INV_X1 U425 ( .A(KEYINPUT90), .ZN(n506) );
  XOR2_X1 U426 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n507) );
  XNOR2_X1 U427 ( .A(n419), .B(G125), .ZN(n504) );
  AND2_X1 U428 ( .A1(n782), .A2(n644), .ZN(n645) );
  INV_X1 U429 ( .A(n687), .ZN(n644) );
  INV_X1 U430 ( .A(G902), .ZN(n423) );
  NAND2_X1 U431 ( .A1(G472), .A2(G902), .ZN(n425) );
  XNOR2_X1 U432 ( .A(n547), .B(n458), .ZN(n457) );
  XNOR2_X1 U433 ( .A(n510), .B(n529), .ZN(n512) );
  XNOR2_X1 U434 ( .A(n511), .B(n459), .ZN(n458) );
  INV_X1 U435 ( .A(KEYINPUT45), .ZN(n441) );
  NAND2_X1 U436 ( .A1(n413), .A2(n416), .ZN(n368) );
  NAND2_X1 U437 ( .A1(n414), .A2(n363), .ZN(n413) );
  NAND2_X1 U438 ( .A1(n415), .A2(n722), .ZN(n414) );
  INV_X1 U439 ( .A(KEYINPUT115), .ZN(n435) );
  INV_X1 U440 ( .A(n606), .ZN(n433) );
  XNOR2_X1 U441 ( .A(n452), .B(KEYINPUT22), .ZN(n575) );
  NAND2_X1 U442 ( .A1(n389), .A2(n387), .ZN(n622) );
  XNOR2_X1 U443 ( .A(n619), .B(n388), .ZN(n387) );
  INV_X1 U444 ( .A(n620), .ZN(n389) );
  NOR2_X1 U445 ( .A1(n745), .A2(G902), .ZN(n393) );
  INV_X1 U446 ( .A(KEYINPUT6), .ZN(n427) );
  XNOR2_X1 U447 ( .A(n390), .B(G131), .ZN(n538) );
  NOR2_X1 U448 ( .A1(G952), .A2(n771), .ZN(n753) );
  INV_X1 U449 ( .A(KEYINPUT83), .ZN(n405) );
  AND2_X1 U450 ( .A1(n374), .A2(n377), .ZN(n373) );
  NAND2_X1 U451 ( .A1(n378), .A2(n382), .ZN(n377) );
  XNOR2_X1 U452 ( .A(n522), .B(KEYINPUT92), .ZN(n590) );
  NAND2_X1 U453 ( .A1(G953), .A2(n431), .ZN(n430) );
  INV_X1 U454 ( .A(G900), .ZN(n431) );
  XOR2_X1 U455 ( .A(G137), .B(KEYINPUT5), .Z(n466) );
  XNOR2_X1 U456 ( .A(G110), .B(KEYINPUT71), .ZN(n511) );
  INV_X1 U457 ( .A(KEYINPUT16), .ZN(n459) );
  XNOR2_X1 U458 ( .A(n407), .B(G113), .ZN(n406) );
  INV_X1 U459 ( .A(G101), .ZN(n407) );
  NOR2_X1 U460 ( .A1(n585), .A2(n582), .ZN(n583) );
  INV_X1 U461 ( .A(KEYINPUT94), .ZN(n482) );
  XNOR2_X1 U462 ( .A(n504), .B(n409), .ZN(n528) );
  INV_X1 U463 ( .A(KEYINPUT10), .ZN(n409) );
  XNOR2_X1 U464 ( .A(n519), .B(KEYINPUT14), .ZN(n521) );
  NAND2_X1 U465 ( .A1(G234), .A2(G237), .ZN(n519) );
  INV_X1 U466 ( .A(n588), .ZN(n693) );
  INV_X1 U467 ( .A(KEYINPUT30), .ZN(n388) );
  AND2_X1 U468 ( .A1(n450), .A2(n449), .ZN(n448) );
  NAND2_X1 U469 ( .A1(n446), .A2(n365), .ZN(n447) );
  XNOR2_X1 U470 ( .A(n499), .B(n498), .ZN(n500) );
  NOR2_X1 U471 ( .A1(n748), .A2(G902), .ZN(n501) );
  NAND2_X1 U472 ( .A1(n646), .A2(n645), .ZN(n765) );
  XNOR2_X1 U473 ( .A(G110), .B(KEYINPUT93), .ZN(n489) );
  XNOR2_X1 U474 ( .A(KEYINPUT85), .B(KEYINPUT8), .ZN(n480) );
  XOR2_X1 U475 ( .A(G116), .B(G107), .Z(n547) );
  XOR2_X1 U476 ( .A(KEYINPUT7), .B(KEYINPUT100), .Z(n549) );
  XNOR2_X1 U477 ( .A(G134), .B(G122), .ZN(n545) );
  XOR2_X1 U478 ( .A(KEYINPUT101), .B(KEYINPUT9), .Z(n546) );
  XOR2_X1 U479 ( .A(G104), .B(G122), .Z(n529) );
  XNOR2_X1 U480 ( .A(G113), .B(G140), .ZN(n531) );
  XNOR2_X1 U481 ( .A(n477), .B(n478), .ZN(n732) );
  XNOR2_X1 U482 ( .A(n456), .B(n455), .ZN(n454) );
  XNOR2_X1 U483 ( .A(n509), .B(n504), .ZN(n455) );
  XNOR2_X1 U484 ( .A(n505), .B(n508), .ZN(n456) );
  NAND2_X1 U485 ( .A1(n645), .A2(KEYINPUT2), .ZN(n437) );
  INV_X1 U486 ( .A(n416), .ZN(n725) );
  XNOR2_X1 U487 ( .A(n399), .B(n398), .ZN(n637) );
  INV_X1 U488 ( .A(KEYINPUT110), .ZN(n398) );
  NAND2_X1 U489 ( .A1(n636), .A2(n688), .ZN(n399) );
  XNOR2_X1 U490 ( .A(n682), .B(n394), .ZN(n642) );
  INV_X1 U491 ( .A(KEYINPUT103), .ZN(n394) );
  XNOR2_X1 U492 ( .A(n598), .B(KEYINPUT28), .ZN(n385) );
  OR2_X1 U493 ( .A1(n657), .A2(n422), .ZN(n421) );
  AND2_X1 U494 ( .A1(n426), .A2(n425), .ZN(n424) );
  NAND2_X1 U495 ( .A1(n471), .A2(n423), .ZN(n422) );
  XNOR2_X1 U496 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U497 ( .A(n444), .B(n442), .ZN(n745) );
  XNOR2_X1 U498 ( .A(n550), .B(n443), .ZN(n442) );
  XNOR2_X1 U499 ( .A(n552), .B(n445), .ZN(n444) );
  INV_X1 U500 ( .A(n547), .ZN(n443) );
  BUF_X1 U501 ( .A(n652), .Z(n392) );
  XNOR2_X1 U502 ( .A(n432), .B(n380), .ZN(n376) );
  INV_X1 U503 ( .A(KEYINPUT36), .ZN(n380) );
  AND2_X1 U504 ( .A1(n576), .A2(n396), .ZN(n578) );
  AND2_X1 U505 ( .A1(n618), .A2(n623), .ZN(n412) );
  BUF_X1 U506 ( .A(G143), .Z(n390) );
  NOR2_X1 U507 ( .A1(n553), .A2(n566), .ZN(n673) );
  BUF_X1 U508 ( .A(n678), .Z(n400) );
  NOR2_X1 U509 ( .A1(n742), .A2(n753), .ZN(n743) );
  XNOR2_X1 U510 ( .A(n731), .B(n410), .ZN(G75) );
  XNOR2_X1 U511 ( .A(KEYINPUT121), .B(KEYINPUT53), .ZN(n410) );
  XNOR2_X1 U512 ( .A(n606), .B(n518), .ZN(n600) );
  AND2_X1 U513 ( .A1(n602), .A2(n672), .ZN(n362) );
  AND2_X1 U514 ( .A1(n440), .A2(KEYINPUT74), .ZN(n363) );
  AND2_X1 U515 ( .A1(n555), .A2(n588), .ZN(n364) );
  XNOR2_X1 U516 ( .A(n698), .B(KEYINPUT89), .ZN(n397) );
  NOR2_X1 U517 ( .A1(n524), .A2(n451), .ZN(n365) );
  NOR2_X1 U518 ( .A1(n615), .A2(n614), .ZN(n366) );
  INV_X1 U519 ( .A(G146), .ZN(n419) );
  AND2_X1 U520 ( .A1(n628), .A2(n412), .ZN(n676) );
  XOR2_X1 U521 ( .A(G902), .B(KEYINPUT15), .Z(n513) );
  INV_X1 U522 ( .A(KEYINPUT80), .ZN(n382) );
  AND2_X1 U523 ( .A1(n513), .A2(G475), .ZN(n367) );
  NAND2_X1 U524 ( .A1(n368), .A2(n367), .ZN(n740) );
  NAND2_X1 U525 ( .A1(n373), .A2(n369), .ZN(n381) );
  NAND2_X1 U526 ( .A1(n370), .A2(n383), .ZN(n369) );
  INV_X1 U527 ( .A(n408), .ZN(n371) );
  NAND2_X1 U528 ( .A1(n611), .A2(KEYINPUT80), .ZN(n372) );
  NAND2_X1 U529 ( .A1(n375), .A2(n382), .ZN(n374) );
  NAND2_X1 U530 ( .A1(n408), .A2(n611), .ZN(n375) );
  INV_X1 U531 ( .A(n378), .ZN(n383) );
  NAND2_X1 U532 ( .A1(n381), .A2(n379), .ZN(n428) );
  INV_X1 U533 ( .A(n601), .ZN(n624) );
  XNOR2_X2 U534 ( .A(n384), .B(KEYINPUT113), .ZN(n601) );
  NAND2_X1 U535 ( .A1(n385), .A2(n391), .ZN(n384) );
  INV_X1 U536 ( .A(n599), .ZN(n391) );
  AND2_X1 U537 ( .A1(n418), .A2(n586), .ZN(n417) );
  XNOR2_X2 U538 ( .A(n386), .B(n441), .ZN(n754) );
  NAND2_X1 U539 ( .A1(n453), .A2(n417), .ZN(n386) );
  NOR2_X1 U540 ( .A1(n738), .A2(G902), .ZN(n544) );
  XNOR2_X1 U541 ( .A(n540), .B(n541), .ZN(n738) );
  XNOR2_X1 U542 ( .A(n759), .B(n454), .ZN(n652) );
  NOR2_X1 U543 ( .A1(n404), .A2(n366), .ZN(n408) );
  NOR2_X2 U544 ( .A1(n698), .A2(n697), .ZN(n556) );
  NAND2_X1 U545 ( .A1(n556), .A2(n605), .ZN(n559) );
  XNOR2_X2 U546 ( .A(n581), .B(KEYINPUT106), .ZN(n781) );
  NAND2_X1 U547 ( .A1(n649), .A2(n648), .ZN(n416) );
  XNOR2_X1 U548 ( .A(n676), .B(n405), .ZN(n404) );
  NOR2_X2 U549 ( .A1(n575), .A2(n571), .ZN(n580) );
  AND2_X2 U550 ( .A1(n580), .A2(n579), .ZN(n581) );
  NAND2_X1 U551 ( .A1(n617), .A2(n688), .ZN(n606) );
  NAND2_X1 U552 ( .A1(n551), .A2(G217), .ZN(n552) );
  XNOR2_X1 U553 ( .A(n481), .B(n480), .ZN(n551) );
  XNOR2_X1 U554 ( .A(n554), .B(KEYINPUT102), .ZN(n678) );
  XNOR2_X1 U555 ( .A(n636), .B(n435), .ZN(n434) );
  XNOR2_X2 U556 ( .A(n599), .B(KEYINPUT1), .ZN(n698) );
  NAND2_X1 U557 ( .A1(n780), .A2(KEYINPUT44), .ZN(n573) );
  BUF_X1 U558 ( .A(n595), .Z(n395) );
  NAND2_X1 U559 ( .A1(n594), .A2(n595), .ZN(n596) );
  AND2_X1 U560 ( .A1(n397), .A2(n577), .ZN(n396) );
  XNOR2_X1 U561 ( .A(n583), .B(KEYINPUT65), .ZN(n453) );
  NAND2_X1 U562 ( .A1(n401), .A2(n640), .ZN(n641) );
  XNOR2_X1 U563 ( .A(n638), .B(n639), .ZN(n401) );
  NAND2_X1 U564 ( .A1(n403), .A2(n402), .ZN(n697) );
  INV_X1 U565 ( .A(n595), .ZN(n403) );
  NOR2_X1 U566 ( .A1(n754), .A2(n437), .ZN(n436) );
  NOR2_X1 U567 ( .A1(G953), .A2(n728), .ZN(n729) );
  NAND2_X1 U568 ( .A1(n604), .A2(n605), .ZN(n411) );
  XNOR2_X1 U569 ( .A(n544), .B(n543), .ZN(n567) );
  NAND2_X1 U570 ( .A1(n434), .A2(n433), .ZN(n432) );
  XNOR2_X1 U571 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U572 ( .A(n488), .B(n460), .ZN(n492) );
  INV_X1 U573 ( .A(n649), .ZN(n415) );
  XNOR2_X2 U574 ( .A(n548), .B(n420), .ZN(n505) );
  XNOR2_X2 U575 ( .A(n462), .B(G128), .ZN(n548) );
  NAND2_X1 U576 ( .A1(n657), .A2(G472), .ZN(n426) );
  XNOR2_X2 U577 ( .A(n704), .B(n427), .ZN(n605) );
  XNOR2_X2 U578 ( .A(n479), .B(G469), .ZN(n599) );
  XNOR2_X1 U579 ( .A(n428), .B(KEYINPUT69), .ZN(n634) );
  AND2_X2 U580 ( .A1(n438), .A2(n646), .ZN(n649) );
  INV_X1 U581 ( .A(n645), .ZN(n439) );
  NAND2_X1 U582 ( .A1(n436), .A2(n646), .ZN(n440) );
  XNOR2_X1 U583 ( .A(n548), .B(n549), .ZN(n445) );
  INV_X1 U584 ( .A(n600), .ZN(n446) );
  NAND2_X1 U585 ( .A1(n600), .A2(n451), .ZN(n450) );
  NAND2_X1 U586 ( .A1(n524), .A2(n451), .ZN(n449) );
  INV_X1 U587 ( .A(KEYINPUT0), .ZN(n451) );
  NAND2_X1 U588 ( .A1(n569), .A2(n570), .ZN(n452) );
  INV_X2 U589 ( .A(G143), .ZN(n462) );
  NOR2_X1 U590 ( .A1(n704), .A2(n403), .ZN(n579) );
  XOR2_X1 U591 ( .A(G128), .B(G119), .Z(n460) );
  XOR2_X1 U592 ( .A(KEYINPUT68), .B(KEYINPUT48), .Z(n461) );
  XNOR2_X1 U593 ( .A(n466), .B(G116), .ZN(n467) );
  XNOR2_X1 U594 ( .A(n510), .B(n467), .ZN(n469) );
  XNOR2_X1 U595 ( .A(n469), .B(n468), .ZN(n470) );
  INV_X1 U596 ( .A(KEYINPUT25), .ZN(n498) );
  XNOR2_X1 U597 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U598 ( .A(n542), .B(G475), .ZN(n543) );
  XNOR2_X1 U599 ( .A(n748), .B(n749), .ZN(n750) );
  INV_X1 U600 ( .A(KEYINPUT63), .ZN(n663) );
  XNOR2_X1 U601 ( .A(n751), .B(n750), .ZN(n752) );
  XNOR2_X1 U602 ( .A(G134), .B(KEYINPUT67), .ZN(n463) );
  XNOR2_X1 U603 ( .A(n463), .B(G131), .ZN(n464) );
  XNOR2_X1 U604 ( .A(G119), .B(KEYINPUT3), .ZN(n465) );
  NAND2_X1 U605 ( .A1(n533), .A2(G210), .ZN(n468) );
  XNOR2_X1 U606 ( .A(n477), .B(n470), .ZN(n657) );
  INV_X1 U607 ( .A(G472), .ZN(n471) );
  XNOR2_X1 U608 ( .A(n473), .B(n472), .ZN(n474) );
  XOR2_X1 U609 ( .A(n495), .B(n474), .Z(n476) );
  NAND2_X1 U610 ( .A1(G227), .A2(n771), .ZN(n475) );
  XNOR2_X1 U611 ( .A(n476), .B(n475), .ZN(n478) );
  NOR2_X1 U612 ( .A1(n732), .A2(G902), .ZN(n479) );
  NAND2_X1 U613 ( .A1(n771), .A2(G234), .ZN(n481) );
  NAND2_X1 U614 ( .A1(n551), .A2(G221), .ZN(n494) );
  NAND2_X1 U615 ( .A1(KEYINPUT84), .A2(n482), .ZN(n485) );
  NAND2_X1 U616 ( .A1(n483), .A2(KEYINPUT94), .ZN(n484) );
  NAND2_X1 U617 ( .A1(n485), .A2(n484), .ZN(n487) );
  XNOR2_X1 U618 ( .A(n487), .B(n486), .ZN(n488) );
  XOR2_X1 U619 ( .A(KEYINPUT75), .B(KEYINPUT24), .Z(n490) );
  XNOR2_X1 U620 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U621 ( .A(n493), .B(n494), .ZN(n496) );
  XOR2_X1 U622 ( .A(n495), .B(n528), .Z(n766) );
  XNOR2_X1 U623 ( .A(n496), .B(n766), .ZN(n748) );
  INV_X1 U624 ( .A(n513), .ZN(n650) );
  NAND2_X1 U625 ( .A1(G234), .A2(n650), .ZN(n497) );
  XNOR2_X1 U626 ( .A(KEYINPUT20), .B(n497), .ZN(n502) );
  NAND2_X1 U627 ( .A1(G217), .A2(n502), .ZN(n499) );
  NAND2_X1 U628 ( .A1(n502), .A2(G221), .ZN(n503) );
  XNOR2_X1 U629 ( .A(n503), .B(KEYINPUT21), .ZN(n700) );
  NAND2_X1 U630 ( .A1(n704), .A2(n556), .ZN(n707) );
  NAND2_X1 U631 ( .A1(G224), .A2(n771), .ZN(n509) );
  NOR2_X1 U632 ( .A1(n652), .A2(n513), .ZN(n516) );
  XNOR2_X1 U633 ( .A(n514), .B(KEYINPUT73), .ZN(n517) );
  NAND2_X1 U634 ( .A1(G210), .A2(n517), .ZN(n515) );
  XNOR2_X1 U635 ( .A(n516), .B(n515), .ZN(n617) );
  NAND2_X1 U636 ( .A1(G214), .A2(n517), .ZN(n688) );
  XOR2_X1 U637 ( .A(KEYINPUT19), .B(KEYINPUT66), .Z(n518) );
  NAND2_X1 U638 ( .A1(G952), .A2(n521), .ZN(n716) );
  NOR2_X1 U639 ( .A1(G953), .A2(n716), .ZN(n592) );
  NOR2_X1 U640 ( .A1(G898), .A2(n771), .ZN(n520) );
  XNOR2_X1 U641 ( .A(KEYINPUT91), .B(n520), .ZN(n760) );
  NAND2_X1 U642 ( .A1(n521), .A2(G902), .ZN(n522) );
  NOR2_X1 U643 ( .A1(n760), .A2(n590), .ZN(n523) );
  NOR2_X1 U644 ( .A1(n592), .A2(n523), .ZN(n524) );
  INV_X1 U645 ( .A(n569), .ZN(n560) );
  NOR2_X1 U646 ( .A1(n707), .A2(n560), .ZN(n525) );
  XNOR2_X1 U647 ( .A(n525), .B(KEYINPUT31), .ZN(n681) );
  NOR2_X1 U648 ( .A1(n560), .A2(n620), .ZN(n526) );
  INV_X1 U649 ( .A(n704), .ZN(n597) );
  NAND2_X1 U650 ( .A1(n526), .A2(n597), .ZN(n667) );
  NAND2_X1 U651 ( .A1(n681), .A2(n667), .ZN(n527) );
  XNOR2_X1 U652 ( .A(n527), .B(KEYINPUT96), .ZN(n555) );
  INV_X1 U653 ( .A(n528), .ZN(n530) );
  XNOR2_X1 U654 ( .A(n530), .B(n529), .ZN(n541) );
  XNOR2_X1 U655 ( .A(n532), .B(n531), .ZN(n537) );
  NAND2_X1 U656 ( .A1(G214), .A2(n533), .ZN(n534) );
  XNOR2_X1 U657 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U658 ( .A(n536), .B(n537), .ZN(n539) );
  XNOR2_X1 U659 ( .A(KEYINPUT13), .B(KEYINPUT99), .ZN(n542) );
  INV_X1 U660 ( .A(n567), .ZN(n553) );
  XNOR2_X1 U661 ( .A(n546), .B(n545), .ZN(n550) );
  INV_X1 U662 ( .A(n673), .ZN(n682) );
  NAND2_X1 U663 ( .A1(n566), .A2(n553), .ZN(n554) );
  NAND2_X1 U664 ( .A1(n642), .A2(n678), .ZN(n588) );
  XNOR2_X1 U665 ( .A(KEYINPUT35), .B(KEYINPUT76), .ZN(n565) );
  XOR2_X1 U666 ( .A(KEYINPUT33), .B(KEYINPUT87), .Z(n557) );
  XNOR2_X1 U667 ( .A(n561), .B(KEYINPUT34), .ZN(n563) );
  NOR2_X1 U668 ( .A1(n567), .A2(n566), .ZN(n623) );
  XOR2_X1 U669 ( .A(n623), .B(KEYINPUT77), .Z(n562) );
  NAND2_X1 U670 ( .A1(n563), .A2(n562), .ZN(n564) );
  NAND2_X1 U671 ( .A1(n567), .A2(n566), .ZN(n691) );
  NOR2_X1 U672 ( .A1(n700), .A2(n691), .ZN(n568) );
  XNOR2_X1 U673 ( .A(KEYINPUT104), .B(n568), .ZN(n570) );
  INV_X1 U674 ( .A(n698), .ZN(n571) );
  XOR2_X1 U675 ( .A(KEYINPUT105), .B(n395), .Z(n701) );
  NOR2_X1 U676 ( .A1(n605), .A2(n701), .ZN(n572) );
  NAND2_X1 U677 ( .A1(n580), .A2(n572), .ZN(n665) );
  NAND2_X1 U678 ( .A1(n573), .A2(n665), .ZN(n587) );
  XOR2_X1 U679 ( .A(KEYINPUT78), .B(n605), .Z(n577) );
  INV_X1 U680 ( .A(n701), .ZN(n574) );
  NOR2_X1 U681 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U682 ( .A1(n783), .A2(n781), .ZN(n585) );
  INV_X1 U683 ( .A(KEYINPUT44), .ZN(n582) );
  NOR2_X1 U684 ( .A1(KEYINPUT44), .A2(n780), .ZN(n584) );
  NAND2_X1 U685 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U686 ( .A1(n693), .A2(KEYINPUT47), .ZN(n589) );
  XNOR2_X1 U687 ( .A(KEYINPUT72), .B(n589), .ZN(n602) );
  NOR2_X1 U688 ( .A1(n700), .A2(n621), .ZN(n594) );
  NAND2_X2 U689 ( .A1(n601), .A2(n446), .ZN(n613) );
  INV_X1 U690 ( .A(n613), .ZN(n672) );
  NOR2_X1 U691 ( .A1(n678), .A2(n603), .ZN(n604) );
  NAND2_X1 U692 ( .A1(n613), .A2(KEYINPUT47), .ZN(n607) );
  NAND2_X1 U693 ( .A1(n607), .A2(KEYINPUT81), .ZN(n611) );
  INV_X1 U694 ( .A(KEYINPUT82), .ZN(n609) );
  NAND2_X1 U695 ( .A1(n693), .A2(KEYINPUT47), .ZN(n608) );
  NAND2_X1 U696 ( .A1(n609), .A2(n608), .ZN(n610) );
  INV_X1 U697 ( .A(KEYINPUT47), .ZN(n615) );
  NOR2_X1 U698 ( .A1(KEYINPUT81), .A2(n615), .ZN(n612) );
  NAND2_X1 U699 ( .A1(n613), .A2(n612), .ZN(n616) );
  NAND2_X1 U700 ( .A1(KEYINPUT82), .A2(n693), .ZN(n614) );
  BUF_X1 U701 ( .A(n617), .Z(n618) );
  INV_X1 U702 ( .A(n618), .ZN(n640) );
  NAND2_X1 U703 ( .A1(n704), .A2(n688), .ZN(n619) );
  XNOR2_X1 U704 ( .A(n640), .B(KEYINPUT38), .ZN(n689) );
  NAND2_X1 U705 ( .A1(n689), .A2(n688), .ZN(n692) );
  NOR2_X1 U706 ( .A1(n691), .A2(n692), .ZN(n626) );
  XNOR2_X1 U707 ( .A(KEYINPUT114), .B(KEYINPUT41), .ZN(n625) );
  XNOR2_X1 U708 ( .A(n626), .B(n625), .ZN(n718) );
  NOR2_X1 U709 ( .A1(n624), .A2(n718), .ZN(n627) );
  XNOR2_X1 U710 ( .A(n627), .B(KEYINPUT42), .ZN(n779) );
  AND2_X1 U711 ( .A1(n689), .A2(n628), .ZN(n629) );
  XNOR2_X1 U712 ( .A(KEYINPUT39), .B(n629), .ZN(n643) );
  NOR2_X1 U713 ( .A1(n643), .A2(n400), .ZN(n630) );
  XNOR2_X1 U714 ( .A(n630), .B(KEYINPUT40), .ZN(n778) );
  NOR2_X1 U715 ( .A1(n779), .A2(n778), .ZN(n632) );
  XNOR2_X1 U716 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n631) );
  XNOR2_X1 U717 ( .A(n632), .B(n631), .ZN(n633) );
  NAND2_X1 U718 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X2 U719 ( .A(n635), .B(n461), .ZN(n646) );
  XOR2_X1 U720 ( .A(KEYINPUT43), .B(KEYINPUT111), .Z(n639) );
  NAND2_X1 U721 ( .A1(n637), .A2(n698), .ZN(n638) );
  XNOR2_X1 U722 ( .A(n641), .B(KEYINPUT112), .ZN(n782) );
  NOR2_X1 U723 ( .A1(n643), .A2(n642), .ZN(n687) );
  INV_X1 U724 ( .A(KEYINPUT74), .ZN(n647) );
  AND2_X1 U725 ( .A1(KEYINPUT2), .A2(n647), .ZN(n648) );
  NAND2_X1 U726 ( .A1(n739), .A2(G210), .ZN(n654) );
  XOR2_X1 U727 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n651) );
  XNOR2_X1 U728 ( .A(n654), .B(n653), .ZN(n655) );
  NOR2_X2 U729 ( .A1(n655), .A2(n753), .ZN(n656) );
  XNOR2_X1 U730 ( .A(n656), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U731 ( .A1(n739), .A2(G472), .ZN(n661) );
  XOR2_X1 U732 ( .A(n657), .B(KEYINPUT116), .Z(n659) );
  XOR2_X1 U733 ( .A(KEYINPUT88), .B(KEYINPUT62), .Z(n658) );
  XNOR2_X1 U734 ( .A(n661), .B(n660), .ZN(n662) );
  NOR2_X2 U735 ( .A1(n662), .A2(n753), .ZN(n664) );
  XNOR2_X1 U736 ( .A(n664), .B(n663), .ZN(G57) );
  XNOR2_X1 U737 ( .A(G101), .B(n665), .ZN(G3) );
  NOR2_X1 U738 ( .A1(n400), .A2(n667), .ZN(n666) );
  XOR2_X1 U739 ( .A(G104), .B(n666), .Z(G6) );
  NOR2_X1 U740 ( .A1(n667), .A2(n682), .ZN(n671) );
  XOR2_X1 U741 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n669) );
  XNOR2_X1 U742 ( .A(G107), .B(KEYINPUT117), .ZN(n668) );
  XNOR2_X1 U743 ( .A(n669), .B(n668), .ZN(n670) );
  XNOR2_X1 U744 ( .A(n671), .B(n670), .ZN(G9) );
  XOR2_X1 U745 ( .A(G128), .B(KEYINPUT29), .Z(n675) );
  NAND2_X1 U746 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U747 ( .A(n675), .B(n674), .ZN(G30) );
  XOR2_X1 U748 ( .A(n390), .B(n676), .Z(G45) );
  OR2_X1 U749 ( .A1(n400), .A2(n613), .ZN(n677) );
  XNOR2_X1 U750 ( .A(n677), .B(G146), .ZN(G48) );
  NOR2_X1 U751 ( .A1(n400), .A2(n681), .ZN(n679) );
  XOR2_X1 U752 ( .A(KEYINPUT118), .B(n679), .Z(n680) );
  XNOR2_X1 U753 ( .A(G113), .B(n680), .ZN(G15) );
  NOR2_X1 U754 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U755 ( .A(G116), .B(n683), .Z(G18) );
  XOR2_X1 U756 ( .A(KEYINPUT37), .B(KEYINPUT119), .Z(n686) );
  XNOR2_X1 U757 ( .A(G125), .B(n684), .ZN(n685) );
  XNOR2_X1 U758 ( .A(n686), .B(n685), .ZN(G27) );
  XOR2_X1 U759 ( .A(G134), .B(n687), .Z(G36) );
  NOR2_X1 U760 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U761 ( .A1(n691), .A2(n690), .ZN(n695) );
  NOR2_X1 U762 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U763 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U764 ( .A1(n696), .A2(n717), .ZN(n712) );
  NAND2_X1 U765 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U766 ( .A(n699), .B(KEYINPUT50), .ZN(n706) );
  NAND2_X1 U767 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U768 ( .A(KEYINPUT49), .B(n702), .ZN(n703) );
  NOR2_X1 U769 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U770 ( .A1(n706), .A2(n705), .ZN(n708) );
  NAND2_X1 U771 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U772 ( .A(KEYINPUT51), .B(n709), .ZN(n710) );
  NOR2_X1 U773 ( .A1(n718), .A2(n710), .ZN(n711) );
  NOR2_X1 U774 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U775 ( .A(n713), .B(KEYINPUT52), .ZN(n714) );
  XNOR2_X1 U776 ( .A(KEYINPUT120), .B(n714), .ZN(n715) );
  NOR2_X1 U777 ( .A1(n716), .A2(n715), .ZN(n720) );
  NOR2_X1 U778 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X1 U779 ( .A1(n720), .A2(n719), .ZN(n730) );
  INV_X1 U780 ( .A(KEYINPUT2), .ZN(n722) );
  NAND2_X1 U781 ( .A1(n765), .A2(n722), .ZN(n721) );
  XNOR2_X1 U782 ( .A(n721), .B(KEYINPUT86), .ZN(n724) );
  NAND2_X1 U783 ( .A1(n754), .A2(n722), .ZN(n723) );
  NAND2_X1 U784 ( .A1(n724), .A2(n723), .ZN(n727) );
  NOR2_X1 U785 ( .A1(n725), .A2(n363), .ZN(n726) );
  NOR2_X1 U786 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U787 ( .A1(n730), .A2(n729), .ZN(n731) );
  XOR2_X1 U788 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n734) );
  XNOR2_X1 U789 ( .A(n732), .B(KEYINPUT122), .ZN(n733) );
  XNOR2_X1 U790 ( .A(n734), .B(n733), .ZN(n736) );
  NAND2_X1 U791 ( .A1(n747), .A2(G469), .ZN(n735) );
  XNOR2_X1 U792 ( .A(n736), .B(n735), .ZN(n737) );
  NOR2_X1 U793 ( .A1(n753), .A2(n737), .ZN(G54) );
  XOR2_X1 U794 ( .A(n738), .B(KEYINPUT59), .Z(n741) );
  XNOR2_X1 U795 ( .A(n741), .B(n740), .ZN(n742) );
  XNOR2_X1 U796 ( .A(n743), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U797 ( .A1(G478), .A2(n747), .ZN(n744) );
  XNOR2_X1 U798 ( .A(n745), .B(n744), .ZN(n746) );
  NOR2_X1 U799 ( .A1(n753), .A2(n746), .ZN(G63) );
  NAND2_X1 U800 ( .A1(n747), .A2(G217), .ZN(n751) );
  INV_X1 U801 ( .A(KEYINPUT123), .ZN(n749) );
  NOR2_X1 U802 ( .A1(n753), .A2(n752), .ZN(G66) );
  OR2_X1 U803 ( .A1(G953), .A2(n754), .ZN(n758) );
  NAND2_X1 U804 ( .A1(G953), .A2(G224), .ZN(n755) );
  XNOR2_X1 U805 ( .A(KEYINPUT61), .B(n755), .ZN(n756) );
  NAND2_X1 U806 ( .A1(n756), .A2(G898), .ZN(n757) );
  NAND2_X1 U807 ( .A1(n758), .A2(n757), .ZN(n764) );
  XNOR2_X1 U808 ( .A(n759), .B(KEYINPUT124), .ZN(n761) );
  NAND2_X1 U809 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U810 ( .A(n762), .B(KEYINPUT125), .ZN(n763) );
  XNOR2_X1 U811 ( .A(n764), .B(n763), .ZN(G69) );
  XNOR2_X1 U812 ( .A(KEYINPUT127), .B(n765), .ZN(n770) );
  XNOR2_X1 U813 ( .A(n766), .B(KEYINPUT126), .ZN(n768) );
  XOR2_X1 U814 ( .A(n767), .B(n768), .Z(n773) );
  INV_X1 U815 ( .A(n773), .ZN(n769) );
  XOR2_X1 U816 ( .A(n770), .B(n769), .Z(n772) );
  NAND2_X1 U817 ( .A1(n772), .A2(n771), .ZN(n777) );
  XOR2_X1 U818 ( .A(G227), .B(n773), .Z(n774) );
  NAND2_X1 U819 ( .A1(n774), .A2(G900), .ZN(n775) );
  NAND2_X1 U820 ( .A1(n775), .A2(G953), .ZN(n776) );
  NAND2_X1 U821 ( .A1(n777), .A2(n776), .ZN(G72) );
  XOR2_X1 U822 ( .A(G131), .B(n778), .Z(G33) );
  XOR2_X1 U823 ( .A(G137), .B(n779), .Z(G39) );
  XOR2_X1 U824 ( .A(n780), .B(G122), .Z(G24) );
  XOR2_X1 U825 ( .A(n781), .B(G110), .Z(G12) );
  XNOR2_X1 U826 ( .A(G140), .B(n782), .ZN(G42) );
  XOR2_X1 U827 ( .A(G119), .B(n783), .Z(G21) );
endmodule

