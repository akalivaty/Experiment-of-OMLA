//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 0 1 1 1 1 1 0 1 0 1 1 1 1 0 1 0 0 1 0 0 1 1 1 1 1 0 1 0 1 1 1 1 0 0 1 0 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:45 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1267,
    new_n1268, new_n1269, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(new_n206), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT64), .Z(new_n214));
  NAND2_X1  g0014(.A1(new_n202), .A2(G50), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT65), .Z(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n220));
  NAND3_X1  g0020(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n208), .B1(new_n217), .B2(new_n221), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n211), .B1(new_n214), .B2(new_n215), .C1(new_n222), .C2(KEYINPUT1), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XOR2_X1   g0024(.A(G238), .B(G244), .Z(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(G232), .ZN(new_n226));
  XOR2_X1   g0026(.A(KEYINPUT2), .B(G226), .Z(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(G250), .B(G257), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G264), .B(G270), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n228), .B(new_n231), .Z(G358));
  XOR2_X1   g0032(.A(G58), .B(G77), .Z(new_n233));
  XNOR2_X1  g0033(.A(G50), .B(G68), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G87), .B(G97), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G107), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n235), .B(new_n238), .Z(G351));
  XNOR2_X1  g0039(.A(G58), .B(G68), .ZN(new_n240));
  NOR2_X1   g0040(.A1(G20), .A2(G33), .ZN(new_n241));
  AOI22_X1  g0041(.A1(new_n240), .A2(G20), .B1(G159), .B2(new_n241), .ZN(new_n242));
  INV_X1    g0042(.A(G33), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(KEYINPUT3), .ZN(new_n244));
  INV_X1    g0044(.A(KEYINPUT3), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g0047(.A(KEYINPUT7), .B1(new_n247), .B2(new_n206), .ZN(new_n248));
  NOR2_X1   g0048(.A1(new_n243), .A2(KEYINPUT3), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n245), .A2(KEYINPUT72), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT72), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n249), .B1(new_n253), .B2(new_n243), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT7), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n255), .A2(G20), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  OAI21_X1  g0057(.A(KEYINPUT74), .B1(new_n254), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT74), .ZN(new_n259));
  AOI21_X1  g0059(.A(G33), .B1(new_n250), .B2(new_n252), .ZN(new_n260));
  OAI211_X1 g0060(.A(new_n259), .B(new_n256), .C1(new_n260), .C2(new_n249), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n248), .B1(new_n258), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G68), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n242), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT16), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n244), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT72), .B(KEYINPUT3), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n267), .B1(new_n268), .B2(G33), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n269), .A2(new_n257), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n250), .A2(new_n252), .A3(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(new_n244), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT73), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n271), .A2(KEYINPUT73), .A3(new_n244), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n274), .A2(new_n206), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n270), .B1(new_n276), .B2(new_n255), .ZN(new_n277));
  OAI211_X1 g0077(.A(KEYINPUT16), .B(new_n242), .C1(new_n277), .C2(new_n263), .ZN(new_n278));
  NAND3_X1  g0078(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n212), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n266), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT8), .B(G58), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n282), .B1(new_n205), .B2(G20), .ZN(new_n283));
  INV_X1    g0083(.A(G13), .ZN(new_n284));
  NOR3_X1   g0084(.A1(new_n284), .A2(new_n206), .A3(G1), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n285), .A2(new_n280), .ZN(new_n286));
  AOI22_X1  g0086(.A1(new_n283), .A2(new_n286), .B1(new_n285), .B2(new_n282), .ZN(new_n287));
  AND2_X1   g0087(.A1(new_n281), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n212), .B1(G33), .B2(G41), .ZN(new_n289));
  INV_X1    g0089(.A(G41), .ZN(new_n290));
  INV_X1    g0090(.A(G45), .ZN(new_n291));
  AOI21_X1  g0091(.A(G1), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G232), .ZN(new_n294));
  OAI211_X1 g0094(.A(G1), .B(G13), .C1(new_n243), .C2(new_n290), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n295), .A2(G274), .A3(new_n292), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G223), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n298), .A2(G1698), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n271), .A2(new_n244), .A3(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT75), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n271), .A2(KEYINPUT75), .A3(new_n244), .A4(new_n299), .ZN(new_n303));
  NAND2_X1  g0103(.A1(G33), .A2(G87), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n271), .A2(G226), .A3(G1698), .A4(new_n244), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n302), .A2(new_n303), .A3(new_n304), .A4(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n297), .B1(new_n306), .B2(new_n289), .ZN(new_n307));
  INV_X1    g0107(.A(G169), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G179), .ZN(new_n310));
  AOI211_X1 g0110(.A(new_n310), .B(new_n297), .C1(new_n306), .C2(new_n289), .ZN(new_n311));
  OAI21_X1  g0111(.A(KEYINPUT76), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n307), .A2(G179), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT76), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n313), .B(new_n314), .C1(new_n308), .C2(new_n307), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(KEYINPUT18), .B1(new_n288), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT17), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT77), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n306), .A2(new_n289), .ZN(new_n320));
  INV_X1    g0120(.A(new_n297), .ZN(new_n321));
  AOI21_X1  g0121(.A(G200), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  AOI211_X1 g0122(.A(G190), .B(new_n297), .C1(new_n306), .C2(new_n289), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n319), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G190), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n320), .A2(new_n325), .A3(new_n321), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n326), .B(KEYINPUT77), .C1(G200), .C2(new_n307), .ZN(new_n327));
  AND2_X1   g0127(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n281), .A2(new_n287), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n318), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n324), .A2(new_n327), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n331), .A2(KEYINPUT17), .A3(new_n281), .A4(new_n287), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT18), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n329), .A2(new_n333), .A3(new_n312), .A4(new_n315), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n317), .A2(new_n330), .A3(new_n332), .A4(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n247), .A2(G1698), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(G222), .ZN(new_n337));
  INV_X1    g0137(.A(G77), .ZN(new_n338));
  INV_X1    g0138(.A(new_n247), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(G1698), .ZN(new_n340));
  OAI221_X1 g0140(.A(new_n337), .B1(new_n338), .B2(new_n339), .C1(new_n298), .C2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n289), .ZN(new_n342));
  INV_X1    g0142(.A(new_n296), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n343), .B1(G226), .B2(new_n293), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(G200), .ZN(new_n346));
  INV_X1    g0146(.A(new_n280), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n206), .A2(G33), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n282), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n349), .B1(G150), .B2(new_n241), .ZN(new_n350));
  OAI21_X1  g0150(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n347), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n205), .A2(G20), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n286), .A2(G50), .A3(new_n353), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n284), .A2(G1), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(G20), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n354), .B1(G50), .B2(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n352), .A2(new_n357), .ZN(new_n358));
  OR2_X1    g0158(.A1(new_n358), .A2(KEYINPUT9), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n342), .A2(G190), .A3(new_n344), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n358), .A2(KEYINPUT9), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n346), .A2(new_n359), .A3(new_n360), .A4(new_n361), .ZN(new_n362));
  XNOR2_X1  g0162(.A(new_n362), .B(KEYINPUT10), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n358), .B1(new_n345), .B2(new_n308), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(G179), .B2(new_n345), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n241), .A2(G50), .ZN(new_n367));
  XNOR2_X1  g0167(.A(new_n367), .B(KEYINPUT71), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n348), .A2(new_n338), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n369), .B1(G20), .B2(new_n263), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n347), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  OR2_X1    g0171(.A1(new_n371), .A2(KEYINPUT11), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n356), .A2(KEYINPUT68), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT68), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n285), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n376), .A2(new_n280), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n377), .A2(G68), .A3(new_n353), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n371), .A2(KEYINPUT11), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n356), .A2(KEYINPUT68), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n285), .A2(new_n374), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(KEYINPUT12), .B1(new_n382), .B2(G68), .ZN(new_n383));
  NOR3_X1   g0183(.A1(new_n206), .A2(KEYINPUT12), .A3(G68), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n355), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n372), .A2(new_n378), .A3(new_n379), .A4(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n343), .B1(G238), .B2(new_n293), .ZN(new_n388));
  INV_X1    g0188(.A(G1698), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n244), .A2(new_n246), .A3(G226), .A4(new_n389), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n244), .A2(new_n246), .A3(G232), .A4(G1698), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G33), .A2(G97), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  AND3_X1   g0193(.A1(new_n393), .A2(KEYINPUT70), .A3(new_n289), .ZN(new_n394));
  AOI21_X1  g0194(.A(KEYINPUT70), .B1(new_n393), .B2(new_n289), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n388), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(KEYINPUT13), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT13), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n398), .B(new_n388), .C1(new_n394), .C2(new_n395), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT14), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n400), .A2(new_n401), .A3(G169), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n397), .A2(G179), .A3(new_n399), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n401), .B1(new_n400), .B2(G169), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n387), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n387), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(new_n400), .B2(new_n325), .ZN(new_n408));
  INV_X1    g0208(.A(G200), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n409), .B1(new_n397), .B2(new_n399), .ZN(new_n410));
  OR2_X1    g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n406), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n336), .A2(G232), .ZN(new_n413));
  OR2_X1    g0213(.A1(KEYINPUT67), .A2(G107), .ZN(new_n414));
  NAND2_X1  g0214(.A1(KEYINPUT67), .A2(G107), .ZN(new_n415));
  AND2_X1   g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(G238), .ZN(new_n417));
  OAI221_X1 g0217(.A(new_n413), .B1(new_n339), .B2(new_n416), .C1(new_n417), .C2(new_n340), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n289), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n293), .A2(G244), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n296), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT66), .ZN(new_n422));
  OR2_X1    g0222(.A1(new_n421), .A2(KEYINPUT66), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n419), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  OR2_X1    g0224(.A1(new_n424), .A2(G179), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n382), .A2(G77), .ZN(new_n426));
  XNOR2_X1  g0226(.A(new_n426), .B(KEYINPUT69), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n338), .B1(new_n205), .B2(G20), .ZN(new_n428));
  INV_X1    g0228(.A(new_n282), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n429), .A2(new_n241), .B1(G20), .B2(G77), .ZN(new_n430));
  XNOR2_X1  g0230(.A(KEYINPUT15), .B(G87), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n430), .B1(new_n348), .B2(new_n431), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n377), .A2(new_n428), .B1(new_n432), .B2(new_n280), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n427), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n424), .A2(new_n308), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n425), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n424), .A2(G200), .ZN(new_n437));
  INV_X1    g0237(.A(new_n434), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n437), .B(new_n438), .C1(new_n325), .C2(new_n424), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  NOR4_X1   g0240(.A1(new_n335), .A2(new_n366), .A3(new_n412), .A4(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  AND2_X1   g0242(.A1(KEYINPUT5), .A2(G41), .ZN(new_n443));
  NOR2_X1   g0243(.A1(KEYINPUT5), .A2(G41), .ZN(new_n444));
  OR2_X1    g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n291), .A2(G1), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n445), .A2(new_n295), .A3(G274), .A4(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n446), .B1(new_n443), .B2(new_n444), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n295), .ZN(new_n449));
  INV_X1    g0249(.A(G257), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n447), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT4), .ZN(new_n452));
  INV_X1    g0252(.A(G244), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n453), .A2(G1698), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n452), .B1(new_n272), .B2(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n452), .A2(new_n453), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n457), .A2(new_n389), .A3(new_n244), .A4(new_n246), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n244), .A2(new_n246), .A3(G250), .A4(G1698), .ZN(new_n459));
  NAND2_X1  g0259(.A1(G33), .A2(G283), .ZN(new_n460));
  AND3_X1   g0260(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n295), .B1(new_n462), .B2(KEYINPUT79), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT79), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n456), .A2(new_n461), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n451), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n310), .ZN(new_n467));
  AOI21_X1  g0267(.A(KEYINPUT4), .B1(new_n269), .B2(new_n454), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n469));
  OAI21_X1  g0269(.A(KEYINPUT79), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n470), .A2(new_n289), .A3(new_n465), .ZN(new_n471));
  INV_X1    g0271(.A(new_n451), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n308), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n356), .A2(G97), .ZN(new_n475));
  AOI211_X1 g0275(.A(new_n280), .B(new_n285), .C1(new_n205), .C2(G33), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n475), .B1(new_n476), .B2(G97), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n241), .A2(G77), .ZN(new_n478));
  OR2_X1    g0278(.A1(KEYINPUT78), .A2(G97), .ZN(new_n479));
  NAND2_X1  g0279(.A1(KEYINPUT78), .A2(G97), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(G107), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n481), .A2(KEYINPUT6), .A3(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT6), .ZN(new_n484));
  INV_X1    g0284(.A(G97), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n485), .A2(new_n482), .ZN(new_n486));
  NOR2_X1   g0286(.A1(G97), .A2(G107), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n484), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n483), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n478), .B1(new_n489), .B2(new_n206), .ZN(new_n490));
  INV_X1    g0290(.A(new_n248), .ZN(new_n491));
  INV_X1    g0291(.A(new_n261), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n246), .B1(new_n268), .B2(G33), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n259), .B1(new_n493), .B2(new_n256), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n491), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n414), .A2(new_n415), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n490), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n477), .B1(new_n497), .B2(new_n347), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n467), .A2(new_n474), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n466), .A2(G190), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n473), .A2(G200), .ZN(new_n501));
  INV_X1    g0301(.A(new_n477), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n483), .A2(new_n488), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n503), .A2(G20), .B1(G77), .B2(new_n241), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n504), .B1(new_n262), .B2(new_n416), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n502), .B1(new_n505), .B2(new_n280), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n500), .A2(new_n501), .A3(new_n506), .ZN(new_n507));
  AND2_X1   g0307(.A1(new_n499), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT24), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT22), .ZN(new_n510));
  INV_X1    g0310(.A(G87), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n510), .B1(new_n247), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(KEYINPUT22), .B1(KEYINPUT23), .B2(G107), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(G20), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n271), .A2(KEYINPUT22), .A3(G87), .A4(new_n244), .ZN(new_n517));
  AOI21_X1  g0317(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n518));
  AND2_X1   g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n206), .B1(new_n496), .B2(KEYINPUT23), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n509), .B(new_n516), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n520), .B1(new_n517), .B2(new_n518), .ZN(new_n522));
  OAI21_X1  g0322(.A(KEYINPUT24), .B1(new_n522), .B2(new_n515), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n280), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n285), .A2(new_n482), .ZN(new_n526));
  OR2_X1    g0326(.A1(new_n526), .A2(KEYINPUT84), .ZN(new_n527));
  XOR2_X1   g0327(.A(KEYINPUT83), .B(KEYINPUT25), .Z(new_n528));
  AOI21_X1  g0328(.A(new_n528), .B1(new_n526), .B2(KEYINPUT84), .ZN(new_n529));
  OR2_X1    g0329(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n476), .A2(G107), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n527), .A2(new_n529), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  NOR2_X1   g0334(.A1(G250), .A2(G1698), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n535), .B1(new_n450), .B2(G1698), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n536), .A2(new_n271), .A3(new_n244), .ZN(new_n537));
  NAND2_X1  g0337(.A1(G33), .A2(G294), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n289), .ZN(new_n540));
  INV_X1    g0340(.A(G264), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n449), .A2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n540), .A2(new_n543), .A3(new_n325), .A4(new_n447), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n540), .A2(new_n447), .A3(new_n543), .ZN(new_n545));
  AOI22_X1  g0345(.A1(KEYINPUT85), .A2(new_n544), .B1(new_n545), .B2(new_n409), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n545), .A2(KEYINPUT85), .A3(new_n409), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n525), .B(new_n534), .C1(new_n546), .C2(new_n547), .ZN(new_n548));
  AND3_X1   g0348(.A1(new_n540), .A2(new_n447), .A3(new_n543), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n310), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n545), .A2(new_n308), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n347), .B1(new_n521), .B2(new_n523), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n550), .B(new_n551), .C1(new_n552), .C2(new_n533), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n548), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  AND2_X1   g0355(.A1(KEYINPUT78), .A2(G97), .ZN(new_n556));
  NOR2_X1   g0356(.A1(KEYINPUT78), .A2(G97), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NOR3_X1   g0358(.A1(new_n558), .A2(KEYINPUT19), .A3(new_n348), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n392), .A2(new_n206), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n414), .A2(new_n511), .A3(new_n415), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n560), .B1(new_n561), .B2(new_n481), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n559), .B1(new_n562), .B2(KEYINPUT19), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n269), .A2(new_n206), .A3(G68), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n280), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(G238), .A2(G1698), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n567), .B1(new_n453), .B2(G1698), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n568), .A2(new_n271), .A3(new_n244), .ZN(new_n569));
  NAND2_X1  g0369(.A1(G33), .A2(G116), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n295), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n446), .A2(KEYINPUT80), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n205), .A2(G45), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT80), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n572), .A2(new_n295), .A3(new_n575), .A4(G250), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n295), .A2(G274), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n576), .B1(new_n577), .B2(new_n573), .ZN(new_n578));
  OAI21_X1  g0378(.A(G200), .B1(new_n571), .B2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n431), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n382), .A2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n476), .A2(G87), .ZN(new_n583));
  AND4_X1   g0383(.A1(new_n566), .A2(new_n579), .A3(new_n582), .A4(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(KEYINPUT81), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n571), .A2(new_n578), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(G190), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n566), .A2(new_n579), .A3(new_n582), .A4(new_n583), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT81), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NOR3_X1   g0391(.A1(new_n571), .A2(new_n578), .A3(G179), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n562), .A2(KEYINPUT19), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n564), .B1(new_n593), .B2(new_n559), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n581), .B1(new_n594), .B2(new_n280), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n476), .A2(new_n580), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n592), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n308), .B1(new_n571), .B2(new_n578), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n585), .A2(new_n591), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT21), .ZN(new_n600));
  INV_X1    g0400(.A(G116), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n380), .A2(new_n381), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n601), .B1(new_n205), .B2(G33), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n347), .B(new_n603), .C1(new_n373), .C2(new_n375), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n279), .A2(new_n212), .B1(G20), .B2(new_n601), .ZN(new_n605));
  AOI21_X1  g0405(.A(G33), .B1(new_n479), .B2(new_n480), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n460), .A2(new_n206), .ZN(new_n607));
  OAI211_X1 g0407(.A(KEYINPUT20), .B(new_n605), .C1(new_n606), .C2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n607), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n610), .B1(new_n558), .B2(G33), .ZN(new_n611));
  AOI21_X1  g0411(.A(KEYINPUT20), .B1(new_n611), .B2(new_n605), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n602), .B(new_n604), .C1(new_n609), .C2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(G169), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n448), .A2(G270), .A3(new_n295), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n447), .A2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT82), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n447), .A2(KEYINPUT82), .A3(new_n615), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n541), .A2(G1698), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n620), .B1(G257), .B2(G1698), .ZN(new_n621));
  INV_X1    g0421(.A(G303), .ZN(new_n622));
  OAI22_X1  g0422(.A1(new_n272), .A2(new_n621), .B1(new_n622), .B2(new_n339), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n618), .A2(new_n619), .B1(new_n289), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n600), .B1(new_n614), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n613), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n623), .A2(new_n289), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n447), .A2(KEYINPUT82), .A3(new_n615), .ZN(new_n628));
  AOI21_X1  g0428(.A(KEYINPUT82), .B1(new_n447), .B2(new_n615), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n627), .B(G190), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n626), .B(new_n630), .C1(new_n624), .C2(new_n409), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n632), .A2(KEYINPUT21), .A3(new_n613), .A4(G169), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n624), .A2(new_n613), .A3(G179), .ZN(new_n634));
  AND4_X1   g0434(.A1(new_n625), .A2(new_n631), .A3(new_n633), .A4(new_n634), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n508), .A2(new_n555), .A3(new_n599), .A4(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n442), .A2(new_n636), .ZN(G372));
  OAI21_X1  g0437(.A(new_n313), .B1(new_n308), .B2(new_n307), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n329), .A2(new_n333), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n333), .B1(new_n329), .B2(new_n638), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n405), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n642), .A2(new_n403), .A3(new_n402), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n425), .A2(new_n434), .A3(new_n435), .ZN(new_n644));
  AOI22_X1  g0444(.A1(new_n387), .A2(new_n643), .B1(new_n411), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n330), .A2(new_n332), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n641), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n363), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n648), .A2(new_n365), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n634), .A2(new_n633), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n650), .A2(new_n553), .A3(new_n625), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n598), .A2(KEYINPUT86), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT86), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n653), .B(new_n308), .C1(new_n571), .C2(new_n578), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n597), .A2(new_n655), .B1(new_n584), .B2(new_n587), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n651), .A2(new_n548), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n499), .A2(new_n507), .ZN(new_n658));
  OAI21_X1  g0458(.A(KEYINPUT87), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n584), .A2(new_n587), .ZN(new_n660));
  INV_X1    g0460(.A(new_n592), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n566), .A2(new_n582), .A3(new_n596), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n655), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n548), .A2(new_n660), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT87), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n508), .A2(new_n664), .A3(new_n665), .A4(new_n651), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n659), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n505), .A2(new_n280), .ZN(new_n668));
  AOI22_X1  g0468(.A1(new_n668), .A2(new_n477), .B1(new_n473), .B2(new_n308), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n669), .A2(new_n467), .A3(new_n660), .A4(new_n663), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n663), .B1(new_n670), .B2(KEYINPUT26), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT26), .ZN(new_n672));
  INV_X1    g0472(.A(new_n499), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n672), .B1(new_n599), .B2(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n667), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n441), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n649), .A2(new_n677), .ZN(G369));
  NAND2_X1  g0478(.A1(new_n650), .A2(new_n625), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n355), .A2(new_n206), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(G213), .A3(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(G343), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n626), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n679), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n635), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n688), .B1(new_n689), .B2(new_n687), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(G330), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n686), .B1(new_n525), .B2(new_n534), .ZN(new_n693));
  OAI22_X1  g0493(.A1(new_n554), .A2(new_n693), .B1(new_n553), .B2(new_n686), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n685), .B1(new_n650), .B2(new_n625), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n696), .A2(new_n548), .A3(new_n553), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n553), .A2(new_n685), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n695), .A2(new_n699), .ZN(G399));
  INV_X1    g0500(.A(new_n209), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(G41), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G1), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n416), .A2(new_n511), .A3(new_n601), .A4(new_n558), .ZN(new_n705));
  OAI22_X1  g0505(.A1(new_n704), .A2(new_n705), .B1(new_n215), .B2(new_n703), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT28), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT29), .ZN(new_n708));
  INV_X1    g0508(.A(new_n663), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n709), .B1(new_n670), .B2(KEYINPUT26), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n599), .A2(new_n673), .A3(new_n672), .ZN(new_n711));
  OAI211_X1 g0511(.A(new_n710), .B(new_n711), .C1(new_n658), .C2(new_n657), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n708), .B1(new_n712), .B2(new_n686), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n685), .B1(new_n667), .B2(new_n675), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n713), .B1(new_n714), .B2(new_n708), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(G330), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT31), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n686), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n586), .A2(new_n543), .A3(new_n540), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n721), .A2(new_n632), .A3(new_n310), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(new_n466), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT30), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n722), .A2(KEYINPUT30), .A3(new_n466), .ZN(new_n726));
  AND2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(KEYINPUT89), .B1(new_n466), .B2(new_n549), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT89), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n473), .A2(new_n729), .A3(new_n545), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n586), .A2(KEYINPUT88), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT88), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n732), .B1(new_n571), .B2(new_n578), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n731), .A2(new_n632), .A3(new_n310), .A4(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n728), .A2(new_n730), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n720), .B1(new_n727), .B2(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n635), .A2(new_n499), .A3(new_n507), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n585), .A2(new_n591), .ZN(new_n739));
  INV_X1    g0539(.A(new_n598), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n662), .A2(new_n661), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n738), .A2(new_n742), .A3(new_n554), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n737), .B1(new_n743), .B2(new_n686), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n725), .A2(new_n726), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT90), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n736), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n473), .A2(new_n545), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n734), .B1(new_n748), .B2(KEYINPUT89), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n749), .A2(KEYINPUT90), .A3(new_n730), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n745), .B1(new_n747), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n718), .B1(new_n751), .B2(new_n686), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n717), .B1(new_n744), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n716), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n707), .B1(new_n754), .B2(G1), .ZN(G364));
  NOR2_X1   g0555(.A1(new_n284), .A2(G20), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n205), .B1(new_n756), .B2(G45), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n702), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n206), .A2(new_n310), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G190), .A2(G200), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n760), .ZN(new_n763));
  NOR3_X1   g0563(.A1(new_n763), .A2(new_n325), .A3(G200), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(G58), .ZN(new_n766));
  OAI221_X1 g0566(.A(new_n339), .B1(new_n338), .B2(new_n762), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n206), .A2(G179), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n761), .ZN(new_n769));
  INV_X1    g0569(.A(G159), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT32), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n768), .A2(G190), .A3(G200), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n768), .A2(new_n325), .A3(G200), .ZN(new_n774));
  OAI221_X1 g0574(.A(new_n772), .B1(new_n511), .B2(new_n773), .C1(new_n482), .C2(new_n774), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n760), .A2(G190), .A3(G200), .ZN(new_n776));
  INV_X1    g0576(.A(KEYINPUT93), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n776), .A2(new_n777), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n767), .B(new_n775), .C1(G50), .C2(new_n782), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n310), .A2(new_n409), .A3(G190), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G20), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G97), .ZN(new_n786));
  NOR3_X1   g0586(.A1(new_n763), .A2(new_n409), .A3(G190), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n786), .B1(new_n788), .B2(new_n263), .ZN(new_n789));
  XOR2_X1   g0589(.A(new_n789), .B(KEYINPUT94), .Z(new_n790));
  INV_X1    g0590(.A(G311), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n247), .B1(new_n762), .B2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n785), .ZN(new_n793));
  INV_X1    g0593(.A(G294), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n793), .A2(new_n794), .B1(new_n773), .B2(new_n622), .ZN(new_n795));
  INV_X1    g0595(.A(new_n774), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n792), .B(new_n795), .C1(G283), .C2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(G317), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(KEYINPUT33), .ZN(new_n799));
  OR2_X1    g0599(.A1(new_n798), .A2(KEYINPUT33), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n787), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n769), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G329), .ZN(new_n803));
  INV_X1    g0603(.A(G322), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n801), .B(new_n803), .C1(new_n804), .C2(new_n765), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n805), .B1(G326), .B2(new_n782), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n783), .A2(new_n790), .B1(new_n797), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n206), .B1(KEYINPUT92), .B2(new_n308), .ZN(new_n808));
  OR2_X1    g0608(.A1(new_n308), .A2(KEYINPUT92), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n212), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n759), .B1(new_n807), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(G13), .A2(G33), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(G20), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n810), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n274), .A2(new_n275), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n818), .A2(new_n701), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT91), .ZN(new_n820));
  INV_X1    g0620(.A(new_n215), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(new_n291), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n820), .B(new_n822), .C1(new_n291), .C2(new_n235), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n701), .A2(new_n247), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n824), .A2(G355), .B1(new_n601), .B2(new_n701), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n817), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n812), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT95), .ZN(new_n828));
  INV_X1    g0628(.A(new_n815), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n828), .B1(new_n690), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n692), .A2(new_n759), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(G330), .B2(new_n690), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(G396));
  NAND2_X1  g0634(.A1(new_n434), .A2(new_n685), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n439), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n436), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n644), .A2(new_n686), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n714), .B(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n753), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n759), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n841), .B2(new_n840), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n764), .A2(G143), .ZN(new_n844));
  INV_X1    g0644(.A(new_n762), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n787), .A2(G150), .B1(G159), .B2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(G137), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n844), .B(new_n846), .C1(new_n781), .C2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  AND2_X1   g0649(.A1(new_n849), .A2(KEYINPUT34), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n849), .A2(KEYINPUT34), .ZN(new_n851));
  INV_X1    g0651(.A(new_n818), .ZN(new_n852));
  INV_X1    g0652(.A(G50), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n793), .A2(new_n766), .B1(new_n773), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(G132), .ZN(new_n855));
  OAI22_X1  g0655(.A1(new_n774), .A2(new_n263), .B1(new_n769), .B2(new_n855), .ZN(new_n856));
  OR2_X1    g0656(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NOR4_X1   g0657(.A1(new_n850), .A2(new_n851), .A3(new_n852), .A4(new_n857), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n787), .A2(G283), .B1(G116), .B2(new_n845), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n781), .B2(new_n622), .ZN(new_n860));
  XOR2_X1   g0660(.A(new_n860), .B(KEYINPUT97), .Z(new_n861));
  OAI221_X1 g0661(.A(new_n247), .B1(new_n769), .B2(new_n791), .C1(new_n765), .C2(new_n794), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n796), .A2(G87), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n863), .B(new_n786), .C1(new_n482), .C2(new_n773), .ZN(new_n864));
  NOR3_X1   g0664(.A1(new_n861), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n810), .B1(new_n858), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n759), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n811), .A2(new_n814), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n868), .B(KEYINPUT96), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n867), .B1(new_n870), .B2(new_n338), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n866), .B(new_n871), .C1(new_n839), .C2(new_n814), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n843), .A2(new_n872), .ZN(G384));
  NOR2_X1   g0673(.A1(new_n756), .A2(new_n205), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n743), .A2(new_n686), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n736), .A2(new_n746), .ZN(new_n876));
  AOI21_X1  g0676(.A(KEYINPUT90), .B1(new_n749), .B2(new_n730), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n727), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n719), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n875), .A2(new_n752), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n837), .A2(new_n838), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n408), .A2(new_n410), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n387), .B(new_n685), .C1(new_n643), .C2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n387), .A2(new_n685), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n406), .A2(new_n411), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n881), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n880), .A2(KEYINPUT40), .A3(new_n886), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n683), .B(KEYINPUT99), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n329), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT101), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n330), .A2(new_n891), .A3(new_n332), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n641), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n891), .B1(new_n330), .B2(new_n332), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n890), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n331), .A2(new_n281), .A3(new_n287), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(KEYINPUT100), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT100), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n288), .A2(new_n898), .A3(new_n331), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n329), .B1(new_n638), .B2(new_n888), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n897), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(KEYINPUT37), .ZN(new_n902));
  INV_X1    g0702(.A(new_n316), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n329), .B1(new_n903), .B2(new_n888), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT37), .B1(new_n288), .B2(new_n331), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n902), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n895), .A2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT38), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n242), .B1(new_n277), .B2(new_n263), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n911), .A2(new_n265), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n278), .A2(new_n280), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n287), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n683), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n914), .A2(new_n638), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n916), .A2(new_n917), .A3(new_n896), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(KEYINPUT37), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n906), .ZN(new_n920));
  INV_X1    g0720(.A(new_n916), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n335), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n920), .A2(new_n922), .A3(KEYINPUT38), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n887), .B1(new_n910), .B2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT40), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n406), .A2(new_n411), .A3(new_n884), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n884), .B1(new_n406), .B2(new_n411), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n839), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n743), .A2(new_n686), .B1(new_n878), .B2(new_n719), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n928), .B1(new_n752), .B2(new_n929), .ZN(new_n930));
  AND3_X1   g0730(.A1(new_n920), .A2(new_n922), .A3(KEYINPUT38), .ZN(new_n931));
  AOI21_X1  g0731(.A(KEYINPUT38), .B1(new_n920), .B2(new_n922), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n924), .B1(new_n925), .B2(new_n933), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n441), .A2(new_n880), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n717), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n934), .B2(new_n935), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT39), .ZN(new_n938));
  AOI21_X1  g0738(.A(KEYINPUT38), .B1(new_n895), .B2(new_n907), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n938), .B1(new_n939), .B2(new_n931), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n643), .A2(new_n387), .A3(new_n686), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n335), .A2(new_n921), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n918), .A2(KEYINPUT37), .B1(new_n904), .B2(new_n905), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n909), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n945), .A2(KEYINPUT39), .A3(new_n923), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n940), .A2(new_n942), .A3(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n641), .A2(new_n888), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n926), .A2(new_n927), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n714), .A2(new_n839), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n949), .B1(new_n950), .B2(new_n838), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n945), .A2(new_n923), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n948), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n947), .A2(new_n953), .ZN(new_n954));
  AOI211_X1 g0754(.A(KEYINPUT29), .B(new_n685), .C1(new_n667), .C2(new_n675), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n441), .B1(new_n955), .B2(new_n713), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(new_n649), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n954), .B(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n874), .B1(new_n937), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n958), .B2(new_n937), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n214), .A2(new_n601), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n489), .B(KEYINPUT98), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT35), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n961), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(new_n963), .B2(new_n962), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT36), .Z(new_n966));
  OAI21_X1  g0766(.A(G77), .B1(new_n766), .B2(new_n263), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n215), .A2(new_n967), .B1(G50), .B2(new_n263), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n968), .A2(G1), .A3(new_n284), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n960), .A2(new_n966), .A3(new_n969), .ZN(G367));
  OAI21_X1  g0770(.A(new_n816), .B1(new_n209), .B2(new_n431), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n971), .B1(new_n820), .B2(new_n231), .ZN(new_n972));
  INV_X1    g0772(.A(G150), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n765), .A2(new_n973), .B1(new_n762), .B2(new_n853), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(G137), .B2(new_n802), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n339), .B1(new_n788), .B2(new_n770), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n976), .B1(G77), .B2(new_n796), .ZN(new_n977));
  INV_X1    g0777(.A(new_n773), .ZN(new_n978));
  AOI22_X1  g0778(.A1(new_n978), .A2(G58), .B1(new_n785), .B2(G68), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n782), .A2(G143), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n975), .A2(new_n977), .A3(new_n979), .A4(new_n980), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n852), .B1(new_n798), .B2(new_n769), .C1(new_n558), .C2(new_n774), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT106), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n787), .A2(G294), .B1(G283), .B2(new_n845), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n984), .B1(new_n622), .B2(new_n765), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(new_n496), .B2(new_n785), .ZN(new_n986));
  OAI21_X1  g0786(.A(KEYINPUT105), .B1(new_n773), .B2(new_n601), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT46), .Z(new_n988));
  OAI211_X1 g0788(.A(new_n986), .B(new_n988), .C1(new_n791), .C2(new_n781), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n981), .B1(new_n983), .B2(new_n989), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT47), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n867), .B(new_n972), .C1(new_n991), .C2(new_n810), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n686), .B1(new_n595), .B2(new_n583), .ZN(new_n993));
  MUX2_X1   g0793(.A(new_n656), .B(new_n709), .S(new_n993), .Z(new_n994));
  OAI21_X1  g0794(.A(new_n992), .B1(new_n829), .B2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n697), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n694), .B2(new_n696), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(new_n692), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n754), .A2(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT104), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n499), .B(new_n507), .C1(new_n506), .C2(new_n686), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n499), .B2(new_n686), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n699), .A2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT103), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT45), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n699), .A2(new_n1002), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT44), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1006), .A2(new_n1007), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n695), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1010), .B(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n754), .B1(new_n1000), .B2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n702), .B(KEYINPUT41), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n758), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n994), .B(KEYINPUT43), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1002), .A2(new_n697), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT42), .Z(new_n1018));
  OAI21_X1  g0818(.A(new_n499), .B1(new_n1001), .B2(new_n553), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(new_n686), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1016), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT102), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n994), .A2(KEYINPUT43), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1018), .A2(new_n1020), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1023), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1011), .A2(new_n1002), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1027), .B(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n995), .B1(new_n1015), .B2(new_n1029), .ZN(G387));
  NOR2_X1   g0830(.A1(new_n754), .A2(new_n998), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1031), .A2(new_n703), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1000), .A2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n793), .A2(new_n431), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(G97), .B2(new_n796), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n338), .B2(new_n773), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(G68), .A2(new_n845), .B1(new_n802), .B2(G150), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1037), .B1(new_n765), .B2(new_n853), .C1(new_n282), .C2(new_n788), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n781), .A2(new_n770), .ZN(new_n1039));
  NOR4_X1   g0839(.A1(new_n1036), .A2(new_n1038), .A3(new_n852), .A4(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(G326), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n774), .A2(new_n601), .B1(new_n769), .B2(new_n1041), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(G311), .A2(new_n787), .B1(new_n764), .B2(G317), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1043), .B1(new_n622), .B2(new_n762), .C1(new_n781), .C2(new_n804), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT48), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n978), .A2(G294), .B1(new_n785), .B2(G283), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n818), .B(new_n1042), .C1(new_n1050), .C2(KEYINPUT49), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n1050), .A2(KEYINPUT49), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1040), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n759), .B1(new_n1053), .B2(new_n811), .ZN(new_n1054));
  AOI211_X1 g0854(.A(G45), .B(new_n705), .C1(G68), .C2(G77), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n282), .A2(G50), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT50), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n820), .A2(new_n1058), .ZN(new_n1059));
  OR2_X1    g0859(.A1(new_n1059), .A2(KEYINPUT107), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(KEYINPUT107), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1060), .B(new_n1061), .C1(new_n291), .C2(new_n228), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n824), .A2(new_n705), .B1(new_n482), .B2(new_n701), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n817), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1054), .A2(new_n1064), .ZN(new_n1065));
  OR2_X1    g0865(.A1(new_n694), .A2(new_n829), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n998), .A2(new_n758), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1033), .A2(new_n1067), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n1068), .A2(KEYINPUT108), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1068), .A2(KEYINPUT108), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1069), .A2(new_n1070), .ZN(G393));
  OR2_X1    g0871(.A1(new_n1000), .A2(new_n1012), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1000), .A2(new_n1012), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1072), .A2(new_n702), .A3(new_n1073), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n781), .A2(new_n973), .B1(new_n770), .B2(new_n765), .ZN(new_n1075));
  XOR2_X1   g0875(.A(new_n1075), .B(KEYINPUT51), .Z(new_n1076));
  AOI22_X1  g0876(.A1(new_n787), .A2(G50), .B1(G143), .B2(new_n802), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n282), .B2(new_n762), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n863), .B1(new_n263), .B2(new_n773), .C1(new_n338), .C2(new_n793), .ZN(new_n1079));
  OR4_X1    g0879(.A1(new_n852), .A2(new_n1076), .A3(new_n1078), .A4(new_n1079), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n781), .A2(new_n798), .B1(new_n791), .B2(new_n765), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT52), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n339), .B1(new_n787), .B2(G303), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(G294), .A2(new_n845), .B1(new_n802), .B2(G322), .ZN(new_n1084));
  INV_X1    g0884(.A(G283), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n482), .A2(new_n774), .B1(new_n773), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(G116), .B2(new_n785), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .A4(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n811), .B1(new_n1080), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n820), .A2(new_n238), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n817), .B1(new_n701), .B2(new_n481), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n867), .B(new_n1089), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n829), .B2(new_n1002), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1074), .B(new_n1093), .C1(new_n757), .C2(new_n1012), .ZN(G390));
  NAND2_X1  g0894(.A1(new_n950), .A2(new_n838), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n949), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n753), .B2(new_n839), .ZN(new_n1097));
  AND3_X1   g0897(.A1(new_n880), .A2(G330), .A3(new_n886), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1095), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n880), .A2(G330), .A3(new_n839), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n949), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n753), .A2(new_n839), .A3(new_n1096), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n712), .A2(new_n686), .A3(new_n837), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n838), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1101), .A2(new_n1102), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1099), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n441), .A2(new_n880), .A3(G330), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n649), .B(new_n1108), .C1(new_n715), .C2(new_n442), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n956), .A2(KEYINPUT109), .A3(new_n649), .A4(new_n1108), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1107), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1098), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n940), .A2(new_n946), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n685), .B(new_n881), .C1(new_n667), .C2(new_n675), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n838), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1096), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n941), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1115), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n942), .B1(new_n1104), .B2(new_n1096), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(new_n931), .B2(new_n939), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1114), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n940), .A2(new_n946), .B1(new_n941), .B2(new_n1118), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1122), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1102), .ZN(new_n1126));
  NOR3_X1   g0926(.A1(new_n1124), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1113), .B1(new_n1123), .B2(new_n1127), .ZN(new_n1128));
  AND3_X1   g0928(.A1(new_n1107), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1129));
  NOR3_X1   g0929(.A1(new_n931), .A2(new_n932), .A3(new_n938), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n646), .A2(KEYINPUT101), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1131), .A2(new_n641), .A3(new_n892), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n1132), .A2(new_n890), .B1(new_n906), .B2(new_n902), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n923), .B1(new_n1133), .B2(KEYINPUT38), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1130), .B1(new_n938), .B2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n951), .A2(new_n942), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1122), .B(new_n1102), .C1(new_n1135), .C2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1098), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1129), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1128), .A2(new_n702), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT111), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1138), .A2(new_n1137), .A3(new_n758), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n759), .B1(new_n869), .B2(new_n429), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n788), .A2(new_n416), .B1(new_n762), .B2(new_n558), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(G116), .B2(new_n764), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n247), .B1(new_n769), .B2(new_n794), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(G87), .B2(new_n978), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n796), .A2(G68), .B1(new_n785), .B2(G77), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n782), .A2(G283), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1145), .A2(new_n1147), .A3(new_n1148), .A4(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(G128), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n781), .A2(new_n1151), .B1(new_n855), .B2(new_n765), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT110), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n978), .A2(G150), .ZN(new_n1154));
  XOR2_X1   g0954(.A(new_n1154), .B(KEYINPUT53), .Z(new_n1155));
  XNOR2_X1  g0955(.A(KEYINPUT54), .B(G143), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n247), .B1(new_n845), .B2(new_n1157), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n787), .A2(G137), .B1(G125), .B2(new_n802), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n796), .A2(G50), .B1(new_n785), .B2(G159), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1155), .A2(new_n1158), .A3(new_n1159), .A4(new_n1160), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1150), .B1(new_n1153), .B2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1143), .B1(new_n1162), .B2(new_n810), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(new_n1135), .B2(new_n814), .ZN(new_n1164));
  AND2_X1   g0964(.A1(new_n1142), .A2(new_n1164), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n1140), .A2(new_n1141), .A3(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1141), .B1(new_n1140), .B2(new_n1165), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1166), .A2(new_n1167), .ZN(G378));
  AND2_X1   g0968(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1139), .A2(new_n1169), .ZN(new_n1170));
  AND2_X1   g0970(.A1(new_n947), .A2(new_n953), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n636), .A2(new_n685), .B1(new_n751), .B2(new_n720), .ZN(new_n1172));
  AOI21_X1  g0972(.A(KEYINPUT31), .B1(new_n878), .B2(new_n685), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n886), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(new_n945), .B2(new_n923), .ZN(new_n1175));
  OAI21_X1  g0975(.A(G330), .B1(new_n1175), .B2(KEYINPUT40), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n358), .A2(new_n683), .ZN(new_n1177));
  AND2_X1   g0977(.A1(new_n366), .A2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n366), .A2(new_n1177), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  OR3_X1    g0981(.A1(new_n1178), .A2(new_n1179), .A3(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1181), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NOR3_X1   g0984(.A1(new_n1176), .A2(new_n924), .A3(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1184), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n717), .B1(new_n933), .B2(new_n925), .ZN(new_n1187));
  OAI211_X1 g0987(.A(KEYINPUT40), .B(new_n930), .C1(new_n939), .C2(new_n931), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1186), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1171), .B1(new_n1185), .B2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1184), .B1(new_n1176), .B2(new_n924), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1187), .A2(new_n1188), .A3(new_n1186), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1191), .A2(new_n954), .A3(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1190), .A2(KEYINPUT115), .A3(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT115), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1195), .A2(new_n1196), .A3(new_n1171), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1170), .A2(new_n1194), .A3(KEYINPUT57), .A4(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1193), .A2(KEYINPUT113), .ZN(new_n1199));
  AOI211_X1 g0999(.A(KEYINPUT114), .B(new_n954), .C1(new_n1192), .C2(new_n1191), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT114), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(new_n1195), .B2(new_n1171), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1199), .B1(new_n1200), .B2(new_n1202), .ZN(new_n1203));
  AND2_X1   g1003(.A1(new_n1193), .A2(KEYINPUT113), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1190), .A2(KEYINPUT114), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1195), .A2(new_n1201), .A3(new_n1171), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n1203), .A2(new_n1207), .B1(new_n1169), .B2(new_n1139), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n702), .B(new_n1198), .C1(new_n1208), .C2(KEYINPUT57), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1186), .A2(new_n813), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n759), .B1(new_n869), .B2(G50), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n793), .A2(new_n973), .B1(new_n773), .B2(new_n1156), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(G128), .A2(new_n764), .B1(new_n787), .B2(G132), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1213), .B1(new_n847), .B2(new_n762), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n1212), .B(new_n1214), .C1(G125), .C2(new_n782), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1215), .B(KEYINPUT59), .ZN(new_n1216));
  AOI211_X1 g1016(.A(G33), .B(G41), .C1(new_n802), .C2(G124), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1216), .B(new_n1217), .C1(new_n770), .C2(new_n774), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n290), .B1(new_n263), .B2(new_n793), .C1(new_n788), .C2(new_n485), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n764), .A2(G107), .B1(G283), .B2(new_n802), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1220), .B1(new_n431), .B2(new_n762), .C1(new_n781), .C2(new_n601), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1219), .B(new_n1221), .C1(G77), .C2(new_n978), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n796), .A2(G58), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1223), .B(KEYINPUT112), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1222), .A2(new_n852), .A3(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT58), .ZN(new_n1226));
  OR2_X1    g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n290), .B1(new_n852), .B2(new_n243), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n853), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1218), .A2(new_n1227), .A3(new_n1229), .A4(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1211), .B1(new_n1231), .B2(new_n810), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1210), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1203), .A2(new_n1207), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1234), .B1(new_n1235), .B2(new_n758), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1209), .A2(new_n1236), .ZN(G375));
  NAND2_X1  g1037(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1238), .A2(new_n1099), .A3(new_n1106), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1239), .A2(new_n1014), .A3(new_n1113), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n757), .B(KEYINPUT116), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1107), .A2(new_n1241), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n787), .A2(new_n1157), .B1(G150), .B2(new_n845), .ZN(new_n1243));
  OAI221_X1 g1043(.A(new_n1243), .B1(new_n853), .B2(new_n793), .C1(new_n847), .C2(new_n765), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(G132), .B2(new_n782), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n773), .A2(new_n770), .B1(new_n769), .B2(new_n1151), .ZN(new_n1246));
  XOR2_X1   g1046(.A(new_n1246), .B(KEYINPUT118), .Z(new_n1247));
  NAND4_X1  g1047(.A1(new_n1245), .A2(new_n818), .A3(new_n1224), .A4(new_n1247), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n338), .A2(new_n774), .B1(new_n773), .B2(new_n485), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n339), .B1(new_n845), .B2(new_n496), .ZN(new_n1250));
  OAI221_X1 g1050(.A(new_n1250), .B1(new_n622), .B2(new_n769), .C1(new_n788), .C2(new_n601), .ZN(new_n1251));
  AOI211_X1 g1051(.A(new_n1249), .B(new_n1251), .C1(G294), .C2(new_n782), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1034), .B1(G283), .B2(new_n764), .ZN(new_n1253));
  XOR2_X1   g1053(.A(new_n1253), .B(KEYINPUT117), .Z(new_n1254));
  NAND2_X1  g1054(.A1(new_n1252), .A2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n811), .B1(new_n1248), .B2(new_n1255), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n867), .B(new_n1256), .C1(new_n263), .C2(new_n870), .ZN(new_n1257));
  XOR2_X1   g1057(.A(new_n1257), .B(KEYINPUT119), .Z(new_n1258));
  OAI21_X1  g1058(.A(new_n1258), .B1(new_n814), .B2(new_n1096), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1240), .A2(new_n1242), .A3(new_n1259), .ZN(G381));
  OR2_X1    g1060(.A1(G390), .A2(G387), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1069), .A2(new_n833), .A3(new_n1070), .ZN(new_n1262));
  NOR4_X1   g1062(.A1(new_n1261), .A2(G384), .A3(G381), .A4(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1140), .A2(new_n1165), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1263), .A2(new_n1265), .A3(new_n1209), .A4(new_n1236), .ZN(G407));
  NAND2_X1  g1066(.A1(new_n684), .A2(G213), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1265), .A2(new_n1268), .ZN(new_n1269));
  OAI211_X1 g1069(.A(G407), .B(G213), .C1(G375), .C2(new_n1269), .ZN(G409));
  NOR3_X1   g1070(.A1(new_n1200), .A2(new_n1202), .A3(new_n1199), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(new_n1205), .A2(new_n1206), .B1(KEYINPUT113), .B2(new_n1193), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n1014), .B(new_n1170), .C1(new_n1271), .C2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1194), .A2(new_n1197), .A3(new_n1241), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n1233), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(KEYINPUT120), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT120), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1274), .A2(new_n1277), .A3(new_n1233), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1273), .A2(new_n1276), .A3(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n1265), .ZN(new_n1280));
  AOI21_X1  g1080(.A(KEYINPUT57), .B1(new_n1235), .B2(new_n1170), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1198), .A2(new_n702), .ZN(new_n1282));
  OAI211_X1 g1082(.A(G378), .B(new_n1236), .C1(new_n1281), .C2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1280), .A2(new_n1283), .ZN(new_n1284));
  OR2_X1    g1084(.A1(G384), .A2(KEYINPUT122), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n1285), .A2(new_n1242), .A3(new_n1259), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1113), .A2(KEYINPUT60), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n1239), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(KEYINPUT121), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1169), .A2(new_n1107), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n703), .B1(new_n1290), .B2(KEYINPUT60), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1289), .A2(new_n1291), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1288), .A2(KEYINPUT121), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1286), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(G384), .A2(KEYINPUT122), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1294), .A2(new_n1296), .ZN(new_n1297));
  OAI211_X1 g1097(.A(new_n1295), .B(new_n1286), .C1(new_n1292), .C2(new_n1293), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1284), .A2(new_n1267), .A3(new_n1299), .ZN(new_n1300));
  XNOR2_X1  g1100(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT61), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1268), .B1(new_n1280), .B2(new_n1283), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1268), .A2(G2897), .ZN(new_n1305));
  AND3_X1   g1105(.A1(new_n1297), .A2(new_n1298), .A3(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1305), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1303), .B1(new_n1304), .B2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1310), .B1(new_n1304), .B2(new_n1299), .ZN(new_n1311));
  NOR3_X1   g1111(.A1(new_n1302), .A2(new_n1309), .A3(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT124), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1262), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n833), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1313), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1315), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1317), .A2(new_n1262), .A3(KEYINPUT124), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(G390), .A2(G387), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1316), .A2(new_n1318), .A3(new_n1261), .A4(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(G387), .A2(KEYINPUT125), .ZN(new_n1321));
  OR2_X1    g1121(.A1(new_n1321), .A2(G390), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1317), .A2(new_n1262), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1321), .A2(G390), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1322), .A2(new_n1323), .A3(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1320), .A2(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1308), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1284), .A2(new_n1267), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT123), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1327), .A2(new_n1328), .A3(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT63), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1300), .A2(new_n1331), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1304), .A2(KEYINPUT63), .A3(new_n1299), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1330), .A2(new_n1332), .A3(new_n1333), .ZN(new_n1334));
  OAI21_X1  g1134(.A(KEYINPUT123), .B1(new_n1304), .B2(new_n1308), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1335), .A2(new_n1326), .A3(new_n1303), .ZN(new_n1336));
  OAI22_X1  g1136(.A1(new_n1312), .A2(new_n1326), .B1(new_n1334), .B2(new_n1336), .ZN(G405));
  NAND2_X1  g1137(.A1(G375), .A2(new_n1265), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1338), .A2(KEYINPUT127), .A3(new_n1283), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT127), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1283), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1264), .B1(new_n1209), .B2(new_n1236), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1340), .B1(new_n1341), .B2(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1299), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1339), .A2(new_n1343), .A3(new_n1344), .ZN(new_n1345));
  NAND4_X1  g1145(.A1(new_n1338), .A2(KEYINPUT127), .A3(new_n1283), .A4(new_n1299), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1345), .A2(new_n1346), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1347), .A2(new_n1326), .ZN(new_n1348));
  NAND4_X1  g1148(.A1(new_n1345), .A2(new_n1325), .A3(new_n1320), .A4(new_n1346), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1348), .A2(new_n1349), .ZN(G402));
endmodule


