//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 1 0 0 0 0 0 1 0 0 1 1 0 1 1 0 0 1 0 0 0 1 0 1 0 1 1 0 0 0 0 0 1 1 1 0 1 0 0 1 0 1 1 1 0 1 1 1 0 0 1 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:58 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n748, new_n749, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT13), .A3(G128), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT101), .ZN(new_n194));
  XNOR2_X1  g008(.A(new_n193), .B(new_n194), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n192), .A2(G128), .ZN(new_n196));
  XNOR2_X1  g010(.A(new_n196), .B(KEYINPUT100), .ZN(new_n197));
  INV_X1    g011(.A(G128), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(G143), .ZN(new_n199));
  OAI211_X1 g013(.A(new_n195), .B(new_n197), .C1(KEYINPUT13), .C2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G134), .ZN(new_n201));
  INV_X1    g015(.A(new_n199), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n197), .A2(new_n201), .A3(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT102), .ZN(new_n204));
  AOI22_X1  g018(.A1(new_n200), .A2(G134), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  OR2_X1    g019(.A1(new_n203), .A2(new_n204), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT67), .B(G116), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G122), .ZN(new_n208));
  INV_X1    g022(.A(G107), .ZN(new_n209));
  AND2_X1   g023(.A1(KEYINPUT98), .A2(G122), .ZN(new_n210));
  NOR2_X1   g024(.A1(KEYINPUT98), .A2(G122), .ZN(new_n211));
  OAI21_X1  g025(.A(G116), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n208), .A2(new_n209), .A3(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n209), .B1(new_n208), .B2(new_n212), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT99), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(new_n215), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT99), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n218), .A3(new_n213), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n205), .A2(new_n206), .A3(new_n216), .A4(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n197), .A2(new_n202), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G134), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(new_n203), .ZN(new_n223));
  AND2_X1   g037(.A1(new_n208), .A2(KEYINPUT14), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n212), .B1(new_n208), .B2(KEYINPUT14), .ZN(new_n225));
  OAI21_X1  g039(.A(G107), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n223), .A2(new_n226), .A3(new_n213), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n220), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G217), .ZN(new_n229));
  NOR3_X1   g043(.A1(new_n188), .A2(new_n229), .A3(G953), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n220), .A2(new_n227), .A3(new_n230), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(new_n190), .ZN(new_n235));
  INV_X1    g049(.A(G478), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n236), .A2(KEYINPUT15), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n237), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n234), .A2(new_n190), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT103), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n238), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n239), .B1(new_n234), .B2(new_n190), .ZN(new_n243));
  AOI211_X1 g057(.A(G902), .B(new_n237), .C1(new_n232), .C2(new_n233), .ZN(new_n244));
  OAI21_X1  g058(.A(KEYINPUT103), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G953), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n246), .A2(G952), .ZN(new_n247));
  INV_X1    g061(.A(G234), .ZN(new_n248));
  INV_X1    g062(.A(G237), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  AOI211_X1 g065(.A(new_n190), .B(new_n246), .C1(G234), .C2(G237), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT21), .B(G898), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n242), .A2(new_n245), .A3(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT97), .ZN(new_n257));
  XNOR2_X1  g071(.A(G125), .B(G140), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(KEYINPUT16), .ZN(new_n259));
  INV_X1    g073(.A(G125), .ZN(new_n260));
  OR3_X1    g074(.A1(new_n260), .A2(KEYINPUT16), .A3(G140), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G146), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT77), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n259), .A2(G146), .A3(new_n261), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n262), .A2(KEYINPUT77), .A3(new_n263), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n257), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n249), .A2(new_n246), .A3(G143), .A4(G214), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n272), .A2(KEYINPUT96), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n272), .A2(KEYINPUT96), .ZN(new_n274));
  AND3_X1   g088(.A1(new_n249), .A2(new_n246), .A3(G214), .ZN(new_n275));
  OAI22_X1  g089(.A1(new_n273), .A2(new_n274), .B1(G143), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G131), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n276), .B(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT17), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n276), .A2(KEYINPUT17), .A3(G131), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n266), .A2(KEYINPUT97), .A3(new_n269), .A4(new_n267), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n271), .A2(new_n280), .A3(new_n281), .A4(new_n282), .ZN(new_n283));
  XNOR2_X1  g097(.A(G113), .B(G122), .ZN(new_n284));
  INV_X1    g098(.A(G104), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n284), .B(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n276), .A2(KEYINPUT18), .A3(G131), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n258), .B(new_n263), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT18), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n289), .A2(new_n277), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n287), .B(new_n288), .C1(new_n276), .C2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n283), .A2(new_n286), .A3(new_n291), .ZN(new_n292));
  XOR2_X1   g106(.A(new_n258), .B(KEYINPUT19), .Z(new_n293));
  OAI21_X1  g107(.A(new_n267), .B1(new_n293), .B2(G146), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n291), .B1(new_n278), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n286), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT20), .ZN(new_n299));
  NOR2_X1   g113(.A1(G475), .A2(G902), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n299), .B1(new_n298), .B2(new_n300), .ZN(new_n303));
  INV_X1    g117(.A(G475), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n283), .A2(new_n291), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n296), .ZN(new_n306));
  AOI21_X1  g120(.A(G902), .B1(new_n306), .B2(new_n292), .ZN(new_n307));
  OAI22_X1  g121(.A1(new_n302), .A2(new_n303), .B1(new_n304), .B2(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n256), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT4), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n209), .B(G104), .C1(KEYINPUT83), .C2(KEYINPUT3), .ZN(new_n311));
  NAND2_X1  g125(.A1(KEYINPUT83), .A2(KEYINPUT3), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT84), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n285), .A2(G107), .ZN(new_n315));
  OR2_X1    g129(.A1(KEYINPUT83), .A2(KEYINPUT3), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT84), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n315), .A2(new_n316), .A3(new_n317), .A4(new_n312), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n314), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n285), .A2(KEYINPUT82), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT82), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G104), .ZN(new_n322));
  AND3_X1   g136(.A1(new_n320), .A2(new_n322), .A3(G107), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(KEYINPUT82), .B(G104), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT3), .B1(new_n325), .B2(G107), .ZN(new_n326));
  AND4_X1   g140(.A1(KEYINPUT85), .A2(new_n319), .A3(new_n324), .A4(new_n326), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n321), .A2(G104), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n285), .A2(KEYINPUT82), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n209), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n323), .B1(KEYINPUT3), .B2(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(KEYINPUT85), .B1(new_n331), .B2(new_n319), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n310), .B(G101), .C1(new_n327), .C2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT68), .ZN(new_n334));
  INV_X1    g148(.A(G116), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n335), .A2(G119), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n336), .B1(new_n207), .B2(G119), .ZN(new_n337));
  XOR2_X1   g151(.A(KEYINPUT2), .B(G113), .Z(new_n338));
  AOI21_X1  g152(.A(new_n334), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n335), .A2(KEYINPUT67), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT67), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G116), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n340), .A2(new_n342), .A3(G119), .ZN(new_n343));
  INV_X1    g157(.A(new_n336), .ZN(new_n344));
  AND4_X1   g158(.A1(new_n334), .A2(new_n338), .A3(new_n343), .A4(new_n344), .ZN(new_n345));
  OAI22_X1  g159(.A1(new_n339), .A2(new_n345), .B1(new_n337), .B2(new_n338), .ZN(new_n346));
  INV_X1    g160(.A(G101), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT85), .ZN(new_n348));
  INV_X1    g162(.A(new_n319), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n324), .A2(new_n326), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n348), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n331), .A2(KEYINPUT85), .A3(new_n319), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n347), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n319), .A2(new_n347), .A3(new_n324), .A4(new_n326), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT4), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n333), .B(new_n346), .C1(new_n353), .C2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n337), .A2(KEYINPUT5), .ZN(new_n357));
  OAI211_X1 g171(.A(new_n357), .B(G113), .C1(KEYINPUT5), .C2(new_n344), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n358), .B1(new_n345), .B2(new_n339), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n330), .B1(G104), .B2(new_n209), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G101), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n354), .A2(new_n361), .ZN(new_n362));
  OR2_X1    g176(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n356), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(G110), .B(G122), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n356), .A2(new_n363), .A3(new_n365), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n367), .A2(KEYINPUT6), .A3(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT65), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n370), .B1(new_n263), .B2(G143), .ZN(new_n371));
  OAI21_X1  g185(.A(KEYINPUT64), .B1(new_n192), .B2(G146), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT64), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(new_n263), .A3(G143), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n192), .A2(KEYINPUT65), .A3(G146), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n371), .A2(new_n372), .A3(new_n374), .A4(new_n375), .ZN(new_n376));
  AND2_X1   g190(.A1(KEYINPUT0), .A2(G128), .ZN(new_n377));
  NOR2_X1   g191(.A1(KEYINPUT0), .A2(G128), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n192), .A2(G146), .ZN(new_n380));
  OAI21_X1  g194(.A(KEYINPUT66), .B1(new_n263), .B2(G143), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT66), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(new_n192), .A3(G146), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n380), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  AOI22_X1  g198(.A1(new_n376), .A2(new_n379), .B1(new_n384), .B2(new_n377), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G125), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT1), .ZN(new_n387));
  OAI21_X1  g201(.A(G128), .B1(new_n380), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n376), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n381), .A2(new_n383), .ZN(new_n390));
  INV_X1    g204(.A(new_n380), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n390), .A2(new_n387), .A3(G128), .A4(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n386), .B1(new_n394), .B2(G125), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n246), .A2(G224), .ZN(new_n396));
  XOR2_X1   g210(.A(new_n396), .B(KEYINPUT94), .Z(new_n397));
  XNOR2_X1  g211(.A(new_n395), .B(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT6), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n364), .A2(new_n399), .A3(new_n366), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n369), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n396), .A2(KEYINPUT7), .ZN(new_n402));
  XOR2_X1   g216(.A(new_n395), .B(new_n402), .Z(new_n403));
  INV_X1    g217(.A(KEYINPUT95), .ZN(new_n404));
  OR3_X1    g218(.A1(new_n359), .A2(new_n404), .A3(new_n362), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n404), .B1(new_n359), .B2(new_n362), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n359), .A2(new_n362), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n405), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n365), .B(KEYINPUT8), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n403), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(G902), .B1(new_n410), .B2(new_n368), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n401), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(G210), .B1(G237), .B2(G902), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n401), .A2(new_n413), .A3(new_n411), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(G214), .B1(G237), .B2(G902), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n309), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  XNOR2_X1  g233(.A(G110), .B(G140), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n246), .A2(G227), .ZN(new_n421));
  XOR2_X1   g235(.A(new_n420), .B(new_n421), .Z(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT11), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n424), .B1(new_n201), .B2(G137), .ZN(new_n425));
  INV_X1    g239(.A(G137), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n426), .A2(KEYINPUT11), .A3(G134), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n201), .A2(G137), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n425), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(G131), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n425), .A2(new_n427), .A3(new_n277), .A4(new_n428), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n333), .B(new_n385), .C1(new_n353), .C2(new_n355), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT10), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n435), .B1(new_n389), .B2(new_n392), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n436), .A2(new_n354), .A3(new_n361), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT86), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n436), .A2(new_n354), .A3(KEYINPUT86), .A4(new_n361), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n390), .A2(new_n391), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n388), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n392), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n354), .A2(new_n443), .A3(new_n361), .ZN(new_n444));
  AOI22_X1  g258(.A1(new_n439), .A2(new_n440), .B1(new_n435), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n434), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT91), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT91), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n434), .A2(new_n445), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n433), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  XOR2_X1   g264(.A(new_n432), .B(KEYINPUT87), .Z(new_n451));
  NAND3_X1  g265(.A1(new_n434), .A2(new_n445), .A3(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n423), .B1(new_n450), .B2(new_n453), .ZN(new_n454));
  AND3_X1   g268(.A1(new_n354), .A2(new_n443), .A3(new_n361), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n393), .B1(new_n354), .B2(new_n361), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(KEYINPUT88), .B(KEYINPUT12), .ZN(new_n458));
  NOR3_X1   g272(.A1(new_n457), .A2(new_n433), .A3(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT89), .ZN(new_n460));
  NOR3_X1   g274(.A1(new_n455), .A2(new_n456), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n362), .A2(new_n394), .ZN(new_n462));
  AOI21_X1  g276(.A(KEYINPUT89), .B1(new_n462), .B2(new_n444), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n432), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT12), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n459), .B1(new_n466), .B2(KEYINPUT90), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT90), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n464), .A2(new_n468), .A3(new_n465), .ZN(new_n469));
  AOI21_X1  g283(.A(KEYINPUT93), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n460), .B1(new_n455), .B2(new_n456), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n462), .A2(KEYINPUT89), .A3(new_n444), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n433), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(KEYINPUT90), .B1(new_n473), .B2(KEYINPUT12), .ZN(new_n474));
  INV_X1    g288(.A(new_n459), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n469), .A2(new_n474), .A3(KEYINPUT93), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n452), .A2(new_n422), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n454), .B1(new_n470), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(G469), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n480), .A2(new_n481), .A3(new_n190), .ZN(new_n482));
  INV_X1    g296(.A(new_n449), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n448), .B1(new_n434), .B2(new_n445), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n432), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n478), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n453), .B1(new_n467), .B2(new_n469), .ZN(new_n487));
  OAI211_X1 g301(.A(G469), .B(new_n486), .C1(new_n487), .C2(new_n422), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT92), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n481), .A2(new_n190), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n488), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n447), .A2(new_n449), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n477), .B1(new_n493), .B2(new_n432), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n469), .A2(new_n474), .A3(new_n475), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n452), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n494), .B1(new_n496), .B2(new_n423), .ZN(new_n497));
  OAI211_X1 g311(.A(KEYINPUT92), .B(G469), .C1(new_n497), .C2(G902), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n492), .A2(new_n498), .ZN(new_n499));
  AOI211_X1 g313(.A(new_n191), .B(new_n419), .C1(new_n482), .C2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT81), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT79), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n502), .A2(KEYINPUT25), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT23), .ZN(new_n504));
  INV_X1    g318(.A(G119), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n504), .B1(new_n505), .B2(G128), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n198), .A2(KEYINPUT23), .A3(G119), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n506), .B(new_n507), .C1(G119), .C2(new_n198), .ZN(new_n508));
  XNOR2_X1  g322(.A(G119), .B(G128), .ZN(new_n509));
  XOR2_X1   g323(.A(KEYINPUT24), .B(G110), .Z(new_n510));
  AOI22_X1  g324(.A1(new_n508), .A2(G110), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n511), .B1(new_n268), .B2(new_n270), .ZN(new_n512));
  XOR2_X1   g326(.A(KEYINPUT78), .B(G110), .Z(new_n513));
  OAI22_X1  g327(.A1(new_n508), .A2(new_n513), .B1(new_n509), .B2(new_n510), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n258), .A2(new_n263), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n514), .A2(new_n267), .A3(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(KEYINPUT22), .B(G137), .ZN(new_n517));
  NOR3_X1   g331(.A1(new_n187), .A2(new_n248), .A3(G953), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n517), .B(new_n518), .ZN(new_n519));
  AND3_X1   g333(.A1(new_n512), .A2(new_n516), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n519), .B1(new_n512), .B2(new_n516), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n502), .A2(KEYINPUT25), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n523), .A2(new_n190), .A3(new_n524), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n502), .B(KEYINPUT25), .C1(new_n522), .C2(G902), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n503), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n229), .B1(G234), .B2(new_n190), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n529), .A2(G902), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n530), .B(KEYINPUT80), .ZN(new_n531));
  AOI22_X1  g345(.A1(new_n528), .A2(new_n529), .B1(new_n531), .B2(new_n523), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT31), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n201), .A2(G137), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n426), .A2(G134), .ZN(new_n536));
  OAI21_X1  g350(.A(G131), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n431), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n393), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT69), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n540), .A2(new_n541), .B1(new_n432), .B2(new_n385), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT70), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n346), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n337), .A2(new_n338), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n338), .A2(new_n343), .A3(new_n344), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(KEYINPUT68), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n337), .A2(new_n334), .A3(new_n338), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n545), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT70), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n538), .B1(new_n389), .B2(new_n392), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(KEYINPUT69), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n542), .A2(new_n544), .A3(new_n550), .A4(new_n552), .ZN(new_n553));
  XNOR2_X1  g367(.A(KEYINPUT26), .B(G101), .ZN(new_n554));
  XNOR2_X1  g368(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n554), .B(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n249), .A2(new_n246), .A3(G210), .ZN(new_n557));
  XOR2_X1   g371(.A(new_n557), .B(KEYINPUT72), .Z(new_n558));
  XNOR2_X1  g372(.A(new_n556), .B(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n385), .A2(new_n432), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT30), .ZN(new_n561));
  AND3_X1   g375(.A1(new_n540), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n540), .A2(new_n541), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n563), .A2(new_n552), .A3(new_n560), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n562), .B1(new_n564), .B2(KEYINPUT30), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n553), .B(new_n559), .C1(new_n565), .C2(new_n549), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n534), .B1(new_n566), .B2(KEYINPUT73), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n544), .A2(new_n550), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n568), .A2(new_n564), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n560), .B1(new_n551), .B2(KEYINPUT69), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n393), .A2(KEYINPUT69), .A3(new_n539), .ZN(new_n571));
  OAI21_X1  g385(.A(KEYINPUT30), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n562), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n569), .B1(new_n346), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT73), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n575), .A2(new_n576), .A3(KEYINPUT31), .A4(new_n559), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n567), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n559), .B(KEYINPUT74), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT28), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n540), .A2(new_n560), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n580), .B1(new_n568), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n346), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n580), .B1(new_n553), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT75), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n582), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  AOI211_X1 g400(.A(KEYINPUT75), .B(new_n580), .C1(new_n553), .C2(new_n583), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n579), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(G902), .B1(new_n578), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(G472), .ZN(new_n590));
  AOI21_X1  g404(.A(KEYINPUT32), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n549), .B1(new_n572), .B2(new_n573), .ZN(new_n592));
  INV_X1    g406(.A(new_n559), .ZN(new_n593));
  NOR3_X1   g407(.A1(new_n592), .A2(new_n569), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(KEYINPUT31), .B1(new_n594), .B2(new_n576), .ZN(new_n595));
  NOR3_X1   g409(.A1(new_n566), .A2(KEYINPUT73), .A3(new_n534), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n588), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n597), .A2(KEYINPUT32), .A3(new_n590), .A4(new_n190), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT76), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n589), .A2(KEYINPUT76), .A3(KEYINPUT32), .A4(new_n590), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n591), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n593), .B1(new_n592), .B2(new_n569), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT29), .ZN(new_n604));
  OR2_X1    g418(.A1(new_n584), .A2(new_n585), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n584), .A2(new_n585), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n605), .A2(new_n606), .A3(new_n582), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n603), .B(new_n604), .C1(new_n607), .C2(new_n579), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n568), .A2(new_n564), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n553), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(KEYINPUT28), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n611), .A2(new_n582), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n593), .A2(new_n604), .ZN(new_n613));
  AOI21_X1  g427(.A(G902), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n590), .B1(new_n608), .B2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  AOI211_X1 g430(.A(new_n501), .B(new_n533), .C1(new_n602), .C2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n600), .A2(new_n601), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n589), .A2(new_n590), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT32), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n618), .A2(new_n616), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(KEYINPUT81), .B1(new_n622), .B2(new_n532), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n500), .B1(new_n617), .B2(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G101), .ZN(G3));
  AOI22_X1  g439(.A1(new_n607), .A2(new_n579), .B1(new_n567), .B2(new_n577), .ZN(new_n626));
  OAI21_X1  g440(.A(KEYINPUT104), .B1(new_n626), .B2(G902), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT104), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n589), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT105), .ZN(new_n631));
  AOI22_X1  g445(.A1(new_n630), .A2(G472), .B1(new_n631), .B2(new_n619), .ZN(new_n632));
  AOI211_X1 g446(.A(KEYINPUT105), .B(new_n590), .C1(new_n627), .C2(new_n629), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n191), .B1(new_n499), .B2(new_n482), .ZN(new_n635));
  AND3_X1   g449(.A1(new_n634), .A2(new_n532), .A3(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT106), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n416), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n401), .A2(KEYINPUT106), .A3(new_n413), .A4(new_n411), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n638), .A2(new_n415), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n418), .ZN(new_n641));
  INV_X1    g455(.A(new_n303), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n306), .A2(new_n292), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n190), .ZN(new_n644));
  AOI22_X1  g458(.A1(new_n642), .A2(new_n301), .B1(new_n644), .B2(G475), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n234), .A2(KEYINPUT33), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT33), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n647), .B1(new_n232), .B2(new_n233), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n190), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(G478), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n235), .A2(G478), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NOR4_X1   g467(.A1(new_n641), .A2(new_n645), .A3(new_n254), .A4(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n636), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT34), .B(G104), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G6));
  INV_X1    g471(.A(KEYINPUT107), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n301), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(new_n303), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n644), .A2(G475), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n241), .B1(new_n238), .B2(new_n240), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n243), .A2(new_n244), .A3(KEYINPUT103), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  OR2_X1    g478(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n665), .A2(new_n641), .A3(new_n254), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n636), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT35), .B(G107), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G9));
  INV_X1    g483(.A(new_n419), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n512), .A2(new_n516), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n519), .A2(KEYINPUT36), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n531), .ZN(new_n674));
  INV_X1    g488(.A(new_n529), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n674), .B1(new_n527), .B2(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n634), .A2(new_n635), .A3(new_n670), .A4(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(KEYINPUT108), .ZN(new_n678));
  XNOR2_X1  g492(.A(KEYINPUT37), .B(G110), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G12));
  INV_X1    g494(.A(new_n676), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n681), .B1(new_n602), .B2(new_n616), .ZN(new_n682));
  INV_X1    g496(.A(new_n641), .ZN(new_n683));
  INV_X1    g497(.A(G900), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n252), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n250), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n665), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n682), .A2(new_n635), .A3(new_n683), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G128), .ZN(G30));
  XNOR2_X1  g504(.A(new_n686), .B(KEYINPUT39), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n635), .A2(new_n691), .ZN(new_n692));
  OR2_X1    g506(.A1(new_n692), .A2(KEYINPUT40), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(KEYINPUT40), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n594), .B1(new_n579), .B2(new_n610), .ZN(new_n695));
  OAI21_X1  g509(.A(G472), .B1(new_n695), .B2(G902), .ZN(new_n696));
  AND2_X1   g510(.A1(new_n602), .A2(new_n696), .ZN(new_n697));
  XOR2_X1   g511(.A(KEYINPUT109), .B(KEYINPUT38), .Z(new_n698));
  XNOR2_X1  g512(.A(new_n417), .B(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n662), .A2(new_n663), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n700), .A2(new_n645), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n681), .A2(new_n418), .ZN(new_n703));
  NOR4_X1   g517(.A1(new_n697), .A2(new_n699), .A3(new_n702), .A4(new_n703), .ZN(new_n704));
  AND3_X1   g518(.A1(new_n693), .A2(new_n694), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(new_n192), .ZN(G45));
  AOI21_X1  g520(.A(new_n651), .B1(new_n649), .B2(G478), .ZN(new_n707));
  AND3_X1   g521(.A1(new_n308), .A2(new_n707), .A3(new_n686), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n682), .A2(new_n635), .A3(new_n683), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G146), .ZN(G48));
  AOI21_X1  g524(.A(new_n422), .B1(new_n485), .B2(new_n452), .ZN(new_n711));
  AND2_X1   g525(.A1(new_n476), .A2(new_n478), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT93), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n495), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n711), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g529(.A(G469), .B1(new_n715), .B2(G902), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT110), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n716), .A2(new_n717), .A3(new_n482), .ZN(new_n718));
  OAI211_X1 g532(.A(KEYINPUT110), .B(G469), .C1(new_n715), .C2(G902), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n191), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n533), .B1(new_n602), .B2(new_n616), .ZN(new_n721));
  AND2_X1   g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AND2_X1   g536(.A1(new_n722), .A2(new_n654), .ZN(new_n723));
  XOR2_X1   g537(.A(KEYINPUT41), .B(G113), .Z(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(G15));
  AND2_X1   g539(.A1(new_n722), .A2(new_n666), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(new_n335), .ZN(G18));
  NAND4_X1  g541(.A1(new_n720), .A2(new_n309), .A3(new_n683), .A4(new_n682), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G119), .ZN(G21));
  NAND3_X1  g543(.A1(new_n640), .A2(new_n701), .A3(new_n418), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT111), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n640), .A2(new_n701), .A3(KEYINPUT111), .A4(new_n418), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g548(.A(G472), .B1(new_n626), .B2(G902), .ZN(new_n735));
  INV_X1    g549(.A(new_n579), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n578), .B1(new_n736), .B2(new_n612), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n737), .A2(new_n590), .A3(new_n190), .ZN(new_n738));
  AND2_X1   g552(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n532), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(new_n254), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n734), .A2(new_n720), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(KEYINPUT112), .B(G122), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n742), .B(new_n743), .ZN(G24));
  NAND2_X1  g558(.A1(new_n718), .A2(new_n719), .ZN(new_n745));
  INV_X1    g559(.A(new_n191), .ZN(new_n746));
  AND4_X1   g560(.A1(new_n676), .A2(new_n708), .A3(new_n735), .A4(new_n738), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n745), .A2(new_n746), .A3(new_n683), .A4(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(KEYINPUT113), .B(G125), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n748), .B(new_n749), .ZN(G27));
  INV_X1    g564(.A(new_n418), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n417), .A2(new_n191), .A3(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n490), .B1(new_n497), .B2(G469), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n482), .A2(new_n753), .A3(KEYINPUT114), .ZN(new_n754));
  AOI21_X1  g568(.A(KEYINPUT114), .B1(new_n482), .B2(new_n753), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n708), .B(new_n752), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT115), .ZN(new_n757));
  OAI211_X1 g571(.A(new_n616), .B(new_n598), .C1(new_n621), .C2(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n591), .A2(KEYINPUT115), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n532), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g574(.A(KEYINPUT42), .B1(new_n756), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n482), .A2(new_n753), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT114), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n482), .A2(new_n753), .A3(KEYINPUT114), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR4_X1   g580(.A1(new_n653), .A2(new_n645), .A3(KEYINPUT42), .A4(new_n687), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n766), .A2(new_n721), .A3(new_n752), .A4(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n761), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(new_n277), .ZN(G33));
  NAND4_X1  g584(.A1(new_n766), .A2(new_n721), .A3(new_n688), .A4(new_n752), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G134), .ZN(G36));
  NOR2_X1   g586(.A1(new_n417), .A2(new_n751), .ZN(new_n773));
  INV_X1    g587(.A(new_n634), .ZN(new_n774));
  OAI21_X1  g588(.A(KEYINPUT43), .B1(new_n653), .B2(new_n308), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT43), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n645), .A2(new_n776), .A3(new_n707), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n774), .A2(new_n676), .A3(new_n775), .A4(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT44), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n773), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n780), .B1(new_n779), .B2(new_n778), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT117), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT45), .ZN(new_n783));
  AOI211_X1 g597(.A(new_n783), .B(new_n494), .C1(new_n423), .C2(new_n496), .ZN(new_n784));
  OAI21_X1  g598(.A(G469), .B1(new_n497), .B2(KEYINPUT45), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n784), .B1(new_n785), .B2(KEYINPUT116), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT116), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n787), .B(G469), .C1(new_n497), .C2(KEYINPUT45), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n782), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(KEYINPUT45), .A2(G469), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n488), .A2(KEYINPUT116), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n497), .A2(KEYINPUT45), .ZN(new_n792));
  AND4_X1   g606(.A1(new_n782), .A2(new_n791), .A3(new_n788), .A4(new_n792), .ZN(new_n793));
  OAI211_X1 g607(.A(KEYINPUT46), .B(new_n491), .C1(new_n789), .C2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n482), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n786), .A2(new_n782), .A3(new_n788), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n791), .A2(new_n788), .A3(new_n792), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(KEYINPUT117), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(KEYINPUT46), .B1(new_n799), .B2(new_n491), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n746), .B1(new_n795), .B2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n691), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n781), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G137), .ZN(G39));
  AOI211_X1 g619(.A(new_n615), .B(new_n591), .C1(new_n600), .C2(new_n601), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n806), .A2(new_n533), .A3(new_n708), .A4(new_n773), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT47), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n801), .A2(new_n808), .ZN(new_n809));
  OAI211_X1 g623(.A(KEYINPUT47), .B(new_n746), .C1(new_n795), .C2(new_n800), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n807), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  XOR2_X1   g625(.A(new_n811), .B(G140), .Z(G42));
  NOR2_X1   g626(.A1(G952), .A2(G953), .ZN(new_n813));
  XOR2_X1   g627(.A(new_n813), .B(KEYINPUT123), .Z(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT121), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n745), .A2(new_n191), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n809), .A2(new_n810), .A3(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n775), .A2(new_n251), .A3(new_n777), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n740), .A2(new_n819), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n820), .A2(new_n773), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n816), .B1(new_n818), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n745), .A2(new_n752), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n602), .A2(new_n696), .ZN(new_n824));
  NOR4_X1   g638(.A1(new_n823), .A2(new_n533), .A3(new_n250), .A4(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n825), .A2(new_n645), .A3(new_n653), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n823), .A2(new_n819), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n739), .A2(new_n676), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n820), .A2(new_n751), .A3(new_n699), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n830), .A2(KEYINPUT50), .A3(new_n720), .ZN(new_n831));
  AOI21_X1  g645(.A(KEYINPUT50), .B1(new_n830), .B2(new_n720), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n826), .B(new_n829), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n833), .B1(new_n818), .B2(new_n821), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n822), .A2(new_n834), .A3(KEYINPUT51), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n836));
  AOI221_X4 g650(.A(new_n833), .B1(new_n816), .B2(new_n836), .C1(new_n818), .C2(new_n821), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n825), .A2(new_n308), .A3(new_n707), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n720), .A2(new_n683), .A3(new_n820), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n838), .A2(new_n247), .A3(new_n839), .ZN(new_n840));
  OR2_X1    g654(.A1(new_n840), .A2(KEYINPUT122), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(KEYINPUT122), .ZN(new_n842));
  INV_X1    g656(.A(new_n760), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n827), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(KEYINPUT48), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n841), .A2(new_n842), .A3(new_n845), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n835), .A2(new_n837), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n238), .A2(new_n240), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n661), .B(new_n848), .C1(new_n303), .C2(new_n302), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n849), .B1(new_n645), .B2(new_n653), .ZN(new_n850));
  AND4_X1   g664(.A1(new_n255), .A2(new_n850), .A3(new_n418), .A4(new_n417), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n634), .A2(new_n635), .A3(new_n532), .A4(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n677), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n499), .A2(new_n482), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n854), .A2(new_n670), .A3(new_n746), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n501), .B1(new_n806), .B2(new_n533), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n622), .A2(KEYINPUT81), .A3(new_n532), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n855), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(KEYINPUT118), .B1(new_n853), .B2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT118), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n624), .A2(new_n860), .A3(new_n677), .A4(new_n852), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n720), .B(new_n721), .C1(new_n654), .C2(new_n666), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n863), .A2(new_n728), .A3(new_n742), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n766), .A2(new_n708), .A3(new_n828), .A4(new_n752), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n848), .A2(new_n687), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n676), .A2(new_n661), .A3(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n867), .A2(new_n660), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n635), .A2(new_n622), .A3(new_n773), .A4(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n771), .A2(new_n865), .A3(new_n869), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n864), .A2(new_n769), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n734), .A2(new_n824), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT119), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n681), .A2(new_n746), .A3(new_n686), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n766), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n875), .B1(new_n754), .B2(new_n755), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(KEYINPUT119), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n872), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n689), .A2(new_n709), .A3(new_n748), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT52), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n689), .A2(new_n709), .A3(new_n748), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n697), .B1(new_n732), .B2(new_n733), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n873), .B1(new_n766), .B2(new_n875), .ZN(new_n885));
  AOI211_X1 g699(.A(KEYINPUT119), .B(new_n874), .C1(new_n764), .C2(new_n765), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n884), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT52), .B1(new_n883), .B2(new_n887), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n862), .B(new_n871), .C1(new_n882), .C2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT53), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT54), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n881), .B1(new_n879), .B2(new_n880), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n883), .A2(KEYINPUT52), .A3(new_n887), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n895), .A2(KEYINPUT53), .A3(new_n862), .A4(new_n871), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n891), .A2(new_n892), .A3(new_n896), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n862), .A2(new_n871), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n898), .A2(KEYINPUT120), .A3(KEYINPUT53), .A4(new_n895), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT120), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n896), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n899), .A2(new_n901), .A3(new_n891), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n897), .B1(KEYINPUT54), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n815), .B1(new_n847), .B2(new_n903), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n745), .B(KEYINPUT49), .Z(new_n905));
  NAND3_X1  g719(.A1(new_n532), .A2(new_n746), .A3(new_n418), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n906), .A2(new_n308), .A3(new_n653), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n699), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n905), .A2(new_n824), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(KEYINPUT124), .B1(new_n904), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n902), .A2(KEYINPUT54), .ZN(new_n911));
  INV_X1    g725(.A(new_n897), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n818), .A2(new_n821), .ZN(new_n914));
  AOI21_X1  g728(.A(KEYINPUT51), .B1(new_n914), .B2(KEYINPUT121), .ZN(new_n915));
  INV_X1    g729(.A(new_n834), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n846), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(new_n837), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n814), .B1(new_n913), .B2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT124), .ZN(new_n921));
  INV_X1    g735(.A(new_n909), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n910), .A2(new_n923), .ZN(G75));
  AND2_X1   g738(.A1(new_n891), .A2(new_n896), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n925), .A2(new_n190), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(G210), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT56), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n369), .A2(new_n400), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(new_n398), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT55), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n927), .A2(new_n928), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n931), .B1(new_n927), .B2(new_n928), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n246), .A2(G952), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(G51));
  XNOR2_X1  g749(.A(new_n490), .B(KEYINPUT57), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n925), .A2(new_n892), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n936), .B1(new_n937), .B2(new_n897), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n480), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n926), .A2(new_n796), .A3(new_n798), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n934), .B1(new_n939), .B2(new_n940), .ZN(G54));
  NAND3_X1  g755(.A1(new_n926), .A2(KEYINPUT58), .A3(G475), .ZN(new_n942));
  INV_X1    g756(.A(new_n298), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n942), .A2(new_n943), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n944), .A2(new_n945), .A3(new_n934), .ZN(G60));
  NOR2_X1   g760(.A1(new_n646), .A2(new_n648), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(G478), .A2(G902), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT59), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n948), .B(new_n950), .C1(new_n937), .C2(new_n897), .ZN(new_n951));
  INV_X1    g765(.A(new_n934), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n948), .B1(new_n913), .B2(new_n950), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n953), .A2(new_n954), .ZN(G63));
  NAND2_X1  g769(.A1(G217), .A2(G902), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT60), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n925), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n673), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n522), .B1(new_n925), .B2(new_n957), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n959), .A2(new_n952), .A3(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT61), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n961), .B(new_n962), .ZN(G66));
  INV_X1    g777(.A(G224), .ZN(new_n964));
  NOR3_X1   g778(.A1(new_n253), .A2(new_n964), .A3(new_n246), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n864), .B1(new_n859), .B2(new_n861), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n965), .B1(new_n966), .B2(new_n246), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n929), .B1(G898), .B2(new_n246), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n967), .B(new_n968), .ZN(G69));
  NAND3_X1  g783(.A1(new_n803), .A2(new_n734), .A3(new_n843), .ZN(new_n970));
  INV_X1    g784(.A(new_n771), .ZN(new_n971));
  NOR3_X1   g785(.A1(new_n769), .A2(new_n880), .A3(new_n971), .ZN(new_n972));
  AND3_X1   g786(.A1(new_n970), .A2(new_n804), .A3(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(new_n811), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n973), .A2(new_n246), .A3(new_n974), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n574), .B(new_n293), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n976), .B1(G900), .B2(G953), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n850), .B(KEYINPUT126), .Z(new_n979));
  NOR4_X1   g793(.A1(new_n692), .A2(new_n979), .A3(new_n751), .A4(new_n417), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n980), .B1(new_n623), .B2(new_n617), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n804), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n705), .A2(new_n880), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT62), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n982), .A2(new_n984), .A3(new_n974), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT127), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n982), .A2(new_n984), .A3(KEYINPUT127), .A4(new_n974), .ZN(new_n988));
  AOI21_X1  g802(.A(G953), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n976), .B(KEYINPUT125), .Z(new_n990));
  OAI21_X1  g804(.A(new_n978), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n246), .B1(G227), .B2(G900), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(new_n992), .ZN(new_n994));
  OAI211_X1 g808(.A(new_n994), .B(new_n978), .C1(new_n989), .C2(new_n990), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n993), .A2(new_n995), .ZN(G72));
  NAND3_X1  g810(.A1(new_n987), .A2(new_n966), .A3(new_n988), .ZN(new_n997));
  NAND2_X1  g811(.A1(G472), .A2(G902), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n998), .B(KEYINPUT63), .Z(new_n999));
  AOI211_X1 g813(.A(new_n593), .B(new_n575), .C1(new_n997), .C2(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n603), .A2(new_n566), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n902), .A2(new_n999), .A3(new_n1001), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n973), .A2(new_n974), .A3(new_n966), .ZN(new_n1003));
  AND2_X1   g817(.A1(new_n1003), .A2(new_n999), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n575), .A2(new_n593), .ZN(new_n1005));
  OAI211_X1 g819(.A(new_n952), .B(new_n1002), .C1(new_n1004), .C2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n1000), .A2(new_n1006), .ZN(G57));
endmodule


