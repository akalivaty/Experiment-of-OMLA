//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 1 0 1 0 0 1 1 1 1 0 0 0 0 0 1 1 0 0 0 1 1 1 0 0 0 1 1 0 1 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:47 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1190, new_n1191, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(G13), .ZN(new_n209));
  NAND3_X1  g0009(.A1(new_n208), .A2(KEYINPUT64), .A3(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  AOI21_X1  g0011(.A(KEYINPUT64), .B1(new_n208), .B2(new_n209), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XOR2_X1   g0015(.A(new_n215), .B(KEYINPUT0), .Z(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n217));
  INV_X1    g0017(.A(G116), .ZN(new_n218));
  INV_X1    g0018(.A(G270), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G97), .A2(G257), .ZN(new_n222));
  INV_X1    g0022(.A(G68), .ZN(new_n223));
  INV_X1    g0023(.A(G238), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n221), .B(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI211_X1 g0025(.A(new_n220), .B(new_n225), .C1(G58), .C2(G232), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n226), .A2(new_n208), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT1), .Z(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n229), .A2(new_n207), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT65), .Z(new_n231));
  INV_X1    g0031(.A(new_n201), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(G50), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  AOI211_X1 g0034(.A(new_n216), .B(new_n228), .C1(new_n231), .C2(new_n234), .ZN(G361));
  XOR2_X1   g0035(.A(G238), .B(G244), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT2), .ZN(new_n238));
  INV_X1    g0038(.A(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G264), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(new_n219), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT66), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n240), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(G107), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(new_n218), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G351));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n229), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT67), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n206), .A2(G20), .ZN(new_n259));
  OAI211_X1 g0059(.A(new_n258), .B(new_n259), .C1(new_n257), .C2(new_n255), .ZN(new_n260));
  OR2_X1    g0060(.A1(new_n260), .A2(new_n202), .ZN(new_n261));
  INV_X1    g0061(.A(new_n256), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(new_n202), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n203), .A2(G20), .ZN(new_n264));
  INV_X1    g0064(.A(G150), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G20), .A2(G33), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT8), .B(G58), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n207), .A2(G33), .ZN(new_n269));
  OAI221_X1 g0069(.A(new_n264), .B1(new_n265), .B2(new_n267), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n254), .ZN(new_n271));
  AND3_X1   g0071(.A1(new_n261), .A2(new_n263), .A3(new_n271), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT3), .B(G33), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n273), .A2(G223), .A3(G1698), .ZN(new_n274));
  INV_X1    g0074(.A(G77), .ZN(new_n275));
  INV_X1    g0075(.A(G1698), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G222), .ZN(new_n278));
  OAI221_X1 g0078(.A(new_n274), .B1(new_n275), .B2(new_n273), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G33), .ZN(new_n280));
  INV_X1    g0080(.A(G41), .ZN(new_n281));
  OAI211_X1 g0081(.A(G1), .B(G13), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n285));
  INV_X1    g0085(.A(G274), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  AND2_X1   g0088(.A1(new_n282), .A2(new_n285), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G226), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n284), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n272), .A2(KEYINPUT9), .B1(new_n291), .B2(G200), .ZN(new_n292));
  INV_X1    g0092(.A(G190), .ZN(new_n293));
  OAI221_X1 g0093(.A(new_n292), .B1(KEYINPUT9), .B2(new_n272), .C1(new_n293), .C2(new_n291), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n294), .B(KEYINPUT10), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n273), .A2(G232), .A3(G1698), .ZN(new_n296));
  NAND2_X1  g0096(.A1(G33), .A2(G97), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n296), .B(new_n297), .C1(new_n277), .C2(new_n239), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n287), .B1(new_n298), .B2(new_n283), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT13), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n289), .A2(G238), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n300), .B1(new_n299), .B2(new_n301), .ZN(new_n304));
  OR3_X1    g0104(.A1(new_n303), .A2(new_n293), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n223), .A2(G20), .ZN(new_n306));
  OAI221_X1 g0106(.A(new_n306), .B1(new_n269), .B2(new_n275), .C1(new_n267), .C2(new_n202), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n307), .A2(KEYINPUT11), .A3(new_n254), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n255), .A2(new_n259), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n308), .B1(new_n223), .B2(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n256), .A2(G68), .ZN(new_n311));
  XNOR2_X1  g0111(.A(new_n311), .B(KEYINPUT12), .ZN(new_n312));
  AOI21_X1  g0112(.A(KEYINPUT11), .B1(new_n307), .B2(new_n254), .ZN(new_n313));
  NOR3_X1   g0113(.A1(new_n310), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(G200), .B1(new_n303), .B2(new_n304), .ZN(new_n315));
  AND3_X1   g0115(.A1(new_n305), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n303), .A2(new_n304), .ZN(new_n317));
  INV_X1    g0117(.A(G169), .ZN(new_n318));
  OAI21_X1  g0118(.A(KEYINPUT14), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n317), .A2(G179), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT14), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n321), .B(G169), .C1(new_n303), .C2(new_n304), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n319), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n314), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n316), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n272), .ZN(new_n326));
  INV_X1    g0126(.A(new_n291), .ZN(new_n327));
  INV_X1    g0127(.A(G179), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n326), .B(new_n329), .C1(G169), .C2(new_n327), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n273), .A2(G238), .A3(G1698), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n273), .A2(G232), .A3(new_n276), .ZN(new_n332));
  INV_X1    g0132(.A(G107), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n331), .B(new_n332), .C1(new_n333), .C2(new_n273), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n283), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n289), .A2(G244), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n335), .A2(new_n288), .A3(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n328), .ZN(new_n339));
  INV_X1    g0139(.A(new_n268), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n340), .A2(new_n266), .B1(G20), .B2(G77), .ZN(new_n341));
  XOR2_X1   g0141(.A(KEYINPUT15), .B(G87), .Z(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n341), .B1(new_n269), .B2(new_n343), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n344), .A2(new_n254), .B1(new_n275), .B2(new_n262), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n345), .B1(new_n275), .B2(new_n309), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n337), .A2(new_n318), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n339), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n295), .A2(new_n325), .A3(new_n330), .A4(new_n348), .ZN(new_n349));
  AND2_X1   g0149(.A1(KEYINPUT3), .A2(G33), .ZN(new_n350));
  NOR2_X1   g0150(.A1(KEYINPUT3), .A2(G33), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(KEYINPUT7), .B1(new_n352), .B2(new_n207), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT3), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n280), .ZN(new_n355));
  NAND2_X1  g0155(.A1(KEYINPUT3), .A2(G33), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n355), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(G68), .B1(new_n353), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G159), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n267), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(G58), .A2(G68), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n207), .B1(new_n232), .B2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n359), .A2(new_n362), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(KEYINPUT16), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n355), .A2(new_n207), .A3(new_n356), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT7), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n357), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n364), .B1(new_n371), .B2(G68), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT16), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n372), .A2(new_n373), .A3(new_n362), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n255), .B1(new_n367), .B2(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n340), .A2(new_n256), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n260), .A2(new_n268), .ZN(new_n377));
  NOR3_X1   g0177(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n282), .A2(G232), .A3(new_n285), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT69), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n282), .A2(KEYINPUT69), .A3(G232), .A4(new_n285), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n381), .A2(new_n288), .A3(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n273), .A2(G226), .A3(G1698), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n273), .A2(G223), .A3(new_n276), .ZN(new_n386));
  NAND3_X1  g0186(.A1(KEYINPUT68), .A2(G33), .A3(G87), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT68), .ZN(new_n388));
  INV_X1    g0188(.A(G87), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n388), .B1(new_n280), .B2(new_n389), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n385), .A2(new_n386), .A3(new_n387), .A4(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n283), .ZN(new_n392));
  AOI21_X1  g0192(.A(G200), .B1(new_n384), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n383), .A2(KEYINPUT70), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT70), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n381), .A2(new_n395), .A3(new_n288), .A4(new_n382), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n394), .A2(new_n396), .B1(new_n283), .B2(new_n391), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n393), .B1(new_n397), .B2(new_n293), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n378), .A2(new_n399), .A3(KEYINPUT71), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n373), .B1(new_n372), .B2(new_n362), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n223), .B1(new_n370), .B2(new_n357), .ZN(new_n402));
  NOR4_X1   g0202(.A1(new_n402), .A2(KEYINPUT16), .A3(new_n361), .A4(new_n364), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n254), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n376), .ZN(new_n405));
  INV_X1    g0205(.A(new_n377), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT72), .ZN(new_n408));
  NOR3_X1   g0208(.A1(new_n407), .A2(new_n398), .A3(new_n408), .ZN(new_n409));
  OAI211_X1 g0209(.A(KEYINPUT17), .B(new_n400), .C1(new_n409), .C2(KEYINPUT71), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n384), .A2(new_n392), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n318), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n397), .A2(new_n328), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n407), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT18), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n407), .A2(KEYINPUT18), .A3(new_n412), .A4(new_n413), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT71), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT17), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n378), .A2(new_n399), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n419), .B(new_n420), .C1(new_n421), .C2(new_n408), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n410), .A2(new_n418), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n346), .B1(G200), .B2(new_n337), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n338), .A2(G190), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  NOR3_X1   g0227(.A1(new_n349), .A2(new_n423), .A3(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT19), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n207), .B1(new_n297), .B2(new_n429), .ZN(new_n430));
  NOR2_X1   g0230(.A1(G97), .A2(G107), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n389), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n207), .A2(G33), .A3(G97), .ZN(new_n433));
  AOI22_X1  g0233(.A1(new_n430), .A2(new_n432), .B1(new_n429), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n273), .A2(new_n207), .A3(G68), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n254), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n342), .A2(new_n256), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n206), .A2(G33), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n255), .A2(new_n256), .A3(new_n440), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n437), .B(new_n439), .C1(new_n343), .C2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT78), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n255), .B1(new_n434), .B2(new_n435), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n441), .A2(new_n343), .ZN(new_n446));
  NOR3_X1   g0246(.A1(new_n445), .A2(new_n446), .A3(new_n438), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(KEYINPUT78), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n444), .A2(new_n448), .ZN(new_n449));
  OAI211_X1 g0249(.A(G244), .B(G1698), .C1(new_n350), .C2(new_n351), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT77), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT77), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n273), .A2(new_n452), .A3(G244), .A4(G1698), .ZN(new_n453));
  NAND2_X1  g0253(.A1(G33), .A2(G116), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n273), .A2(G238), .A3(new_n276), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n451), .A2(new_n453), .A3(new_n454), .A4(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n283), .ZN(new_n457));
  INV_X1    g0257(.A(G45), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n458), .A2(G1), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n282), .A2(new_n460), .A3(G250), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n461), .B1(new_n286), .B2(new_n460), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n457), .A2(new_n328), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n462), .B1(new_n456), .B2(new_n283), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n464), .B1(G169), .B2(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n441), .A2(new_n389), .ZN(new_n467));
  NOR3_X1   g0267(.A1(new_n445), .A2(new_n467), .A3(new_n438), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n457), .A2(new_n463), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n468), .B1(new_n469), .B2(new_n293), .ZN(new_n470));
  INV_X1    g0270(.A(G200), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n465), .A2(new_n471), .ZN(new_n472));
  OAI22_X1  g0272(.A1(new_n449), .A2(new_n466), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT5), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT74), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n474), .B1(new_n475), .B2(G41), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n281), .A2(KEYINPUT74), .A3(KEYINPUT5), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n476), .A2(new_n477), .A3(new_n459), .A4(G274), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n273), .A2(G257), .A3(new_n276), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n352), .A2(G303), .ZN(new_n481));
  OAI211_X1 g0281(.A(G264), .B(G1698), .C1(new_n350), .C2(new_n351), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n479), .B1(new_n483), .B2(new_n283), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n476), .A2(new_n477), .A3(new_n459), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n485), .A2(G270), .A3(new_n282), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT79), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT79), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n485), .A2(new_n488), .A3(G270), .A4(new_n282), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n484), .A2(new_n490), .ZN(new_n491));
  AND3_X1   g0291(.A1(new_n255), .A2(new_n256), .A3(new_n440), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(G116), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n262), .A2(new_n218), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n253), .A2(new_n229), .B1(G20), .B2(new_n218), .ZN(new_n495));
  NAND2_X1  g0295(.A1(G33), .A2(G283), .ZN(new_n496));
  INV_X1    g0296(.A(G97), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n496), .B(new_n207), .C1(G33), .C2(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(KEYINPUT20), .B1(new_n495), .B2(new_n498), .ZN(new_n499));
  AND3_X1   g0299(.A1(new_n495), .A2(KEYINPUT20), .A3(new_n498), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n493), .B(new_n494), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n491), .A2(new_n501), .A3(G169), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT21), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT80), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI211_X1 g0306(.A(new_n503), .B(new_n318), .C1(new_n484), .C2(new_n490), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n491), .A2(new_n328), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n501), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n502), .A2(KEYINPUT80), .A3(new_n503), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n491), .A2(G200), .ZN(new_n511));
  INV_X1    g0311(.A(new_n501), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n511), .B(new_n512), .C1(new_n293), .C2(new_n491), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n506), .A2(new_n509), .A3(new_n510), .A4(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT81), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n318), .B1(new_n484), .B2(new_n490), .ZN(new_n516));
  AOI211_X1 g0316(.A(new_n505), .B(KEYINPUT21), .C1(new_n516), .C2(new_n501), .ZN(new_n517));
  AOI21_X1  g0317(.A(KEYINPUT80), .B1(new_n502), .B2(new_n503), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT81), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n519), .A2(new_n520), .A3(new_n509), .A4(new_n513), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n473), .B1(new_n515), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n485), .A2(G264), .A3(new_n282), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(KEYINPUT83), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT83), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n485), .A2(new_n525), .A3(G264), .A4(new_n282), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n479), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  OAI211_X1 g0327(.A(G257), .B(G1698), .C1(new_n350), .C2(new_n351), .ZN(new_n528));
  OAI211_X1 g0328(.A(G250), .B(new_n276), .C1(new_n350), .C2(new_n351), .ZN(new_n529));
  NAND2_X1  g0329(.A1(G33), .A2(G294), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT82), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n531), .A2(new_n532), .A3(new_n283), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n531), .A2(new_n283), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(KEYINPUT82), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n527), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G169), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n524), .A2(new_n526), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n538), .A2(G179), .A3(new_n478), .A4(new_n534), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT24), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n207), .B(G87), .C1(new_n350), .C2(new_n351), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(KEYINPUT22), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT22), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n273), .A2(new_n544), .A3(new_n207), .A4(G87), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n454), .A2(G20), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n207), .A2(G107), .ZN(new_n549));
  XNOR2_X1  g0349(.A(new_n549), .B(KEYINPUT23), .ZN(new_n550));
  AND4_X1   g0350(.A1(new_n541), .A2(new_n546), .A3(new_n548), .A4(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n547), .B1(new_n543), .B2(new_n545), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n541), .B1(new_n552), .B2(new_n550), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n254), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n492), .A2(G107), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n256), .A2(G107), .ZN(new_n556));
  XNOR2_X1  g0356(.A(new_n556), .B(KEYINPUT25), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n554), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n540), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n538), .A2(new_n478), .A3(new_n534), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n471), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n527), .A2(new_n293), .A3(new_n533), .A4(new_n535), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n563), .A2(new_n555), .A3(new_n554), .A4(new_n557), .ZN(new_n564));
  AND2_X1   g0364(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n485), .A2(G257), .A3(new_n282), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n478), .ZN(new_n567));
  OAI211_X1 g0367(.A(G244), .B(new_n276), .C1(new_n350), .C2(new_n351), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT4), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n273), .A2(KEYINPUT4), .A3(G244), .A4(new_n276), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n273), .A2(G250), .A3(G1698), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n570), .A2(new_n571), .A3(new_n496), .A4(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n567), .B1(new_n573), .B2(new_n283), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(G179), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n318), .B2(new_n574), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n262), .A2(new_n497), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n492), .A2(G97), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n333), .B1(new_n370), .B2(new_n357), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT6), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n497), .A2(new_n333), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n580), .B1(new_n581), .B2(new_n431), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n333), .A2(KEYINPUT6), .A3(G97), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n207), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n267), .A2(new_n275), .ZN(new_n585));
  NOR3_X1   g0385(.A1(new_n579), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n577), .B(new_n578), .C1(new_n586), .C2(new_n255), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n576), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n573), .A2(new_n283), .ZN(new_n589));
  INV_X1    g0389(.A(new_n567), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(KEYINPUT75), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT75), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n574), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n592), .A2(new_n594), .A3(G200), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT76), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT73), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n587), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n371), .A2(G107), .ZN(new_n600));
  INV_X1    g0400(.A(new_n584), .ZN(new_n601));
  INV_X1    g0401(.A(new_n585), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n254), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n604), .A2(KEYINPUT73), .A3(new_n577), .A4(new_n578), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n599), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n574), .A2(G190), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n592), .A2(new_n594), .A3(KEYINPUT76), .A4(G200), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n597), .A2(new_n606), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n565), .A2(new_n588), .A3(new_n609), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n428), .A2(new_n522), .A3(new_n610), .ZN(G372));
  NAND3_X1  g0411(.A1(new_n599), .A2(new_n605), .A3(new_n576), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT85), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n456), .A2(KEYINPUT84), .A3(new_n283), .ZN(new_n614));
  AOI21_X1  g0414(.A(KEYINPUT84), .B1(new_n456), .B2(new_n283), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n463), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n470), .B1(G200), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n464), .A2(new_n442), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n618), .B1(new_n318), .B2(new_n616), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n613), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n437), .B(new_n439), .C1(new_n389), .C2(new_n441), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n621), .B1(G190), .B2(new_n465), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT84), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n457), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n456), .A2(KEYINPUT84), .A3(new_n283), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n462), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n622), .B1(new_n626), .B2(new_n471), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n447), .B1(new_n328), .B2(new_n465), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n628), .B1(new_n626), .B2(G169), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n627), .A2(new_n629), .A3(KEYINPUT85), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n612), .B1(new_n620), .B2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT26), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(KEYINPUT26), .B1(new_n473), .B2(new_n588), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n629), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n559), .A2(new_n509), .A3(new_n506), .A4(new_n510), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n637), .A2(new_n588), .A3(new_n609), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n627), .A2(new_n629), .A3(KEYINPUT85), .ZN(new_n639));
  AOI21_X1  g0439(.A(KEYINPUT85), .B1(new_n627), .B2(new_n629), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n564), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n633), .B(new_n636), .C1(new_n638), .C2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n428), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n330), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n323), .A2(new_n324), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n645), .B1(new_n316), .B2(new_n348), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n646), .A2(new_n410), .A3(new_n422), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n418), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n644), .B1(new_n648), .B2(new_n295), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n643), .A2(new_n649), .ZN(G369));
  INV_X1    g0450(.A(G330), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n515), .A2(new_n521), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n209), .A2(G20), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(new_n206), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n655), .A2(G213), .A3(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(G343), .ZN(new_n659));
  XNOR2_X1  g0459(.A(new_n659), .B(KEYINPUT86), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n652), .B1(new_n512), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n519), .A2(new_n509), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n660), .A2(new_n512), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n651), .B1(new_n661), .B2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n660), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n558), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n565), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n668), .B1(new_n559), .B2(new_n660), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n666), .B1(new_n519), .B2(new_n509), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n565), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(new_n559), .B2(new_n666), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n671), .A2(new_n674), .ZN(G399));
  NOR2_X1   g0475(.A1(new_n213), .A2(G41), .ZN(new_n676));
  AOI21_X1  g0476(.A(KEYINPUT87), .B1(new_n676), .B2(new_n234), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n431), .A2(new_n389), .A3(new_n218), .ZN(new_n678));
  NOR3_X1   g0478(.A1(new_n676), .A2(new_n206), .A3(new_n678), .ZN(new_n679));
  MUX2_X1   g0479(.A(new_n677), .B(KEYINPUT87), .S(new_n679), .Z(new_n680));
  XNOR2_X1  g0480(.A(new_n680), .B(KEYINPUT88), .ZN(new_n681));
  XOR2_X1   g0481(.A(new_n681), .B(KEYINPUT28), .Z(new_n682));
  INV_X1    g0482(.A(KEYINPUT29), .ZN(new_n683));
  OR3_X1    g0483(.A1(new_n473), .A2(new_n588), .A3(KEYINPUT26), .ZN(new_n684));
  OAI211_X1 g0484(.A(new_n629), .B(new_n684), .C1(new_n631), .C2(new_n632), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n641), .A2(new_n638), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n683), .B1(new_n687), .B2(new_n660), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n609), .A2(new_n588), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n620), .A2(new_n630), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n689), .A2(new_n564), .A3(new_n690), .A4(new_n637), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n635), .B1(new_n631), .B2(new_n632), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n666), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n683), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n522), .A2(new_n610), .A3(new_n660), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n560), .A2(new_n591), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(KEYINPUT89), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n698), .A2(new_n491), .A3(new_n616), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n328), .B1(new_n697), .B2(KEYINPUT89), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n574), .A2(G179), .A3(new_n484), .A4(new_n490), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n465), .A2(new_n534), .A3(new_n538), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT30), .ZN(new_n704));
  OR3_X1    g0504(.A1(new_n702), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n704), .B1(new_n702), .B2(new_n703), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n666), .B1(new_n701), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(KEYINPUT31), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT31), .ZN(new_n710));
  OAI211_X1 g0510(.A(new_n710), .B(new_n666), .C1(new_n701), .C2(new_n707), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n696), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(G330), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR3_X1   g0515(.A1(new_n688), .A2(new_n695), .A3(new_n715), .ZN(new_n716));
  XOR2_X1   g0516(.A(new_n716), .B(KEYINPUT90), .Z(new_n717));
  OAI21_X1  g0517(.A(new_n682), .B1(new_n717), .B2(G1), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT91), .ZN(G364));
  INV_X1    g0519(.A(new_n676), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n653), .A2(G45), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n720), .A2(G1), .A3(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n665), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n661), .A2(new_n664), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n724), .B1(G330), .B2(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n229), .B1(G20), .B2(new_n318), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n207), .A2(new_n328), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(new_n471), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(new_n293), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n293), .A2(G179), .A3(G200), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(new_n207), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AOI22_X1  g0536(.A1(new_n733), .A2(G326), .B1(G294), .B2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(G311), .ZN(new_n738));
  NOR2_X1   g0538(.A1(G190), .A2(G200), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n729), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n737), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  XOR2_X1   g0541(.A(new_n741), .B(KEYINPUT98), .Z(new_n742));
  NOR3_X1   g0542(.A1(new_n730), .A2(new_n293), .A3(G200), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G322), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n207), .A2(G179), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n745), .A2(new_n293), .A3(G200), .ZN(new_n746));
  INV_X1    g0546(.A(G283), .ZN(new_n747));
  INV_X1    g0547(.A(G303), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n745), .A2(G190), .A3(G200), .ZN(new_n749));
  OAI221_X1 g0549(.A(new_n352), .B1(new_n746), .B2(new_n747), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  AND2_X1   g0550(.A1(new_n745), .A2(new_n739), .ZN(new_n751));
  OR2_X1    g0551(.A1(new_n751), .A2(KEYINPUT95), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(KEYINPUT95), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AND2_X1   g0555(.A1(new_n755), .A2(G329), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n731), .A2(KEYINPUT97), .A3(new_n293), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(KEYINPUT97), .B1(new_n731), .B2(new_n293), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  XNOR2_X1  g0561(.A(KEYINPUT33), .B(G317), .ZN(new_n762));
  AOI211_X1 g0562(.A(new_n750), .B(new_n756), .C1(new_n761), .C2(new_n762), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n742), .A2(new_n744), .A3(new_n763), .ZN(new_n764));
  XOR2_X1   g0564(.A(new_n740), .B(KEYINPUT93), .Z(new_n765));
  AOI22_X1  g0565(.A1(new_n765), .A2(G77), .B1(G58), .B2(new_n743), .ZN(new_n766));
  INV_X1    g0566(.A(new_n733), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n766), .B1(new_n202), .B2(new_n767), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n768), .B(KEYINPUT94), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n760), .A2(new_n223), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n273), .B1(new_n749), .B2(new_n389), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n735), .A2(new_n497), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n746), .A2(new_n333), .ZN(new_n773));
  NOR4_X1   g0573(.A1(new_n770), .A2(new_n771), .A3(new_n772), .A4(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n754), .A2(new_n360), .ZN(new_n775));
  XNOR2_X1  g0575(.A(KEYINPUT96), .B(KEYINPUT32), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n769), .A2(new_n774), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n728), .B1(new_n764), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G13), .A2(G33), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(G20), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n727), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n214), .A2(new_n352), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT92), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n248), .A2(G45), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n785), .B(new_n786), .C1(G45), .C2(new_n233), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n214), .A2(G355), .A3(new_n273), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n787), .B(new_n788), .C1(G116), .C2(new_n214), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n779), .B1(new_n783), .B2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n782), .ZN(new_n791));
  OAI211_X1 g0591(.A(new_n790), .B(new_n723), .C1(new_n725), .C2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n726), .A2(new_n792), .ZN(G396));
  AOI22_X1  g0593(.A1(G159), .A2(new_n765), .B1(new_n733), .B2(G137), .ZN(new_n794));
  INV_X1    g0594(.A(G143), .ZN(new_n795));
  INV_X1    g0595(.A(new_n743), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n794), .B1(new_n795), .B2(new_n796), .C1(new_n265), .C2(new_n760), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n797), .B(KEYINPUT34), .Z(new_n798));
  OAI21_X1  g0598(.A(new_n273), .B1(new_n749), .B2(new_n202), .ZN(new_n799));
  INV_X1    g0599(.A(new_n746), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n799), .B1(G68), .B2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(G58), .ZN(new_n802));
  INV_X1    g0602(.A(G132), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n801), .B1(new_n802), .B2(new_n735), .C1(new_n754), .C2(new_n803), .ZN(new_n804));
  XOR2_X1   g0604(.A(new_n804), .B(KEYINPUT100), .Z(new_n805));
  NOR2_X1   g0605(.A1(new_n746), .A2(new_n389), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n767), .A2(new_n748), .B1(new_n749), .B2(new_n333), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n807), .B1(new_n761), .B2(G283), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n772), .B1(new_n755), .B2(G311), .ZN(new_n809));
  INV_X1    g0609(.A(G294), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n352), .B1(new_n796), .B2(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n811), .B1(new_n765), .B2(G116), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n808), .A2(new_n809), .A3(new_n812), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n798), .A2(new_n805), .B1(new_n806), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n348), .A2(new_n660), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT101), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n348), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g0617(.A1(new_n339), .A2(new_n346), .A3(KEYINPUT101), .A4(new_n347), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n817), .A2(new_n818), .B1(new_n425), .B2(new_n424), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n666), .A2(new_n346), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n815), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n727), .A2(new_n814), .B1(new_n821), .B2(new_n780), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n727), .A2(new_n780), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT99), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(new_n275), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n722), .B1(new_n822), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n642), .A2(new_n660), .A3(new_n819), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n821), .B(KEYINPUT102), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n827), .B1(new_n828), .B2(new_n693), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(new_n714), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n826), .B1(new_n830), .B2(new_n722), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT103), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(G384));
  NAND2_X1  g0633(.A1(new_n407), .A2(new_n658), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT105), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n407), .A2(KEYINPUT105), .A3(new_n658), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n423), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n421), .A2(new_n414), .ZN(new_n840));
  OAI21_X1  g0640(.A(KEYINPUT37), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n421), .A2(new_n414), .A3(new_n834), .ZN(new_n842));
  OR2_X1    g0642(.A1(new_n842), .A2(KEYINPUT37), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n839), .A2(new_n844), .A3(KEYINPUT38), .ZN(new_n845));
  INV_X1    g0645(.A(new_n834), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n842), .A2(KEYINPUT37), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n423), .A2(new_n846), .B1(new_n843), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n845), .B1(KEYINPUT38), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n316), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT104), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n645), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n660), .A2(new_n314), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n854), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n325), .A2(new_n852), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n821), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT106), .ZN(new_n859));
  AND3_X1   g0659(.A1(new_n696), .A2(new_n859), .A3(new_n712), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n859), .B1(new_n696), .B2(new_n712), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n858), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(KEYINPUT40), .B1(new_n850), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(KEYINPUT38), .B1(new_n839), .B2(new_n844), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n845), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT40), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n713), .A2(KEYINPUT106), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n696), .A2(new_n859), .A3(new_n712), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n866), .A2(new_n867), .A3(new_n870), .A4(new_n858), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n863), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n870), .A2(new_n428), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n872), .B(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(G330), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n817), .A2(new_n660), .A3(new_n818), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n827), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n855), .A2(new_n857), .ZN(new_n878));
  AND3_X1   g0678(.A1(new_n839), .A2(new_n844), .A3(KEYINPUT38), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n877), .B(new_n878), .C1(new_n879), .C2(new_n864), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n645), .A2(new_n666), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(KEYINPUT39), .B1(new_n879), .B2(new_n864), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT39), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n845), .B(new_n885), .C1(KEYINPUT38), .C2(new_n848), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n883), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n418), .A2(new_n658), .ZN(new_n888));
  NOR3_X1   g0688(.A1(new_n881), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n875), .B(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n428), .B1(new_n695), .B2(new_n688), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n649), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n890), .B(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n206), .B2(new_n653), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n582), .A2(new_n583), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n218), .B1(new_n895), .B2(KEYINPUT35), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n896), .B(new_n231), .C1(KEYINPUT35), .C2(new_n895), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n897), .B(KEYINPUT36), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n363), .A2(G77), .ZN(new_n899));
  OAI22_X1  g0699(.A1(new_n233), .A2(new_n899), .B1(G50), .B2(new_n223), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n900), .A2(G1), .A3(new_n209), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n894), .A2(new_n898), .A3(new_n901), .ZN(G367));
  INV_X1    g0702(.A(new_n690), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n666), .A2(new_n621), .ZN(new_n904));
  MUX2_X1   g0704(.A(new_n629), .B(new_n903), .S(new_n904), .Z(new_n905));
  XOR2_X1   g0705(.A(new_n905), .B(KEYINPUT107), .Z(new_n906));
  INV_X1    g0706(.A(KEYINPUT43), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n689), .B1(new_n606), .B2(new_n660), .ZN(new_n909));
  OR2_X1    g0709(.A1(new_n612), .A2(new_n660), .ZN(new_n910));
  AND3_X1   g0710(.A1(new_n909), .A2(KEYINPUT108), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT108), .B1(new_n909), .B2(new_n910), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n913), .A2(new_n673), .ZN(new_n914));
  XOR2_X1   g0714(.A(new_n914), .B(KEYINPUT42), .Z(new_n915));
  OR2_X1    g0715(.A1(new_n913), .A2(new_n559), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n666), .B1(new_n916), .B2(new_n588), .ZN(new_n917));
  OAI221_X1 g0717(.A(new_n908), .B1(new_n907), .B2(new_n905), .C1(new_n915), .C2(new_n917), .ZN(new_n918));
  OR3_X1    g0718(.A1(new_n915), .A2(new_n917), .A3(new_n908), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n913), .A2(new_n670), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n920), .B(new_n921), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n676), .B(KEYINPUT41), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n913), .A2(new_n674), .B1(KEYINPUT109), .B2(KEYINPUT44), .ZN(new_n925));
  OR2_X1    g0725(.A1(KEYINPUT109), .A2(KEYINPUT44), .ZN(new_n926));
  XOR2_X1   g0726(.A(new_n925), .B(new_n926), .Z(new_n927));
  NOR2_X1   g0727(.A1(new_n913), .A2(new_n674), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n928), .B(KEYINPUT45), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n671), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n927), .A2(new_n670), .A3(new_n929), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n673), .B1(new_n669), .B2(new_n672), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n665), .B(new_n933), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n931), .A2(new_n717), .A3(new_n932), .A4(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n924), .B1(new_n935), .B2(new_n717), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n721), .A2(G1), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n922), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n735), .A2(new_n223), .ZN(new_n939));
  INV_X1    g0739(.A(G137), .ZN(new_n940));
  OAI221_X1 g0740(.A(new_n273), .B1(new_n265), .B2(new_n796), .C1(new_n754), .C2(new_n940), .ZN(new_n941));
  AOI211_X1 g0741(.A(new_n939), .B(new_n941), .C1(G50), .C2(new_n765), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n767), .A2(new_n795), .B1(new_n749), .B2(new_n802), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(new_n761), .B2(G159), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n942), .B(new_n944), .C1(new_n275), .C2(new_n746), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT110), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT46), .ZN(new_n947));
  NOR3_X1   g0747(.A1(new_n749), .A2(new_n947), .A3(new_n218), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n947), .B1(new_n749), .B2(new_n218), .ZN(new_n949));
  INV_X1    g0749(.A(new_n765), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n949), .B1(new_n950), .B2(new_n747), .ZN(new_n951));
  AOI211_X1 g0751(.A(new_n948), .B(new_n951), .C1(G317), .C2(new_n755), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n746), .A2(new_n497), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(G107), .B2(new_n736), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n352), .B(new_n954), .C1(new_n767), .C2(new_n738), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(G294), .B2(new_n761), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n952), .B(new_n956), .C1(new_n748), .C2(new_n796), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n946), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT47), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n722), .B1(new_n959), .B2(new_n727), .ZN(new_n960));
  INV_X1    g0760(.A(new_n785), .ZN(new_n961));
  OAI221_X1 g0761(.A(new_n783), .B1(new_n214), .B2(new_n343), .C1(new_n961), .C2(new_n243), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n905), .A2(new_n782), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n960), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n938), .A2(new_n964), .ZN(G387));
  AND2_X1   g0765(.A1(new_n755), .A2(G326), .ZN(new_n966));
  AOI22_X1  g0766(.A1(G303), .A2(new_n765), .B1(new_n733), .B2(G322), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n738), .B2(new_n760), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n968), .B1(G317), .B2(new_n743), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n969), .B(KEYINPUT48), .Z(new_n970));
  OAI221_X1 g0770(.A(new_n970), .B1(new_n747), .B2(new_n735), .C1(new_n810), .C2(new_n749), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT49), .ZN(new_n972));
  AOI211_X1 g0772(.A(new_n273), .B(new_n966), .C1(new_n971), .C2(new_n972), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n973), .B1(new_n972), .B2(new_n971), .C1(new_n218), .C2(new_n746), .ZN(new_n974));
  AND3_X1   g0774(.A1(new_n733), .A2(KEYINPUT112), .A3(G159), .ZN(new_n975));
  AOI21_X1  g0775(.A(KEYINPUT112), .B1(new_n733), .B2(G159), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n754), .A2(new_n265), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n273), .B1(new_n740), .B2(new_n223), .ZN(new_n978));
  NOR4_X1   g0778(.A1(new_n975), .A2(new_n976), .A3(new_n977), .A4(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n202), .B2(new_n796), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n749), .A2(new_n275), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n760), .A2(new_n268), .B1(new_n343), .B2(new_n735), .ZN(new_n982));
  OR4_X1    g0782(.A1(new_n953), .A2(new_n980), .A3(new_n981), .A4(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n728), .B1(new_n974), .B2(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n669), .A2(new_n791), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n214), .A2(new_n273), .A3(new_n678), .ZN(new_n986));
  OR3_X1    g0786(.A1(new_n268), .A2(KEYINPUT50), .A3(G50), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n678), .B1(G68), .B2(G77), .ZN(new_n988));
  OAI21_X1  g0788(.A(KEYINPUT50), .B1(new_n268), .B2(G50), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n987), .A2(new_n988), .A3(new_n989), .A4(new_n458), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n785), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT111), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n240), .A2(new_n458), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n986), .B1(G107), .B2(new_n214), .C1(new_n992), .C2(new_n993), .ZN(new_n994));
  AND2_X1   g0794(.A1(new_n994), .A2(new_n783), .ZN(new_n995));
  NOR3_X1   g0795(.A1(new_n984), .A2(new_n985), .A3(new_n995), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n996), .A2(new_n723), .B1(new_n937), .B2(new_n934), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n717), .A2(new_n934), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n676), .B1(new_n717), .B2(new_n934), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n997), .B1(new_n999), .B2(new_n1000), .ZN(G393));
  NAND2_X1  g0801(.A1(new_n931), .A2(new_n932), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n720), .B1(new_n1002), .B2(new_n998), .ZN(new_n1003));
  AND2_X1   g0803(.A1(new_n1003), .A2(new_n935), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n913), .A2(new_n782), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n783), .B1(new_n497), .B2(new_n214), .C1(new_n961), .C2(new_n251), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n733), .A2(G317), .B1(G311), .B2(new_n743), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n761), .A2(G303), .B1(new_n1007), .B2(KEYINPUT52), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n735), .A2(new_n218), .B1(new_n749), .B2(new_n747), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1009), .A2(new_n773), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n352), .B1(new_n740), .B2(new_n810), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(new_n755), .B2(G322), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1008), .A2(new_n1010), .A3(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1007), .A2(KEYINPUT52), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n761), .A2(G50), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n735), .A2(new_n275), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n755), .A2(G143), .B1(new_n340), .B2(new_n765), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n749), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n352), .B(new_n806), .C1(G68), .C2(new_n1019), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1015), .A2(new_n1017), .A3(new_n1018), .A4(new_n1020), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n733), .A2(G150), .B1(G159), .B2(new_n743), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT51), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n1013), .A2(new_n1014), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n722), .B1(new_n1024), .B2(new_n727), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1005), .A2(new_n1006), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n937), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1026), .B1(new_n1002), .B2(new_n1027), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n1004), .A2(new_n1028), .ZN(G390));
  OAI211_X1 g0829(.A(new_n660), .B(new_n819), .C1(new_n685), .C2(new_n686), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n876), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n878), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1032), .A2(new_n849), .A3(new_n883), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n715), .A2(new_n858), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n884), .A2(new_n886), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n882), .B1(new_n877), .B2(new_n878), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1033), .B(new_n1034), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(KEYINPUT113), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1033), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1039));
  OAI211_X1 g0839(.A(G330), .B(new_n858), .C1(new_n860), .C2(new_n861), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n876), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(new_n693), .B2(new_n819), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n878), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n883), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1046), .A2(new_n884), .A3(new_n886), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT113), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1047), .A2(new_n1048), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1038), .A2(new_n1042), .A3(new_n1049), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n1050), .A2(new_n1027), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n754), .A2(new_n810), .B1(new_n389), .B2(new_n749), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n352), .B1(new_n218), .B2(new_n796), .C1(new_n950), .C2(new_n497), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n767), .A2(new_n747), .B1(new_n746), .B2(new_n223), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1017), .B1(new_n760), .B2(new_n333), .ZN(new_n1055));
  OR4_X1    g0855(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .A4(new_n1055), .ZN(new_n1056));
  XOR2_X1   g0856(.A(KEYINPUT54), .B(G143), .Z(new_n1057));
  AOI22_X1  g0857(.A1(new_n755), .A2(G125), .B1(new_n765), .B2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n746), .A2(new_n202), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n273), .B1(new_n735), .B2(new_n360), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n1059), .B(new_n1060), .C1(new_n733), .C2(G128), .ZN(new_n1061));
  AND2_X1   g0861(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1062), .B1(new_n803), .B2(new_n796), .C1(new_n940), .C2(new_n760), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n749), .A2(new_n265), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT115), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT53), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1056), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n1067), .A2(new_n727), .B1(new_n268), .B2(new_n824), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n723), .B(new_n1068), .C1(new_n1035), .C2(new_n781), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n651), .B(new_n821), .C1(new_n696), .C2(new_n712), .ZN(new_n1070));
  OAI21_X1  g0870(.A(KEYINPUT114), .B1(new_n1070), .B2(new_n878), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n821), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n713), .A2(G330), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT114), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1073), .A2(new_n1074), .A3(new_n1045), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1071), .A2(new_n1040), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n877), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n828), .B(G330), .C1(new_n860), .C2(new_n861), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n1045), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1031), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1079), .A2(new_n1080), .A3(new_n1034), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1077), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n870), .A2(new_n428), .A3(G330), .ZN(new_n1083));
  AND3_X1   g0883(.A1(new_n891), .A2(new_n1083), .A3(new_n649), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  AND2_X1   g0885(.A1(new_n1050), .A2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n676), .B1(new_n1050), .B2(new_n1085), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1051), .B(new_n1069), .C1(new_n1086), .C2(new_n1087), .ZN(G378));
  OAI21_X1  g0888(.A(new_n1084), .B1(new_n1050), .B2(new_n1085), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(KEYINPUT118), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n295), .A2(new_n330), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n326), .A2(new_n658), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1091), .B(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT55), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT56), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1035), .A2(new_n882), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n888), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1096), .A2(new_n880), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n651), .B1(new_n863), .B2(new_n871), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1095), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT56), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1094), .B(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n872), .A2(G330), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n889), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1104), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1102), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT118), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1110), .B(new_n1084), .C1(new_n1050), .C2(new_n1085), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1090), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT57), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1090), .A2(new_n1109), .A3(KEYINPUT57), .A4(new_n1111), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1114), .A2(new_n676), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1109), .A2(new_n937), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1104), .A2(new_n780), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n733), .A2(G125), .B1(G150), .B2(new_n736), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n743), .A2(G128), .B1(new_n1019), .B2(new_n1057), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n1121), .B1(new_n803), .B2(new_n760), .C1(new_n940), .C2(new_n740), .ZN(new_n1122));
  XOR2_X1   g0922(.A(new_n1122), .B(KEYINPUT59), .Z(new_n1123));
  AOI21_X1  g0923(.A(G41), .B1(new_n755), .B2(G124), .ZN(new_n1124));
  AOI21_X1  g0924(.A(G33), .B1(new_n800), .B2(G159), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1123), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n202), .B1(new_n350), .B2(G41), .ZN(new_n1127));
  AOI21_X1  g0927(.A(G41), .B1(new_n743), .B2(G107), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n740), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n273), .B1(new_n1129), .B2(new_n342), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1128), .B(new_n1130), .C1(new_n754), .C2(new_n747), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n746), .A2(new_n802), .ZN(new_n1132));
  NOR4_X1   g0932(.A1(new_n1131), .A2(new_n939), .A3(new_n981), .A4(new_n1132), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n1133), .B1(new_n497), .B2(new_n760), .C1(new_n218), .C2(new_n767), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT58), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1126), .A2(new_n1127), .A3(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n727), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n722), .B1(new_n202), .B2(new_n823), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT116), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1118), .A2(new_n1137), .A3(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1117), .A2(KEYINPUT117), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT117), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1027), .B1(new_n1102), .B2(new_n1108), .ZN(new_n1143));
  AND3_X1   g0943(.A1(new_n1118), .A2(new_n1137), .A3(new_n1139), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1142), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1141), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1116), .A2(new_n1146), .ZN(G375));
  INV_X1    g0947(.A(KEYINPUT119), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n1078), .A2(new_n1045), .B1(new_n715), .B2(new_n858), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n1080), .A2(new_n1149), .B1(new_n1076), .B2(new_n877), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1148), .B1(new_n1150), .B2(new_n1027), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n343), .A2(new_n735), .B1(new_n497), .B2(new_n749), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(new_n761), .B2(G116), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n733), .A2(G294), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n765), .A2(G107), .B1(G77), .B2(new_n800), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n352), .B1(new_n796), .B2(new_n747), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(new_n755), .B2(G303), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1153), .A2(new_n1154), .A3(new_n1155), .A4(new_n1157), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1132), .A2(new_n352), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n1159), .B(KEYINPUT122), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(new_n761), .B2(new_n1057), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n735), .A2(new_n202), .B1(new_n740), .B2(new_n265), .ZN(new_n1162));
  XOR2_X1   g0962(.A(new_n1162), .B(KEYINPUT121), .Z(new_n1163));
  NAND2_X1  g0963(.A1(new_n733), .A2(G132), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT120), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n749), .A2(new_n360), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(new_n755), .B2(G128), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1161), .A2(new_n1163), .A3(new_n1165), .A4(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n796), .A2(new_n940), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1158), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n1170), .A2(new_n727), .B1(new_n223), .B2(new_n824), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n723), .B(new_n1171), .C1(new_n878), .C2(new_n781), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1082), .A2(KEYINPUT119), .A3(new_n937), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1151), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(KEYINPUT123), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT123), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1151), .A2(new_n1173), .A3(new_n1176), .A4(new_n1172), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1179), .A2(new_n924), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(new_n1085), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1178), .A2(new_n1181), .ZN(G381));
  INV_X1    g0982(.A(KEYINPUT125), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(G375), .B(new_n1183), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1004), .A2(new_n1028), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1185), .A2(new_n964), .A3(new_n938), .ZN(new_n1186));
  NOR4_X1   g0986(.A1(new_n1186), .A2(G396), .A3(G393), .A4(G381), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(G378), .B(KEYINPUT124), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1184), .A2(new_n832), .A3(new_n1187), .A4(new_n1188), .ZN(G407));
  INV_X1    g0989(.A(G343), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1184), .A2(new_n1190), .A3(new_n1188), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(G407), .A2(G213), .A3(new_n1191), .ZN(G409));
  INV_X1    g0992(.A(KEYINPUT127), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1116), .A2(G378), .A3(new_n1146), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1117), .B(new_n1140), .C1(new_n1112), .C2(new_n924), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1188), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1190), .A2(G213), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1190), .A2(KEYINPUT126), .A3(G213), .ZN(new_n1199));
  OR2_X1    g0999(.A1(new_n1179), .A2(KEYINPUT60), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1179), .A2(KEYINPUT60), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1200), .A2(new_n676), .A3(new_n1085), .A4(new_n1201), .ZN(new_n1202));
  AND3_X1   g1002(.A1(new_n1178), .A2(new_n1202), .A3(new_n832), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n832), .B1(new_n1178), .B2(new_n1202), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1199), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1190), .A2(G213), .A3(G2897), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1206), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1208), .B(new_n1199), .C1(new_n1203), .C2(new_n1204), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n1197), .A2(new_n1198), .B1(new_n1207), .B2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1193), .B1(new_n1210), .B2(KEYINPUT61), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT61), .ZN(new_n1212));
  AND2_X1   g1012(.A1(new_n1207), .A2(new_n1209), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n1194), .A2(new_n1196), .B1(G213), .B2(new_n1190), .ZN(new_n1214));
  OAI211_X1 g1014(.A(KEYINPUT127), .B(new_n1212), .C1(new_n1213), .C2(new_n1214), .ZN(new_n1215));
  OR2_X1    g1015(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1214), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(KEYINPUT62), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT62), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1214), .A2(new_n1219), .A3(new_n1216), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1211), .A2(new_n1215), .A3(new_n1218), .A4(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(G387), .A2(G390), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(new_n1186), .ZN(new_n1223));
  XOR2_X1   g1023(.A(G393), .B(G396), .Z(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1224), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1222), .A2(new_n1186), .A3(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1225), .A2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1221), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT63), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1217), .A2(new_n1230), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1231), .A2(new_n1228), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1217), .B1(new_n1210), .B2(new_n1230), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1232), .A2(new_n1212), .A3(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1229), .A2(new_n1234), .ZN(G405));
  NAND2_X1  g1035(.A1(G375), .A2(new_n1188), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1228), .A2(new_n1194), .A3(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1216), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1236), .A2(new_n1194), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1225), .A2(new_n1227), .A3(new_n1239), .ZN(new_n1240));
  AND3_X1   g1040(.A1(new_n1237), .A2(new_n1238), .A3(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1238), .B1(new_n1237), .B2(new_n1240), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1241), .A2(new_n1242), .ZN(G402));
endmodule


