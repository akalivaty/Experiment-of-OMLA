//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 0 1 1 0 0 1 0 0 1 0 0 1 0 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 1 0 1 0 1 0 1 0 1 1 1 1 0 1 1 1 1 1 1 1 1 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:27 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n451, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n555, new_n557, new_n558,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n621, new_n624, new_n625,
    new_n626, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1227, new_n1228;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT65), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT66), .ZN(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT67), .ZN(G217));
  NAND4_X1  g027(.A1(new_n437), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n455), .A2(G567), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n458), .A2(KEYINPUT68), .ZN(new_n459));
  AOI21_X1  g034(.A(new_n459), .B1(new_n454), .B2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(KEYINPUT68), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G101), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(KEYINPUT3), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G137), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n469), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n468), .B1(new_n464), .B2(new_n476), .ZN(G160));
  INV_X1    g052(.A(KEYINPUT69), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n465), .A2(KEYINPUT69), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n479), .A2(new_n480), .A3(G2105), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n479), .A2(new_n480), .A3(new_n464), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n483), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  NAND3_X1  g065(.A1(new_n464), .A2(G102), .A3(G2104), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(new_n470), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n493), .B1(new_n465), .B2(G126), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n491), .B1(new_n494), .B2(new_n464), .ZN(new_n495));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(KEYINPUT70), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n497), .A2(new_n471), .A3(new_n473), .A4(new_n464), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n465), .A2(KEYINPUT4), .A3(new_n464), .A4(new_n497), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n495), .A2(new_n502), .ZN(G164));
  XNOR2_X1  g078(.A(KEYINPUT5), .B(G543), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n504), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OR2_X1    g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G50), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT5), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G543), .ZN(new_n516));
  AND2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  OAI211_X1 g093(.A(new_n514), .B(new_n516), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  OAI22_X1  g095(.A1(new_n511), .A2(new_n512), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n507), .A2(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  NAND2_X1  g098(.A1(new_n514), .A2(new_n516), .ZN(new_n524));
  OAI21_X1  g099(.A(G89), .B1(new_n517), .B2(new_n518), .ZN(new_n525));
  NAND2_X1  g100(.A1(G63), .A2(G651), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  OAI211_X1 g102(.A(G51), .B(G543), .C1(new_n517), .C2(new_n518), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT7), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n530), .B(new_n531), .ZN(new_n532));
  NOR3_X1   g107(.A1(new_n527), .A2(new_n529), .A3(new_n532), .ZN(G168));
  INV_X1    g108(.A(G52), .ZN(new_n534));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n511), .A2(new_n534), .B1(new_n519), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n504), .A2(G64), .ZN(new_n537));
  NAND2_X1  g112(.A1(G77), .A2(G543), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n506), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n536), .A2(new_n539), .ZN(G171));
  AOI22_X1  g115(.A1(new_n504), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n541));
  OAI21_X1  g116(.A(KEYINPUT71), .B1(new_n541), .B2(new_n506), .ZN(new_n542));
  OAI211_X1 g117(.A(G43), .B(G543), .C1(new_n517), .C2(new_n518), .ZN(new_n543));
  INV_X1    g118(.A(G81), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n519), .B2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G56), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n524), .B2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT71), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n549), .A2(new_n550), .A3(G651), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n542), .A2(new_n546), .A3(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  AND3_X1   g129(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G36), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n555), .A2(new_n558), .ZN(G188));
  INV_X1    g134(.A(KEYINPUT73), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT72), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g138(.A1(KEYINPUT72), .A2(KEYINPUT9), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n513), .B1(new_n508), .B2(new_n509), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n565), .B1(G53), .B2(new_n566), .ZN(new_n567));
  OAI211_X1 g142(.A(G53), .B(G543), .C1(new_n517), .C2(new_n518), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n568), .A2(new_n563), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n560), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(G78), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(G65), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n524), .B2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n519), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n573), .A2(G651), .B1(new_n574), .B2(G91), .ZN(new_n575));
  OAI211_X1 g150(.A(new_n566), .B(G53), .C1(new_n561), .C2(new_n562), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n568), .B1(new_n564), .B2(new_n563), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n576), .A2(KEYINPUT73), .A3(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n570), .A2(new_n575), .A3(new_n578), .ZN(G299));
  INV_X1    g154(.A(G171), .ZN(G301));
  NAND2_X1  g155(.A1(G168), .A2(KEYINPUT74), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n530), .B(KEYINPUT7), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n510), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n583));
  OAI211_X1 g158(.A(new_n528), .B(new_n582), .C1(new_n583), .C2(new_n524), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT74), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n581), .A2(new_n586), .ZN(G286));
  NAND2_X1  g162(.A1(new_n574), .A2(G87), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n566), .A2(G49), .ZN(new_n589));
  OAI21_X1  g164(.A(G651), .B1(new_n504), .B2(G74), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(G288));
  AOI22_X1  g166(.A1(new_n504), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n506), .ZN(new_n593));
  INV_X1    g168(.A(G48), .ZN(new_n594));
  INV_X1    g169(.A(G86), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n511), .A2(new_n594), .B1(new_n519), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G305));
  AOI22_X1  g173(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n599), .A2(new_n506), .ZN(new_n600));
  INV_X1    g175(.A(G47), .ZN(new_n601));
  INV_X1    g176(.A(G85), .ZN(new_n602));
  OAI22_X1  g177(.A1(new_n511), .A2(new_n601), .B1(new_n519), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G79), .A2(G543), .ZN(new_n606));
  INV_X1    g181(.A(G66), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n524), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G651), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n566), .A2(G54), .ZN(new_n610));
  INV_X1    g185(.A(G92), .ZN(new_n611));
  OAI21_X1  g186(.A(KEYINPUT10), .B1(new_n519), .B2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT10), .ZN(new_n613));
  NAND4_X1  g188(.A1(new_n510), .A2(new_n504), .A3(new_n613), .A4(G92), .ZN(new_n614));
  NAND4_X1  g189(.A1(new_n609), .A2(new_n610), .A3(new_n612), .A4(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(G868), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(new_n616), .B2(G171), .ZN(G284));
  OAI21_X1  g193(.A(new_n617), .B1(new_n616), .B2(G171), .ZN(G321));
  NAND2_X1  g194(.A1(G299), .A2(new_n616), .ZN(new_n620));
  INV_X1    g195(.A(G286), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(new_n616), .ZN(G280));
  XOR2_X1   g197(.A(G280), .B(KEYINPUT75), .Z(G297));
  INV_X1    g198(.A(new_n615), .ZN(new_n624));
  XNOR2_X1  g199(.A(KEYINPUT76), .B(G559), .ZN(new_n625));
  INV_X1    g200(.A(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n624), .B1(G860), .B2(new_n626), .ZN(G148));
  NAND2_X1  g202(.A1(new_n552), .A2(new_n616), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n615), .A2(new_n625), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n629), .B2(new_n616), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g206(.A1(new_n482), .A2(G123), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n485), .A2(G135), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n634));
  INV_X1    g209(.A(KEYINPUT78), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g211(.A(KEYINPUT77), .B1(new_n464), .B2(G111), .ZN(new_n637));
  OR3_X1    g212(.A1(new_n464), .A2(KEYINPUT77), .A3(G111), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n634), .A2(new_n635), .ZN(new_n639));
  NAND4_X1  g214(.A1(new_n636), .A2(new_n637), .A3(new_n638), .A4(new_n639), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n632), .A2(new_n633), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(G2096), .Z(new_n642));
  NAND3_X1  g217(.A1(new_n464), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT12), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT13), .ZN(new_n645));
  INV_X1    g220(.A(G2100), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n642), .A2(new_n647), .ZN(G156));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2430), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2435), .ZN(new_n650));
  XOR2_X1   g225(.A(G2427), .B(G2438), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(KEYINPUT14), .ZN(new_n653));
  XOR2_X1   g228(.A(G1341), .B(G1348), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2451), .B(G2454), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT16), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT79), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n657), .B(new_n660), .Z(new_n661));
  AND2_X1   g236(.A1(new_n661), .A2(G14), .ZN(G401));
  XNOR2_X1  g237(.A(G2084), .B(G2090), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT80), .Z(new_n664));
  XOR2_X1   g239(.A(G2067), .B(G2678), .Z(new_n665));
  NOR2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2072), .B(G2078), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT18), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n667), .B(KEYINPUT17), .Z(new_n670));
  AOI21_X1  g245(.A(new_n670), .B1(new_n664), .B2(new_n665), .ZN(new_n671));
  INV_X1    g246(.A(new_n665), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n672), .A2(new_n667), .ZN(new_n673));
  AOI211_X1 g248(.A(new_n666), .B(new_n671), .C1(new_n664), .C2(new_n673), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n669), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(G2096), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(new_n646), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(G227));
  XOR2_X1   g253(.A(G1956), .B(G2474), .Z(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  NOR2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1971), .B(G1976), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT19), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n679), .A2(new_n680), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT20), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n685), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n682), .A2(new_n684), .A3(new_n686), .ZN(new_n690));
  OAI211_X1 g265(.A(new_n689), .B(new_n690), .C1(new_n688), .C2(new_n687), .ZN(new_n691));
  XOR2_X1   g266(.A(G1981), .B(G1986), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(G1991), .B(G1996), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT81), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n695), .B(new_n697), .ZN(G229));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G22), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(G166), .B2(new_n699), .ZN(new_n701));
  INV_X1    g276(.A(G1971), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(G16), .A2(G23), .ZN(new_n704));
  INV_X1    g279(.A(G288), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n704), .B1(new_n705), .B2(G16), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT33), .B(G1976), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n699), .A2(G6), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(new_n597), .B2(new_n699), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT32), .B(G1981), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n703), .A2(new_n708), .A3(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT82), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT34), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT36), .ZN(new_n717));
  INV_X1    g292(.A(G29), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n718), .A2(G25), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n482), .A2(G119), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n485), .A2(G131), .ZN(new_n721));
  NOR2_X1   g296(.A1(G95), .A2(G2105), .ZN(new_n722));
  OAI21_X1  g297(.A(G2104), .B1(new_n464), .B2(G107), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n720), .B(new_n721), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n719), .B1(new_n724), .B2(G29), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT35), .B(G1991), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n725), .A2(new_n727), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n699), .A2(G24), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(new_n604), .B2(new_n699), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G1986), .ZN(new_n732));
  NOR3_X1   g307(.A1(new_n728), .A2(new_n729), .A3(new_n732), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n716), .A2(new_n717), .A3(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n717), .B1(new_n716), .B2(new_n733), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n485), .A2(G141), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n482), .A2(G129), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n464), .A2(G105), .A3(G2104), .ZN(new_n740));
  NAND3_X1  g315(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT26), .Z(new_n742));
  NAND4_X1  g317(.A1(new_n738), .A2(new_n739), .A3(new_n740), .A4(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(KEYINPUT91), .ZN(new_n744));
  INV_X1    g319(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n743), .A2(KEYINPUT91), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(G29), .ZN(new_n748));
  INV_X1    g323(.A(G32), .ZN(new_n749));
  AOI21_X1  g324(.A(KEYINPUT92), .B1(new_n718), .B2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(KEYINPUT92), .B2(new_n748), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT27), .B(G1996), .Z(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT24), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n718), .B1(new_n757), .B2(G34), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n758), .A2(KEYINPUT88), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n757), .A2(G34), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(KEYINPUT88), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n759), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n762), .A2(KEYINPUT89), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(KEYINPUT89), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n466), .A2(new_n467), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n765), .A2(G2105), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n476), .A2(new_n464), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n763), .B(new_n764), .C1(new_n768), .C2(new_n718), .ZN(new_n769));
  INV_X1    g344(.A(G2084), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT90), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n699), .A2(G19), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n553), .B2(new_n699), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G1341), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT85), .B(KEYINPUT28), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n718), .A2(G26), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n485), .A2(KEYINPUT84), .A3(G140), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n482), .A2(G128), .ZN(new_n781));
  OR2_X1    g356(.A1(G104), .A2(G2105), .ZN(new_n782));
  OAI211_X1 g357(.A(new_n782), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT84), .ZN(new_n784));
  INV_X1    g359(.A(G140), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n784), .B1(new_n484), .B2(new_n785), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n780), .A2(new_n781), .A3(new_n783), .A4(new_n786), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n779), .B1(new_n787), .B2(G29), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G2067), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n753), .A2(new_n755), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n756), .A2(new_n776), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n699), .A2(KEYINPUT23), .A3(G20), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT23), .ZN(new_n793));
  INV_X1    g368(.A(G20), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n793), .B1(new_n794), .B2(G16), .ZN(new_n795));
  INV_X1    g370(.A(G299), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n792), .B(new_n795), .C1(new_n796), .C2(new_n699), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G1956), .ZN(new_n798));
  NOR2_X1   g373(.A1(G4), .A2(G16), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(new_n624), .B2(G16), .ZN(new_n800));
  XNOR2_X1  g375(.A(KEYINPUT83), .B(G1348), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n769), .A2(new_n770), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n718), .A2(G27), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G164), .B2(new_n718), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT94), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G2078), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  NOR4_X1   g384(.A1(new_n791), .A2(new_n798), .A3(new_n804), .A4(new_n809), .ZN(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT31), .B(G11), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT30), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n812), .A2(G28), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(G28), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n813), .A2(new_n814), .A3(new_n718), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(G171), .A2(G16), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(G5), .B2(G16), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n819), .A2(G1961), .ZN(new_n820));
  INV_X1    g395(.A(G1966), .ZN(new_n821));
  NAND2_X1  g396(.A1(G168), .A2(G16), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(G16), .B2(G21), .ZN(new_n823));
  AOI211_X1 g398(.A(new_n816), .B(new_n820), .C1(new_n821), .C2(new_n823), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n821), .B2(new_n823), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n819), .A2(G1961), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT93), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(new_n718), .B2(new_n641), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT86), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(G29), .B2(G33), .ZN(new_n832));
  OR3_X1    g407(.A1(new_n831), .A2(G29), .A3(G33), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT25), .Z(new_n835));
  AOI22_X1  g410(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n836));
  INV_X1    g411(.A(G139), .ZN(new_n837));
  OAI221_X1 g412(.A(new_n835), .B1(new_n464), .B2(new_n836), .C1(new_n484), .C2(new_n837), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT87), .Z(new_n839));
  OAI211_X1 g414(.A(new_n832), .B(new_n833), .C1(new_n839), .C2(new_n718), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(G2072), .Z(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n810), .A2(new_n811), .A3(new_n830), .A4(new_n842), .ZN(new_n843));
  NOR2_X1   g418(.A1(G29), .A2(G35), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(G162), .B2(G29), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT29), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(G2090), .ZN(new_n847));
  NOR3_X1   g422(.A1(new_n737), .A2(new_n843), .A3(new_n847), .ZN(G311));
  OR2_X1    g423(.A1(new_n735), .A2(new_n736), .ZN(new_n849));
  AND3_X1   g424(.A1(new_n810), .A2(new_n830), .A3(new_n842), .ZN(new_n850));
  INV_X1    g425(.A(new_n847), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n849), .A2(new_n850), .A3(new_n851), .A4(new_n811), .ZN(G150));
  AOI22_X1  g427(.A1(new_n504), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n853), .A2(new_n506), .ZN(new_n854));
  INV_X1    g429(.A(G55), .ZN(new_n855));
  INV_X1    g430(.A(G93), .ZN(new_n856));
  OAI22_X1  g431(.A1(new_n511), .A2(new_n855), .B1(new_n519), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(G860), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(KEYINPUT37), .Z(new_n861));
  NAND2_X1  g436(.A1(new_n624), .A2(G559), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT38), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT39), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n552), .A2(KEYINPUT95), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT95), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n542), .A2(new_n546), .A3(new_n551), .A4(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n865), .A2(new_n858), .A3(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n858), .B1(new_n865), .B2(new_n867), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n864), .B(new_n871), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n861), .B1(new_n872), .B2(G860), .ZN(G145));
  OAI21_X1  g448(.A(new_n839), .B1(new_n745), .B2(new_n746), .ZN(new_n874));
  INV_X1    g449(.A(new_n746), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n838), .B(KEYINPUT87), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n875), .A2(new_n876), .A3(new_n744), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  OR2_X1    g453(.A1(G106), .A2(G2105), .ZN(new_n879));
  OAI211_X1 g454(.A(new_n879), .B(G2104), .C1(G118), .C2(new_n464), .ZN(new_n880));
  INV_X1    g455(.A(G130), .ZN(new_n881));
  INV_X1    g456(.A(G142), .ZN(new_n882));
  OAI221_X1 g457(.A(new_n880), .B1(new_n481), .B2(new_n881), .C1(new_n882), .C2(new_n484), .ZN(new_n883));
  OR2_X1    g458(.A1(new_n883), .A2(G164), .ZN(new_n884));
  INV_X1    g459(.A(new_n644), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(G164), .ZN(new_n886));
  AND3_X1   g461(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n885), .B1(new_n884), .B2(new_n886), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n878), .A2(new_n889), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n874), .B(new_n877), .C1(new_n888), .C2(new_n887), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n787), .B(new_n724), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n890), .A2(new_n893), .A3(new_n891), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(G160), .B(KEYINPUT96), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(new_n489), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n768), .B(KEYINPUT96), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(G162), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(new_n641), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n902), .A2(new_n641), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(G37), .B1(new_n897), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g482(.A(KEYINPUT97), .B1(new_n904), .B2(new_n905), .ZN(new_n908));
  INV_X1    g483(.A(new_n905), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT97), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n909), .A2(new_n910), .A3(new_n903), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n895), .A2(new_n912), .A3(new_n896), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT98), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n895), .A2(new_n912), .A3(KEYINPUT98), .A4(new_n896), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n907), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(KEYINPUT99), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT99), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n907), .A2(new_n915), .A3(new_n919), .A4(new_n916), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n918), .A2(KEYINPUT40), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(KEYINPUT40), .B1(new_n918), .B2(new_n920), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(G395));
  XNOR2_X1  g498(.A(G303), .B(G288), .ZN(new_n924));
  OR2_X1    g499(.A1(new_n924), .A2(G305), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(G305), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n925), .A2(new_n604), .A3(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n604), .B1(new_n925), .B2(new_n926), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT42), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n930), .B1(KEYINPUT102), .B2(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n871), .B(new_n629), .ZN(new_n933));
  NAND2_X1  g508(.A1(G299), .A2(new_n624), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n615), .A2(new_n570), .A3(new_n575), .A4(new_n578), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n933), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT100), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n934), .A2(new_n939), .A3(new_n935), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n796), .A2(KEYINPUT100), .A3(new_n615), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT41), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT101), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n937), .A2(KEYINPUT41), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n940), .A2(new_n941), .A3(KEYINPUT101), .A4(new_n942), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n938), .B1(new_n933), .B2(new_n948), .ZN(new_n949));
  AND2_X1   g524(.A1(new_n932), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n932), .A2(new_n949), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n931), .A2(KEYINPUT102), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  NOR3_X1   g530(.A1(new_n950), .A2(new_n951), .A3(new_n953), .ZN(new_n956));
  OAI21_X1  g531(.A(G868), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n957), .B1(G868), .B2(new_n858), .ZN(G295));
  OAI21_X1  g533(.A(new_n957), .B1(G868), .B2(new_n858), .ZN(G331));
  NOR2_X1   g534(.A1(G171), .A2(new_n584), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n960), .B1(G286), .B2(G171), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n961), .B1(new_n869), .B2(new_n870), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n865), .A2(new_n867), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n859), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n527), .A2(new_n529), .ZN(new_n965));
  AOI21_X1  g540(.A(KEYINPUT74), .B1(new_n965), .B2(new_n582), .ZN(new_n966));
  NOR4_X1   g541(.A1(new_n527), .A2(new_n529), .A3(new_n532), .A4(new_n585), .ZN(new_n967));
  OAI21_X1  g542(.A(G171), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n960), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n964), .A2(new_n970), .A3(new_n868), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n962), .A2(new_n971), .A3(new_n936), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT103), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n937), .A2(new_n942), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n940), .A2(KEYINPUT41), .A3(new_n941), .ZN(new_n976));
  NOR3_X1   g551(.A1(new_n869), .A2(new_n961), .A3(new_n870), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n970), .B1(new_n964), .B2(new_n868), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n975), .B(new_n976), .C1(new_n977), .C2(new_n978), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n962), .A2(new_n971), .A3(KEYINPUT103), .A4(new_n936), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n974), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(new_n930), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n962), .A2(new_n971), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n948), .A2(new_n983), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n924), .B(G305), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(G290), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(new_n927), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n984), .A2(new_n987), .A3(new_n972), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT43), .ZN(new_n989));
  INV_X1    g564(.A(G37), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n982), .A2(new_n988), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(KEYINPUT104), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n988), .A2(new_n990), .ZN(new_n993));
  INV_X1    g568(.A(new_n972), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n994), .B1(new_n948), .B2(new_n983), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n995), .A2(new_n987), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT43), .B1(new_n993), .B2(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(G37), .B1(new_n995), .B2(new_n987), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT104), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n998), .A2(new_n999), .A3(new_n989), .A4(new_n982), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n992), .A2(new_n997), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT44), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(new_n996), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT43), .B1(new_n1004), .B2(new_n998), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n998), .A2(KEYINPUT43), .A3(new_n982), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT44), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1003), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT105), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT105), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1003), .A2(new_n1010), .A3(new_n1007), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1011), .ZN(G397));
  INV_X1    g587(.A(G1384), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1013), .B1(new_n495), .B2(new_n502), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT45), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(G160), .A2(G40), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n747), .B(G1996), .ZN(new_n1019));
  INV_X1    g594(.A(G2067), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n787), .B(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n724), .B(new_n726), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1018), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  NOR2_X1   g600(.A1(G290), .A2(G1986), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1026), .A2(KEYINPUT106), .ZN(new_n1027));
  NAND2_X1  g602(.A1(G290), .A2(G1986), .ZN(new_n1028));
  XOR2_X1   g603(.A(new_n1027), .B(new_n1028), .Z(new_n1029));
  AOI21_X1  g604(.A(new_n1025), .B1(new_n1018), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1017), .B1(KEYINPUT50), .B2(new_n1014), .ZN(new_n1031));
  INV_X1    g606(.A(G126), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n474), .A2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(G2105), .B1(new_n1033), .B2(new_n493), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1034), .A2(new_n491), .A3(new_n500), .A4(new_n501), .ZN(new_n1035));
  XOR2_X1   g610(.A(KEYINPUT108), .B(KEYINPUT50), .Z(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(new_n1013), .A3(new_n1036), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1031), .A2(KEYINPUT113), .A3(new_n770), .A4(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT113), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1014), .A2(KEYINPUT50), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n766), .A2(new_n767), .A3(G40), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1040), .A2(new_n1037), .A3(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1039), .B1(new_n1042), .B2(G2084), .ZN(new_n1043));
  OAI211_X1 g618(.A(KEYINPUT45), .B(new_n1013), .C1(new_n495), .C2(new_n502), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1016), .A2(new_n1041), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(new_n821), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1038), .A2(new_n1043), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(G8), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT121), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT51), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n584), .A2(G8), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1048), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1055));
  OAI211_X1 g630(.A(G8), .B(new_n1051), .C1(new_n1047), .C2(new_n584), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1047), .A2(G8), .A3(new_n584), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1045), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT124), .B1(new_n1061), .B2(G2078), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1060), .B(new_n1062), .C1(KEYINPUT124), .C2(G2078), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1044), .A2(KEYINPUT107), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(new_n1016), .ZN(new_n1065));
  INV_X1    g640(.A(G2078), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1014), .A2(KEYINPUT107), .A3(new_n1015), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1065), .A2(new_n1066), .A3(new_n1041), .A4(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(new_n1061), .ZN(new_n1069));
  INV_X1    g644(.A(G1961), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1042), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT123), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT123), .B1(new_n1042), .B2(new_n1070), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1063), .B(new_n1069), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(G171), .ZN(new_n1076));
  NOR3_X1   g651(.A1(new_n1045), .A2(new_n1061), .A3(G2078), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1077), .B1(new_n1068), .B2(new_n1061), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1078), .A2(G301), .A3(new_n1071), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1076), .A2(KEYINPUT54), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1059), .A2(new_n1080), .ZN(new_n1081));
  XNOR2_X1  g656(.A(KEYINPUT122), .B(KEYINPUT54), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1075), .A2(G171), .ZN(new_n1083));
  AOI21_X1  g658(.A(G301), .B1(new_n1078), .B2(new_n1071), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1082), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT52), .ZN(new_n1086));
  INV_X1    g661(.A(G8), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1014), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1087), .B1(new_n1088), .B2(new_n1041), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n705), .A2(G1976), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1086), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(G1976), .ZN(new_n1092));
  NAND2_X1  g667(.A1(G288), .A2(new_n1092), .ZN(new_n1093));
  AND4_X1   g668(.A1(new_n1086), .A2(new_n1089), .A3(new_n1090), .A4(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(G1981), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n597), .A2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(G1981), .B1(new_n593), .B2(new_n596), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT49), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1096), .A2(KEYINPUT49), .A3(new_n1097), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1100), .A2(new_n1089), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(KEYINPUT110), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT110), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1100), .A2(new_n1089), .A3(new_n1104), .A4(new_n1101), .ZN(new_n1105));
  AOI211_X1 g680(.A(new_n1091), .B(new_n1094), .C1(new_n1103), .C2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1042), .A2(G2090), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1065), .A2(new_n1041), .A3(new_n1067), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1107), .B1(new_n702), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1110), .A2(KEYINPUT55), .ZN(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n1112));
  NAND2_X1  g687(.A1(G303), .A2(G8), .ZN(new_n1113));
  MUX2_X1   g688(.A(new_n1111), .B(new_n1112), .S(new_n1113), .Z(new_n1114));
  NOR3_X1   g689(.A1(new_n1109), .A2(new_n1087), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1041), .B1(new_n1014), .B2(KEYINPUT50), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1036), .B1(new_n1035), .B2(new_n1013), .ZN(new_n1118));
  NOR3_X1   g693(.A1(new_n1117), .A2(new_n1118), .A3(G2090), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1119), .B1(new_n1108), .B2(new_n702), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1114), .B1(new_n1120), .B2(new_n1087), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(KEYINPUT112), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT112), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n1123), .B(new_n1114), .C1(new_n1120), .C2(new_n1087), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1085), .A2(new_n1106), .A3(new_n1116), .A4(new_n1125), .ZN(new_n1126));
  AND2_X1   g701(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT117), .ZN(new_n1128));
  INV_X1    g703(.A(G1996), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1127), .A2(new_n1128), .A3(new_n1129), .A4(new_n1041), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1065), .A2(new_n1129), .A3(new_n1041), .A4(new_n1067), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(KEYINPUT117), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1088), .A2(new_n1041), .ZN(new_n1134));
  XOR2_X1   g709(.A(KEYINPUT58), .B(G1341), .Z(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(KEYINPUT118), .B1(new_n1133), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT118), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1136), .ZN(new_n1139));
  AOI211_X1 g714(.A(new_n1138), .B(new_n1139), .C1(new_n1130), .C2(new_n1132), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1137), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT119), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1142), .A2(KEYINPUT59), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1142), .A2(KEYINPUT59), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1141), .A2(new_n553), .A3(new_n1144), .A4(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(G1348), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1042), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1088), .A2(new_n1020), .A3(new_n1041), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT60), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n624), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1148), .A2(KEYINPUT60), .A3(new_n615), .A4(new_n1149), .ZN(new_n1153));
  AOI22_X1  g728(.A1(new_n1152), .A2(new_n1153), .B1(new_n1151), .B2(new_n1150), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT61), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1155), .A2(KEYINPUT120), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT57), .ZN(new_n1157));
  NOR2_X1   g732(.A1(G299), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(KEYINPUT116), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT116), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n576), .A2(new_n577), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n1161), .B(KEYINPUT115), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(new_n575), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1160), .B1(new_n1163), .B2(new_n1157), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1159), .B1(new_n1164), .B2(new_n1158), .ZN(new_n1165));
  INV_X1    g740(.A(G1956), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1166), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1167));
  XNOR2_X1  g742(.A(KEYINPUT56), .B(G2072), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1127), .A2(new_n1041), .A3(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1165), .A2(new_n1167), .A3(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1170), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1165), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1156), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1170), .B1(KEYINPUT120), .B2(new_n1155), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1154), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  AND2_X1   g750(.A1(new_n1131), .A2(KEYINPUT117), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1131), .A2(KEYINPUT117), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1136), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(new_n1138), .ZN(new_n1179));
  OAI211_X1 g754(.A(KEYINPUT118), .B(new_n1136), .C1(new_n1176), .C2(new_n1177), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1179), .A2(new_n553), .A3(new_n1145), .A4(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1181), .A2(new_n1143), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1146), .A2(new_n1175), .A3(new_n1182), .ZN(new_n1183));
  AND2_X1   g758(.A1(new_n1170), .A2(new_n1150), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1172), .B1(new_n1184), .B2(new_n624), .ZN(new_n1185));
  AOI211_X1 g760(.A(new_n1081), .B(new_n1126), .C1(new_n1183), .C2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1059), .A2(KEYINPUT62), .ZN(new_n1187));
  AND3_X1   g762(.A1(new_n1125), .A2(new_n1106), .A3(new_n1116), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT62), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1057), .A2(new_n1189), .A3(new_n1058), .ZN(new_n1190));
  NAND4_X1  g765(.A1(new_n1187), .A2(new_n1188), .A3(new_n1084), .A4(new_n1190), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT63), .ZN(new_n1192));
  NAND4_X1  g767(.A1(new_n1047), .A2(new_n1192), .A3(G8), .A4(new_n621), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1193), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1106), .B1(new_n1194), .B2(new_n1115), .ZN(new_n1195));
  XNOR2_X1  g770(.A(new_n1089), .B(KEYINPUT111), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1197), .A2(new_n1092), .A3(new_n705), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1196), .B1(new_n1198), .B2(new_n1096), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n1048), .A2(G286), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1114), .B1(new_n1109), .B2(new_n1087), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1200), .A2(new_n1106), .A3(new_n1201), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1199), .B1(new_n1202), .B2(KEYINPUT63), .ZN(new_n1203));
  AND3_X1   g778(.A1(new_n1195), .A2(new_n1203), .A3(KEYINPUT114), .ZN(new_n1204));
  AOI21_X1  g779(.A(KEYINPUT114), .B1(new_n1195), .B2(new_n1203), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1191), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1030), .B1(new_n1186), .B2(new_n1206), .ZN(new_n1207));
  XNOR2_X1  g782(.A(new_n1024), .B(KEYINPUT126), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1018), .A2(new_n1026), .ZN(new_n1209));
  XNOR2_X1  g784(.A(new_n1209), .B(KEYINPUT127), .ZN(new_n1210));
  XNOR2_X1  g785(.A(new_n1210), .B(KEYINPUT48), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1208), .A2(new_n1211), .ZN(new_n1212));
  OR2_X1    g787(.A1(new_n724), .A2(new_n726), .ZN(new_n1213));
  AOI21_X1  g788(.A(new_n1213), .B1(new_n1022), .B2(new_n1018), .ZN(new_n1214));
  NOR2_X1   g789(.A1(new_n787), .A2(G2067), .ZN(new_n1215));
  OR3_X1    g790(.A1(new_n1214), .A2(KEYINPUT125), .A3(new_n1215), .ZN(new_n1216));
  OAI21_X1  g791(.A(KEYINPUT125), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1217));
  NAND3_X1  g792(.A1(new_n1216), .A2(new_n1018), .A3(new_n1217), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1018), .A2(new_n1129), .ZN(new_n1219));
  XOR2_X1   g794(.A(new_n1219), .B(KEYINPUT46), .Z(new_n1220));
  NAND2_X1  g795(.A1(new_n747), .A2(new_n1021), .ZN(new_n1221));
  AOI21_X1  g796(.A(new_n1220), .B1(new_n1221), .B2(new_n1018), .ZN(new_n1222));
  XOR2_X1   g797(.A(new_n1222), .B(KEYINPUT47), .Z(new_n1223));
  AND3_X1   g798(.A1(new_n1212), .A2(new_n1218), .A3(new_n1223), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1207), .A2(new_n1224), .ZN(G329));
  assign    G231 = 1'b0;
  AND2_X1   g800(.A1(new_n917), .A2(G319), .ZN(new_n1227));
  NOR2_X1   g801(.A1(G401), .A2(G229), .ZN(new_n1228));
  NAND4_X1  g802(.A1(new_n1227), .A2(new_n677), .A3(new_n1001), .A4(new_n1228), .ZN(G225));
  INV_X1    g803(.A(G225), .ZN(G308));
endmodule


