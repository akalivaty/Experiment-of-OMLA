//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 0 1 0 0 0 1 0 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 1 1 1 0 0 0 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 1 0 1 1 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:25 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  OR3_X1    g003(.A1(new_n189), .A2(KEYINPUT78), .A3(G107), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT78), .B1(new_n189), .B2(G107), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT77), .B(G107), .ZN(new_n192));
  OAI211_X1 g006(.A(new_n190), .B(new_n191), .C1(new_n192), .C2(G104), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G101), .ZN(new_n194));
  INV_X1    g008(.A(G113), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT2), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT2), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G113), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(G116), .B(G119), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n189), .A2(KEYINPUT3), .ZN(new_n202));
  INV_X1    g016(.A(G107), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT77), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT77), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G107), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n202), .A2(new_n204), .A3(new_n206), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT3), .B1(new_n189), .B2(G107), .ZN(new_n208));
  AOI21_X1  g022(.A(G101), .B1(new_n189), .B2(G107), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G119), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G116), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT5), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G116), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G119), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n212), .A2(new_n217), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n215), .B(G113), .C1(new_n218), .C2(new_n214), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n194), .A2(new_n201), .A3(new_n210), .A4(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(G110), .B(G122), .ZN(new_n221));
  INV_X1    g035(.A(G101), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n223), .B1(G104), .B2(new_n203), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n224), .B1(new_n192), .B2(new_n202), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n189), .A2(G107), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n222), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n210), .A2(KEYINPUT4), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n207), .A2(new_n208), .A3(new_n226), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n222), .A2(KEYINPUT4), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT2), .B(G113), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n218), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(new_n201), .A3(KEYINPUT67), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT67), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n218), .A2(new_n233), .A3(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n232), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n220), .B(new_n221), .C1(new_n229), .C2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT79), .ZN(new_n240));
  AND2_X1   g054(.A1(new_n235), .A2(new_n237), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n230), .A2(G101), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n242), .A2(KEYINPUT4), .A3(new_n210), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n241), .A2(new_n243), .A3(new_n232), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT79), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n244), .A2(new_n245), .A3(new_n220), .A4(new_n221), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n240), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT6), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n244), .A2(new_n220), .ZN(new_n249));
  INV_X1    g063(.A(new_n221), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT80), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n247), .A2(new_n251), .A3(KEYINPUT80), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n249), .A2(new_n248), .A3(new_n250), .ZN(new_n256));
  INV_X1    g070(.A(G128), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n257), .A2(KEYINPUT1), .ZN(new_n258));
  INV_X1    g072(.A(G146), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G143), .ZN(new_n260));
  INV_X1    g074(.A(G143), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G146), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n258), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n261), .A2(G146), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT64), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n265), .B1(new_n259), .B2(G143), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n261), .A2(KEYINPUT64), .A3(G146), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n264), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n257), .B1(new_n260), .B2(KEYINPUT1), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n263), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  OR2_X1    g084(.A1(new_n270), .A2(G125), .ZN(new_n271));
  AND2_X1   g085(.A1(KEYINPUT0), .A2(G128), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n260), .A2(new_n262), .A3(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(KEYINPUT0), .A2(G128), .ZN(new_n274));
  OR2_X1    g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n273), .B1(new_n268), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G125), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n271), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G953), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G224), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n278), .B(new_n281), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n254), .A2(new_n255), .A3(new_n256), .A4(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT81), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n256), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n286), .B1(new_n252), .B2(new_n253), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n287), .A2(KEYINPUT81), .A3(new_n255), .A4(new_n282), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  XOR2_X1   g103(.A(new_n221), .B(KEYINPUT8), .Z(new_n290));
  AND2_X1   g104(.A1(new_n194), .A2(new_n210), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n219), .A2(new_n201), .ZN(new_n292));
  OR2_X1    g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n290), .B1(new_n293), .B2(new_n220), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT7), .ZN(new_n295));
  NOR3_X1   g109(.A1(new_n278), .A2(new_n295), .A3(new_n281), .ZN(new_n296));
  AOI22_X1  g110(.A1(new_n271), .A2(new_n277), .B1(KEYINPUT7), .B2(new_n280), .ZN(new_n297));
  NOR3_X1   g111(.A1(new_n294), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(G902), .B1(new_n298), .B2(new_n247), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n289), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(G210), .B1(G237), .B2(G902), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n289), .A2(new_n301), .A3(new_n299), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n188), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  AND3_X1   g119(.A1(new_n261), .A2(KEYINPUT64), .A3(G146), .ZN(new_n306));
  AOI21_X1  g120(.A(KEYINPUT64), .B1(new_n261), .B2(G146), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n260), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n272), .A2(new_n274), .ZN(new_n309));
  AND2_X1   g123(.A1(new_n260), .A2(new_n262), .ZN(new_n310));
  AOI22_X1  g124(.A1(new_n308), .A2(new_n309), .B1(new_n310), .B2(new_n272), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n243), .A2(new_n311), .A3(new_n232), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n263), .B1(new_n310), .B2(new_n269), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n194), .A2(new_n210), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT10), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G134), .ZN(new_n317));
  OAI21_X1  g131(.A(KEYINPUT11), .B1(new_n317), .B2(G137), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT11), .ZN(new_n319));
  INV_X1    g133(.A(G137), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(new_n320), .A3(G134), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  XOR2_X1   g136(.A(KEYINPUT65), .B(G131), .Z(new_n323));
  OAI21_X1  g137(.A(KEYINPUT66), .B1(new_n320), .B2(G134), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT66), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n325), .A2(new_n317), .A3(G137), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NOR3_X1   g141(.A1(new_n322), .A2(new_n323), .A3(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G131), .ZN(new_n329));
  AND2_X1   g143(.A1(new_n324), .A2(new_n326), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n318), .A2(new_n321), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n194), .A2(KEYINPUT10), .A3(new_n270), .A4(new_n210), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n312), .A2(new_n316), .A3(new_n333), .A4(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n314), .B1(new_n291), .B2(new_n270), .ZN(new_n336));
  INV_X1    g150(.A(new_n333), .ZN(new_n337));
  AND3_X1   g151(.A1(new_n336), .A2(KEYINPUT12), .A3(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(KEYINPUT12), .B1(new_n336), .B2(new_n337), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n335), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(G110), .B(G140), .ZN(new_n341));
  AND2_X1   g155(.A1(new_n279), .A2(G227), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n341), .B(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n312), .A2(new_n316), .A3(new_n334), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(new_n337), .ZN(new_n345));
  INV_X1    g159(.A(new_n343), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n335), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  AOI22_X1  g162(.A1(new_n340), .A2(new_n343), .B1(new_n345), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(G469), .B1(new_n349), .B2(G902), .ZN(new_n350));
  INV_X1    g164(.A(G469), .ZN(new_n351));
  INV_X1    g165(.A(G902), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n336), .A2(new_n337), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT12), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n336), .A2(KEYINPUT12), .A3(new_n337), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n347), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n346), .B1(new_n345), .B2(new_n335), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n351), .B(new_n352), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n350), .A2(new_n359), .ZN(new_n360));
  XNOR2_X1  g174(.A(KEYINPUT9), .B(G234), .ZN(new_n361));
  OAI21_X1  g175(.A(G221), .B1(new_n361), .B2(G902), .ZN(new_n362));
  XOR2_X1   g176(.A(new_n362), .B(KEYINPUT76), .Z(new_n363));
  NAND2_X1  g177(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT84), .ZN(new_n366));
  XNOR2_X1  g180(.A(G113), .B(G122), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n367), .B(new_n189), .ZN(new_n368));
  NOR2_X1   g182(.A1(G237), .A2(G953), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n369), .A2(G143), .A3(G214), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(G143), .B1(new_n369), .B2(G214), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n323), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G237), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(new_n279), .A3(G214), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n261), .ZN(new_n376));
  XNOR2_X1  g190(.A(KEYINPUT65), .B(G131), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n376), .A2(new_n377), .A3(new_n370), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(G125), .B(G140), .ZN(new_n380));
  AOI21_X1  g194(.A(KEYINPUT19), .B1(new_n380), .B2(KEYINPUT82), .ZN(new_n381));
  INV_X1    g195(.A(G140), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G125), .ZN(new_n383));
  INV_X1    g197(.A(G125), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G140), .ZN(new_n385));
  AND4_X1   g199(.A1(KEYINPUT82), .A2(new_n383), .A3(new_n385), .A4(KEYINPUT19), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n259), .B1(new_n381), .B2(new_n386), .ZN(new_n387));
  NOR3_X1   g201(.A1(new_n384), .A2(KEYINPUT16), .A3(G140), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n388), .B1(new_n380), .B2(KEYINPUT16), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G146), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n379), .A2(new_n387), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n376), .A2(new_n370), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(KEYINPUT18), .A3(G131), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n380), .B(new_n259), .ZN(new_n394));
  NAND2_X1  g208(.A1(KEYINPUT18), .A2(G131), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n376), .A2(new_n370), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n393), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n368), .B1(new_n391), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(KEYINPUT83), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n379), .A2(KEYINPUT17), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n392), .A2(KEYINPUT17), .A3(new_n323), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT16), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n403), .A2(new_n382), .A3(G125), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n383), .A2(new_n385), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n404), .B1(new_n405), .B2(new_n403), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n259), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n402), .A2(new_n407), .A3(new_n390), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n368), .B(new_n397), .C1(new_n401), .C2(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n409), .B1(new_n398), .B2(KEYINPUT83), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n366), .B1(new_n400), .B2(new_n410), .ZN(new_n411));
  NOR2_X1   g225(.A1(G475), .A2(G902), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT83), .ZN(new_n413));
  AND2_X1   g227(.A1(new_n391), .A2(new_n397), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n413), .B1(new_n414), .B2(new_n368), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n415), .A2(KEYINPUT84), .A3(new_n399), .A4(new_n409), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n411), .A2(new_n412), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(KEYINPUT20), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT85), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n417), .A2(KEYINPUT85), .A3(KEYINPUT20), .ZN(new_n421));
  NOR3_X1   g235(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n422), .B1(new_n400), .B2(new_n410), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n420), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n397), .B1(new_n401), .B2(new_n408), .ZN(new_n425));
  INV_X1    g239(.A(new_n368), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n409), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n352), .ZN(new_n429));
  AND2_X1   g243(.A1(new_n429), .A2(G475), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n424), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(G952), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n433), .A2(KEYINPUT88), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n433), .A2(KEYINPUT88), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n279), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(G234), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n437), .B1(new_n438), .B2(new_n374), .ZN(new_n439));
  OAI211_X1 g253(.A(G902), .B(G953), .C1(new_n438), .C2(new_n374), .ZN(new_n440));
  XOR2_X1   g254(.A(new_n440), .B(KEYINPUT89), .Z(new_n441));
  XOR2_X1   g255(.A(KEYINPUT21), .B(G898), .Z(new_n442));
  OAI21_X1  g256(.A(new_n439), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  XOR2_X1   g257(.A(new_n443), .B(KEYINPUT90), .Z(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n192), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n216), .A2(G122), .ZN(new_n447));
  INV_X1    g261(.A(G122), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(G116), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n446), .A2(new_n450), .ZN(new_n451));
  OR2_X1    g265(.A1(new_n447), .A2(KEYINPUT14), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n447), .A2(KEYINPUT14), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n452), .A2(new_n453), .A3(new_n449), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n451), .B1(G107), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(KEYINPUT86), .B1(new_n257), .B2(G143), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT86), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n457), .A2(new_n261), .A3(G128), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n459), .B1(G128), .B2(new_n261), .ZN(new_n460));
  AND2_X1   g274(.A1(new_n460), .A2(G134), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n460), .A2(G134), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n455), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT87), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n455), .B(KEYINPUT87), .C1(new_n461), .C2(new_n462), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n451), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n446), .A2(new_n450), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n462), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n459), .ZN(new_n471));
  OAI22_X1  g285(.A1(new_n471), .A2(KEYINPUT13), .B1(G128), .B2(new_n261), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n472), .B1(KEYINPUT13), .B2(new_n471), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n470), .B1(new_n473), .B2(new_n317), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n467), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(G217), .ZN(new_n476));
  NOR3_X1   g290(.A1(new_n361), .A2(new_n476), .A3(G953), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n477), .B1(new_n467), .B2(new_n474), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n352), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(G478), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n482), .A2(KEYINPUT15), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n481), .B(new_n483), .ZN(new_n484));
  NOR3_X1   g298(.A1(new_n432), .A2(new_n445), .A3(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n305), .A2(new_n365), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n476), .B1(G234), .B2(new_n352), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n279), .A2(G221), .A3(G234), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n489), .B(KEYINPUT73), .ZN(new_n490));
  XNOR2_X1  g304(.A(KEYINPUT22), .B(G137), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n490), .B(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT23), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n493), .B1(new_n211), .B2(G128), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n257), .A2(KEYINPUT23), .A3(G119), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n494), .B(new_n495), .C1(G119), .C2(new_n257), .ZN(new_n496));
  XNOR2_X1  g310(.A(G119), .B(G128), .ZN(new_n497));
  XOR2_X1   g311(.A(KEYINPUT24), .B(G110), .Z(new_n498));
  OAI22_X1  g312(.A1(new_n496), .A2(G110), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n499), .B(new_n390), .C1(G146), .C2(new_n405), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n496), .A2(G110), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT72), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n496), .A2(KEYINPUT72), .A3(G110), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n498), .A2(new_n497), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n406), .A2(new_n259), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n389), .A2(G146), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OAI211_X1 g323(.A(KEYINPUT74), .B(new_n500), .C1(new_n505), .C2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n503), .A2(new_n504), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n407), .A2(new_n390), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n512), .A2(new_n506), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(KEYINPUT74), .B1(new_n514), .B2(new_n500), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n492), .B1(new_n511), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n500), .B1(new_n505), .B2(new_n509), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT74), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n492), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n516), .A2(new_n352), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT25), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n517), .A2(new_n518), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n510), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n519), .B1(new_n525), .B2(new_n492), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n526), .A2(KEYINPUT25), .A3(new_n352), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n488), .B1(new_n523), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n487), .A2(G902), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n529), .B(KEYINPUT75), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n528), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(G472), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT29), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n311), .B1(new_n328), .B2(new_n332), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT30), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n330), .A2(new_n377), .A3(new_n331), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n317), .A2(G137), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n320), .A2(G134), .ZN(new_n541));
  OAI21_X1  g355(.A(G131), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n270), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n537), .A2(new_n538), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n538), .B1(new_n537), .B2(new_n543), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n241), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n235), .A2(new_n237), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n537), .A2(new_n543), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n369), .A2(G210), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n549), .B(KEYINPUT27), .ZN(new_n550));
  XNOR2_X1  g364(.A(KEYINPUT26), .B(G101), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n550), .B(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n546), .A2(new_n548), .A3(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  AND3_X1   g369(.A1(new_n537), .A2(new_n543), .A3(new_n547), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n547), .B1(new_n537), .B2(new_n543), .ZN(new_n557));
  OAI21_X1  g371(.A(KEYINPUT28), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT28), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n548), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n553), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n536), .B1(new_n555), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n558), .A2(new_n560), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n552), .A2(KEYINPUT29), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n352), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n535), .B1(new_n562), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n548), .A2(new_n552), .ZN(new_n568));
  AND3_X1   g382(.A1(new_n270), .A2(new_n539), .A3(new_n542), .ZN(new_n569));
  OAI21_X1  g383(.A(G131), .B1(new_n322), .B2(new_n327), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n276), .B1(new_n539), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(KEYINPUT30), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n537), .A2(new_n538), .A3(new_n543), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n568), .B1(new_n574), .B2(new_n241), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT31), .ZN(new_n576));
  AOI22_X1  g390(.A1(new_n563), .A2(new_n553), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n568), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n546), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(KEYINPUT68), .B1(new_n579), .B2(KEYINPUT31), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT68), .ZN(new_n581));
  AOI211_X1 g395(.A(new_n581), .B(new_n576), .C1(new_n546), .C2(new_n578), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n577), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n535), .A2(new_n352), .A3(KEYINPUT69), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT69), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n585), .B1(G472), .B2(G902), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT32), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n567), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT71), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n241), .B1(new_n569), .B2(new_n571), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n559), .B1(new_n592), .B2(new_n548), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n548), .A2(new_n559), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n553), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n546), .A2(new_n576), .A3(new_n578), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n547), .B1(new_n572), .B2(new_n573), .ZN(new_n598));
  OAI21_X1  g412(.A(KEYINPUT31), .B1(new_n598), .B2(new_n568), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n581), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n579), .A2(KEYINPUT68), .A3(KEYINPUT31), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n597), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n587), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(new_n589), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  OAI21_X1  g419(.A(KEYINPUT70), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT70), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n583), .A2(new_n607), .A3(new_n604), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n590), .A2(new_n591), .A3(new_n606), .A4(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n606), .A2(new_n608), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n563), .A2(new_n552), .ZN(new_n611));
  AOI21_X1  g425(.A(KEYINPUT29), .B1(new_n611), .B2(new_n554), .ZN(new_n612));
  OAI21_X1  g426(.A(G472), .B1(new_n612), .B2(new_n565), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n600), .A2(new_n601), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n603), .B1(new_n614), .B2(new_n577), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n613), .B1(new_n615), .B2(KEYINPUT32), .ZN(new_n616));
  OAI21_X1  g430(.A(KEYINPUT71), .B1(new_n610), .B2(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n534), .B1(new_n609), .B2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n486), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(new_n222), .ZN(G3));
  OAI21_X1  g435(.A(G472), .B1(new_n602), .B2(G902), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n588), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n534), .A2(new_n364), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(KEYINPUT91), .ZN(new_n625));
  NAND2_X1  g439(.A1(KEYINPUT92), .A2(KEYINPUT33), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n626), .B1(new_n479), .B2(new_n480), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n482), .A2(G902), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n475), .B(new_n478), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT92), .B(KEYINPUT33), .Z(new_n630));
  OAI211_X1 g444(.A(new_n627), .B(new_n628), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT93), .B(G478), .Z(new_n632));
  NAND2_X1  g446(.A1(new_n481), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n432), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n635), .A2(new_n445), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n625), .A2(new_n305), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(KEYINPUT94), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT34), .B(G104), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G6));
  AND2_X1   g454(.A1(new_n411), .A2(new_n416), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n422), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n420), .A2(new_n421), .A3(new_n642), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n643), .A2(new_n444), .A3(new_n484), .A4(new_n431), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n305), .A2(new_n645), .A3(KEYINPUT95), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT95), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n301), .B1(new_n289), .B2(new_n299), .ZN(new_n648));
  INV_X1    g462(.A(new_n299), .ZN(new_n649));
  AOI211_X1 g463(.A(new_n302), .B(new_n649), .C1(new_n285), .C2(new_n288), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n187), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n647), .B1(new_n651), .B2(new_n644), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n646), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n625), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT35), .B(G107), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G9));
  AOI21_X1  g470(.A(KEYINPUT25), .B1(new_n526), .B2(new_n352), .ZN(new_n657));
  AND4_X1   g471(.A1(KEYINPUT25), .A2(new_n516), .A3(new_n352), .A4(new_n520), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n487), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n492), .A2(KEYINPUT36), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n517), .B(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n530), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n663), .A2(new_n588), .A3(new_n622), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n486), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT96), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT37), .B(G110), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G12));
  AND2_X1   g482(.A1(new_n661), .A2(new_n530), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n528), .A2(new_n669), .ZN(new_n670));
  AOI211_X1 g484(.A(new_n364), .B(new_n670), .C1(new_n609), .C2(new_n617), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n303), .A2(new_n304), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n439), .B(KEYINPUT97), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n673), .B1(G900), .B2(new_n441), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n643), .A2(new_n431), .A3(new_n484), .A4(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n672), .A2(KEYINPUT98), .A3(new_n187), .A4(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT98), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n678), .B1(new_n651), .B2(new_n675), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n671), .A2(new_n677), .A3(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT99), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n671), .A2(new_n679), .A3(new_n677), .A4(KEYINPUT99), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G128), .ZN(G30));
  XOR2_X1   g499(.A(new_n672), .B(KEYINPUT38), .Z(new_n686));
  NAND3_X1  g500(.A1(new_n592), .A2(new_n548), .A3(new_n553), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n352), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n552), .B1(new_n598), .B2(new_n556), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n535), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n692), .B1(new_n615), .B2(KEYINPUT32), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n610), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n483), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n481), .B(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n697), .B1(new_n424), .B2(new_n431), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n695), .A2(new_n187), .A3(new_n670), .A4(new_n698), .ZN(new_n699));
  OR2_X1    g513(.A1(new_n686), .A2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT100), .ZN(new_n701));
  OR2_X1    g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n674), .B(KEYINPUT39), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n365), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g519(.A(new_n705), .B(KEYINPUT40), .Z(new_n706));
  NAND3_X1  g520(.A1(new_n702), .A2(new_n703), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G143), .ZN(G45));
  INV_X1    g522(.A(KEYINPUT101), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n432), .A2(new_n634), .A3(new_n674), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n709), .B1(new_n305), .B2(new_n711), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n670), .B1(new_n609), .B2(new_n617), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n365), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n305), .A2(new_n711), .A3(new_n709), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G146), .ZN(G48));
  NOR2_X1   g532(.A1(new_n357), .A2(new_n358), .ZN(new_n719));
  OAI21_X1  g533(.A(G469), .B1(new_n719), .B2(G902), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n720), .A2(new_n362), .A3(new_n359), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(KEYINPUT102), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT102), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n720), .A2(new_n723), .A3(new_n362), .A4(new_n359), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n618), .A2(new_n305), .A3(new_n636), .A4(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(KEYINPUT41), .B(G113), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G15));
  NAND2_X1  g542(.A1(new_n618), .A2(new_n725), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n729), .B1(new_n652), .B2(new_n646), .ZN(new_n730));
  XNOR2_X1  g544(.A(KEYINPUT103), .B(G116), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n730), .B(new_n731), .ZN(G18));
  INV_X1    g546(.A(new_n721), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n713), .A2(new_n305), .A3(new_n485), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G119), .ZN(G21));
  OAI211_X1 g549(.A(new_n698), .B(new_n187), .C1(new_n648), .C2(new_n650), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g551(.A(KEYINPUT105), .B1(new_n528), .B2(new_n532), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT105), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n659), .A2(new_n739), .A3(new_n531), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n577), .A2(new_n599), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n587), .B(KEYINPUT104), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n622), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n741), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n722), .A2(new_n444), .A3(new_n724), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n737), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G122), .ZN(G24));
  NAND2_X1  g564(.A1(new_n745), .A2(new_n663), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n710), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(new_n305), .A3(new_n733), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G125), .ZN(G27));
  AND2_X1   g568(.A1(new_n631), .A2(new_n633), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n755), .B1(new_n424), .B2(new_n431), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n590), .B1(new_n602), .B2(new_n605), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n756), .A2(new_n757), .A3(new_n674), .A4(new_n741), .ZN(new_n758));
  INV_X1    g572(.A(new_n362), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n759), .B1(new_n350), .B2(new_n359), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n303), .A2(new_n187), .A3(new_n304), .A4(new_n760), .ZN(new_n761));
  OAI21_X1  g575(.A(KEYINPUT42), .B1(new_n758), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n360), .A2(new_n362), .ZN(new_n763));
  NOR4_X1   g577(.A1(new_n648), .A2(new_n650), .A3(new_n188), .A4(new_n763), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n710), .A2(KEYINPUT42), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n764), .A2(new_n618), .A3(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT106), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n762), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n767), .B1(new_n762), .B2(new_n766), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G131), .ZN(G33));
  NAND3_X1  g585(.A1(new_n764), .A2(new_n618), .A3(new_n676), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G134), .ZN(G36));
  AND2_X1   g587(.A1(new_n349), .A2(KEYINPUT45), .ZN(new_n774));
  OAI21_X1  g588(.A(G469), .B1(new_n349), .B2(KEYINPUT45), .ZN(new_n775));
  OR2_X1    g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(G469), .A2(G902), .ZN(new_n777));
  AOI21_X1  g591(.A(KEYINPUT46), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n776), .A2(KEYINPUT46), .A3(new_n777), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n359), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n778), .B1(new_n780), .B2(KEYINPUT107), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n781), .B1(KEYINPUT107), .B2(new_n780), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n782), .A2(new_n362), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT108), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n783), .A2(new_n784), .A3(new_n704), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n782), .A2(new_n362), .A3(new_n704), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(KEYINPUT108), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n648), .A2(new_n650), .A3(new_n188), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(KEYINPUT109), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n424), .A2(new_n431), .A3(new_n634), .ZN(new_n791));
  XOR2_X1   g605(.A(new_n791), .B(KEYINPUT43), .Z(new_n792));
  NAND3_X1  g606(.A1(new_n792), .A2(new_n623), .A3(new_n663), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT44), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n790), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n795), .A2(KEYINPUT110), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(KEYINPUT110), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n793), .A2(new_n794), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n788), .A2(new_n796), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G137), .ZN(G39));
  INV_X1    g614(.A(KEYINPUT111), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT47), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n783), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n609), .A2(new_n617), .A3(new_n534), .ZN(new_n804));
  NOR4_X1   g618(.A1(new_n804), .A2(new_n672), .A3(new_n188), .A4(new_n710), .ZN(new_n805));
  XOR2_X1   g619(.A(new_n805), .B(KEYINPUT112), .Z(new_n806));
  OR2_X1    g620(.A1(new_n801), .A2(KEYINPUT47), .ZN(new_n807));
  AOI22_X1  g621(.A1(new_n782), .A2(new_n362), .B1(new_n807), .B2(new_n802), .ZN(new_n808));
  OR3_X1    g622(.A1(new_n803), .A2(new_n806), .A3(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G140), .ZN(G42));
  INV_X1    g624(.A(new_n791), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n720), .A2(new_n359), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(KEYINPUT49), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n363), .A2(new_n187), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n695), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n686), .A2(new_n741), .A3(new_n811), .A4(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n433), .A2(new_n279), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n634), .B1(new_n424), .B2(new_n431), .ZN(new_n818));
  INV_X1    g632(.A(new_n432), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n818), .B1(new_n819), .B2(new_n697), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n534), .A2(new_n623), .A3(new_n445), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n820), .A2(new_n305), .A3(new_n365), .A4(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n726), .A2(new_n734), .A3(new_n749), .A4(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n486), .B1(new_n619), .B2(new_n664), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n823), .A2(new_n730), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n643), .A2(new_n431), .ZN(new_n826));
  INV_X1    g640(.A(new_n674), .ZN(new_n827));
  NOR4_X1   g641(.A1(new_n826), .A2(new_n364), .A3(new_n484), .A4(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n713), .A2(new_n789), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n764), .A2(new_n752), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n772), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT113), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n772), .A2(new_n829), .A3(new_n830), .A4(KEYINPUT113), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n762), .A2(new_n766), .A3(KEYINPUT53), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n825), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n760), .A2(new_n670), .A3(new_n674), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n694), .A2(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n305), .A2(new_n839), .A3(KEYINPUT115), .A4(new_n698), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT115), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n663), .A2(new_n827), .ZN(new_n842));
  OAI211_X1 g656(.A(new_n842), .B(new_n760), .C1(new_n610), .C2(new_n693), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n841), .B1(new_n736), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n845), .B1(new_n715), .B2(new_n716), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n684), .A2(new_n753), .A3(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT52), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n753), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n850), .B1(new_n682), .B2(new_n683), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n851), .A2(KEYINPUT52), .A3(new_n846), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n837), .B1(new_n849), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n849), .A2(new_n852), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n825), .A2(new_n835), .A3(new_n770), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT114), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n825), .A2(new_n835), .A3(new_n770), .A4(KEYINPUT114), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n854), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  XOR2_X1   g673(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n860));
  AOI211_X1 g674(.A(KEYINPUT54), .B(new_n853), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT53), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n863), .B1(new_n860), .B2(new_n859), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n861), .B1(new_n864), .B2(KEYINPUT54), .ZN(new_n865));
  INV_X1    g679(.A(new_n673), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n792), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n867), .A2(new_n746), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n868), .A2(new_n305), .A3(new_n733), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n789), .A2(new_n733), .ZN(new_n870));
  NOR4_X1   g684(.A1(new_n870), .A2(new_n534), .A3(new_n439), .A4(new_n695), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n436), .B1(new_n871), .B2(new_n756), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n867), .A2(new_n870), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT48), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n757), .A2(new_n741), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n874), .B1(new_n873), .B2(new_n875), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n869), .B(new_n872), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  OAI22_X1  g692(.A1(new_n803), .A2(new_n808), .B1(new_n363), .B2(new_n812), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n879), .A2(new_n790), .A3(new_n868), .ZN(new_n880));
  INV_X1    g694(.A(new_n868), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n686), .A2(new_n188), .A3(new_n733), .ZN(new_n882));
  OAI21_X1  g696(.A(KEYINPUT117), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT50), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OR2_X1    g699(.A1(new_n883), .A2(new_n884), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n867), .A2(new_n751), .A3(new_n870), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n432), .A2(new_n634), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n887), .B1(new_n871), .B2(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n880), .A2(new_n885), .A3(new_n886), .A4(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT51), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n878), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n886), .A2(new_n889), .A3(new_n885), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT118), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n886), .A2(new_n889), .A3(KEYINPUT118), .A4(new_n885), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n895), .A2(KEYINPUT51), .A3(new_n896), .A4(new_n880), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n892), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n865), .A2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT119), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n817), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(KEYINPUT119), .B1(new_n865), .B2(new_n898), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n816), .B1(new_n901), .B2(new_n902), .ZN(G75));
  NAND2_X1  g717(.A1(new_n287), .A2(new_n255), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(new_n282), .ZN(new_n905));
  XNOR2_X1  g719(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n905), .B(new_n906), .Z(new_n907));
  NAND2_X1  g721(.A1(new_n857), .A2(new_n858), .ZN(new_n908));
  INV_X1    g722(.A(new_n852), .ZN(new_n909));
  AOI21_X1  g723(.A(KEYINPUT52), .B1(new_n851), .B2(new_n846), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n860), .B1(new_n908), .B2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n853), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n352), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n914), .A2(G210), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n907), .B1(new_n915), .B2(KEYINPUT56), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n279), .A2(G952), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n915), .A2(KEYINPUT56), .A3(new_n907), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n919), .A2(new_n920), .ZN(G51));
  INV_X1    g735(.A(KEYINPUT121), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n912), .A2(new_n913), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(KEYINPUT54), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT54), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n912), .A2(new_n925), .A3(new_n913), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n777), .B(KEYINPUT57), .Z(new_n928));
  AOI21_X1  g742(.A(new_n719), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  AOI211_X1 g743(.A(new_n352), .B(new_n776), .C1(new_n912), .C2(new_n913), .ZN(new_n930));
  OAI211_X1 g744(.A(new_n922), .B(new_n918), .C1(new_n929), .C2(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n925), .B1(new_n912), .B2(new_n913), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n928), .B1(new_n932), .B2(new_n861), .ZN(new_n933));
  INV_X1    g747(.A(new_n719), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n930), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(KEYINPUT121), .B1(new_n935), .B2(new_n917), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n931), .A2(new_n936), .ZN(G54));
  NAND3_X1  g751(.A1(new_n914), .A2(KEYINPUT58), .A3(G475), .ZN(new_n938));
  INV_X1    g752(.A(new_n641), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n938), .A2(new_n939), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n940), .A2(new_n941), .A3(new_n917), .ZN(G60));
  OAI21_X1  g756(.A(new_n627), .B1(new_n629), .B2(new_n630), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT122), .Z(new_n944));
  INV_X1    g758(.A(new_n865), .ZN(new_n945));
  NAND2_X1  g759(.A1(G478), .A2(G902), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT59), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n944), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n927), .A2(new_n944), .A3(new_n947), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n948), .A2(new_n917), .A3(new_n949), .ZN(G63));
  NAND2_X1  g764(.A1(G217), .A2(G902), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT60), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n952), .B1(new_n912), .B2(new_n913), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(new_n661), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n954), .B(new_n918), .C1(new_n526), .C2(new_n953), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT61), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(G66));
  NAND3_X1  g771(.A1(new_n442), .A2(G224), .A3(G953), .ZN(new_n958));
  INV_X1    g772(.A(new_n825), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n958), .B1(new_n959), .B2(G953), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n904), .B1(G898), .B2(new_n279), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT123), .Z(new_n962));
  XNOR2_X1  g776(.A(new_n960), .B(new_n962), .ZN(G69));
  NAND3_X1  g777(.A1(new_n788), .A2(new_n737), .A3(new_n875), .ZN(new_n964));
  AND4_X1   g778(.A1(new_n770), .A2(new_n809), .A3(new_n772), .A4(new_n964), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n851), .A2(new_n717), .ZN(new_n966));
  AOI21_X1  g780(.A(KEYINPUT126), .B1(new_n799), .B2(new_n966), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n799), .A2(KEYINPUT126), .A3(new_n966), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n965), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n381), .A2(new_n386), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT124), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT125), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(new_n574), .Z(new_n973));
  NOR2_X1   g787(.A1(new_n973), .A2(G953), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n969), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g789(.A(G900), .B1(KEYINPUT127), .B2(G227), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(G953), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT127), .ZN(new_n979));
  NAND2_X1  g793(.A1(G227), .A2(G900), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n979), .B1(new_n980), .B2(G953), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n707), .A2(new_n966), .ZN(new_n983));
  OR2_X1    g797(.A1(new_n983), .A2(KEYINPUT62), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(KEYINPUT62), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n619), .A2(new_n705), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n986), .A2(new_n789), .A3(new_n820), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n809), .A2(new_n799), .A3(new_n987), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n984), .A2(new_n985), .A3(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n973), .B1(new_n989), .B2(G953), .ZN(new_n990));
  AND3_X1   g804(.A1(new_n978), .A2(new_n982), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n982), .B1(new_n978), .B2(new_n990), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n991), .A2(new_n992), .ZN(G72));
  OR2_X1    g807(.A1(new_n969), .A2(new_n959), .ZN(new_n994));
  NAND2_X1  g808(.A1(G472), .A2(G902), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n995), .B(KEYINPUT63), .Z(new_n996));
  AOI21_X1  g810(.A(new_n554), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  AND4_X1   g811(.A1(new_n554), .A2(new_n864), .A3(new_n690), .A4(new_n996), .ZN(new_n998));
  NAND4_X1  g812(.A1(new_n984), .A2(new_n825), .A3(new_n988), .A4(new_n985), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n690), .B1(new_n999), .B2(new_n996), .ZN(new_n1000));
  NOR4_X1   g814(.A1(new_n997), .A2(new_n998), .A3(new_n917), .A4(new_n1000), .ZN(G57));
endmodule


