//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 1 1 0 1 1 0 1 1 0 1 1 1 0 0 0 1 1 0 0 0 1 0 0 0 0 1 1 1 0 0 0 0 1 0 1 0 1 1 1 0 0 0 0 1 0 1 0 0 1 0 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:19 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n608, new_n609, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n634, new_n635, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n843, new_n844, new_n845, new_n846, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT73), .ZN(new_n188));
  INV_X1    g002(.A(G137), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G134), .ZN(new_n190));
  INV_X1    g004(.A(G134), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G137), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n190), .B1(new_n193), .B2(KEYINPUT64), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT64), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n192), .A2(new_n195), .ZN(new_n196));
  OAI21_X1  g010(.A(G131), .B1(new_n194), .B2(new_n196), .ZN(new_n197));
  OR3_X1    g011(.A1(new_n191), .A2(KEYINPUT11), .A3(G137), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT11), .B1(new_n191), .B2(G137), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(new_n193), .ZN(new_n200));
  INV_X1    g014(.A(G131), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n197), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G143), .ZN(new_n205));
  INV_X1    g019(.A(G143), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G128), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT65), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT65), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G128), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT1), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n214), .B1(G143), .B2(new_n204), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n208), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT66), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(G143), .B(G146), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(new_n214), .A3(G128), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT1), .B1(new_n206), .B2(G146), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(new_n210), .A3(new_n212), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n222), .A2(KEYINPUT66), .A3(new_n208), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n218), .A2(new_n220), .A3(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n218), .A2(KEYINPUT68), .A3(new_n220), .A4(new_n223), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n203), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  XOR2_X1   g042(.A(G116), .B(G119), .Z(new_n229));
  XNOR2_X1  g043(.A(KEYINPUT2), .B(G113), .ZN(new_n230));
  XNOR2_X1  g044(.A(new_n229), .B(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n232));
  XNOR2_X1  g046(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(new_n200), .B(new_n201), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT0), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n219), .B1(new_n235), .B2(new_n209), .ZN(new_n236));
  XOR2_X1   g050(.A(KEYINPUT0), .B(G128), .Z(new_n237));
  OAI21_X1  g051(.A(new_n236), .B1(new_n219), .B2(new_n237), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n234), .A2(new_n238), .ZN(new_n239));
  NOR3_X1   g053(.A1(new_n228), .A2(new_n233), .A3(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n241));
  INV_X1    g055(.A(G237), .ZN(new_n242));
  INV_X1    g056(.A(G953), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n242), .A2(new_n243), .A3(G210), .ZN(new_n244));
  XNOR2_X1  g058(.A(new_n241), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g059(.A(KEYINPUT26), .B(G101), .ZN(new_n246));
  XNOR2_X1  g060(.A(new_n245), .B(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(KEYINPUT70), .B1(new_n240), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n203), .ZN(new_n250));
  AND3_X1   g064(.A1(new_n222), .A2(KEYINPUT66), .A3(new_n208), .ZN(new_n251));
  AOI21_X1  g065(.A(KEYINPUT66), .B1(new_n222), .B2(new_n208), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(KEYINPUT68), .B1(new_n253), .B2(new_n220), .ZN(new_n254));
  INV_X1    g068(.A(new_n227), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n250), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n234), .A2(new_n238), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n256), .A2(KEYINPUT30), .A3(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n224), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n257), .B1(new_n203), .B2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT30), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n258), .A2(new_n233), .A3(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n233), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n256), .A2(new_n264), .A3(new_n257), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n265), .A2(new_n266), .A3(new_n247), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n249), .A2(new_n263), .A3(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT31), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n249), .A2(new_n263), .A3(new_n267), .A4(KEYINPUT31), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n256), .A2(new_n273), .A3(new_n257), .ZN(new_n274));
  OAI21_X1  g088(.A(KEYINPUT71), .B1(new_n228), .B2(new_n239), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n274), .A2(new_n275), .A3(new_n264), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT28), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n260), .A2(new_n233), .ZN(new_n279));
  OAI21_X1  g093(.A(KEYINPUT28), .B1(new_n240), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n248), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n272), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT72), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n272), .A2(KEYINPUT72), .A3(new_n282), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NOR2_X1   g101(.A1(G472), .A2(G902), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n188), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  AND3_X1   g103(.A1(new_n272), .A2(KEYINPUT72), .A3(new_n282), .ZN(new_n290));
  AOI21_X1  g104(.A(KEYINPUT72), .B1(new_n272), .B2(new_n282), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n188), .B(new_n288), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n187), .B1(new_n289), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n288), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n295), .B1(new_n285), .B2(new_n286), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(KEYINPUT32), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n263), .A2(new_n265), .ZN(new_n298));
  OR2_X1    g112(.A1(new_n298), .A2(new_n247), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n281), .A2(new_n248), .ZN(new_n301));
  NOR3_X1   g115(.A1(new_n300), .A2(KEYINPUT29), .A3(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT74), .B(G902), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n264), .B1(new_n256), .B2(new_n257), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n305), .A2(new_n240), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n278), .B1(new_n306), .B2(new_n277), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n247), .A2(KEYINPUT29), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n304), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(G472), .B1(new_n302), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n294), .A2(new_n297), .A3(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G221), .ZN(new_n312));
  XOR2_X1   g126(.A(KEYINPUT9), .B(G234), .Z(new_n313));
  INV_X1    g127(.A(G902), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G104), .ZN(new_n316));
  NOR3_X1   g130(.A1(new_n316), .A2(KEYINPUT84), .A3(G107), .ZN(new_n317));
  OAI21_X1  g131(.A(KEYINPUT3), .B1(new_n317), .B2(KEYINPUT83), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT84), .ZN(new_n319));
  INV_X1    g133(.A(G107), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(new_n320), .A3(G104), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT83), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT3), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n318), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G101), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n316), .A2(G107), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(KEYINPUT83), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n320), .A2(G104), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n325), .A2(new_n326), .A3(new_n328), .A4(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT86), .ZN(new_n332));
  OAI21_X1  g146(.A(G101), .B1(new_n327), .B2(new_n329), .ZN(new_n333));
  AND3_X1   g147(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n332), .B1(new_n331), .B2(new_n333), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n259), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NOR3_X1   g150(.A1(new_n317), .A2(KEYINPUT83), .A3(KEYINPUT3), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n323), .B1(new_n321), .B2(new_n322), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n328), .B(new_n330), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n333), .B1(new_n339), .B2(G101), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n208), .B1(new_n215), .B2(new_n209), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n220), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n336), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(KEYINPUT12), .B1(new_n345), .B2(new_n234), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT12), .ZN(new_n347));
  INV_X1    g161(.A(new_n234), .ZN(new_n348));
  AOI211_X1 g162(.A(new_n347), .B(new_n348), .C1(new_n336), .C2(new_n344), .ZN(new_n349));
  OAI21_X1  g163(.A(KEYINPUT88), .B1(new_n346), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n340), .A2(KEYINPUT86), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n224), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n340), .B1(new_n220), .B2(new_n342), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n234), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n347), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT88), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n345), .A2(KEYINPUT12), .A3(new_n234), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n356), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n339), .A2(KEYINPUT85), .A3(KEYINPUT4), .A4(G101), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n331), .A2(KEYINPUT4), .ZN(new_n361));
  AND3_X1   g175(.A1(new_n339), .A2(KEYINPUT85), .A3(G101), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n364));
  AOI22_X1  g178(.A1(new_n363), .A2(new_n238), .B1(new_n344), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT87), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n366), .B1(new_n334), .B2(new_n335), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n351), .A2(KEYINPUT87), .A3(new_n352), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n364), .B1(new_n226), .B2(new_n227), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n365), .A2(new_n370), .A3(new_n348), .ZN(new_n371));
  XNOR2_X1  g185(.A(G110), .B(G140), .ZN(new_n372));
  INV_X1    g186(.A(G227), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n373), .A2(G953), .ZN(new_n374));
  XOR2_X1   g188(.A(new_n372), .B(new_n374), .Z(new_n375));
  NAND4_X1  g189(.A1(new_n350), .A2(new_n359), .A3(new_n371), .A4(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n375), .ZN(new_n377));
  INV_X1    g191(.A(new_n371), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n348), .B1(new_n365), .B2(new_n370), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(G469), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(new_n382), .A3(new_n304), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT89), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n303), .B1(new_n376), .B2(new_n380), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(KEYINPUT89), .A3(new_n382), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n378), .B1(new_n358), .B2(new_n356), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n371), .A2(new_n375), .ZN(new_n390));
  OAI22_X1  g204(.A1(new_n389), .A2(new_n375), .B1(new_n390), .B2(new_n379), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n314), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G469), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n315), .B1(new_n388), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(G214), .B1(G237), .B2(G902), .ZN(new_n395));
  XOR2_X1   g209(.A(new_n395), .B(KEYINPUT90), .Z(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  AND2_X1   g211(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(KEYINPUT77), .B1(new_n209), .B2(G119), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT76), .ZN(new_n400));
  OAI21_X1  g214(.A(KEYINPUT23), .B1(new_n209), .B2(G119), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n399), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n209), .A2(KEYINPUT77), .A3(G119), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n402), .B(new_n403), .C1(new_n400), .C2(new_n401), .ZN(new_n404));
  XNOR2_X1  g218(.A(KEYINPUT65), .B(G128), .ZN(new_n405));
  INV_X1    g219(.A(G119), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT23), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n409), .A2(G110), .ZN(new_n410));
  INV_X1    g224(.A(G125), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n411), .A2(G140), .ZN(new_n412));
  XNOR2_X1  g226(.A(G125), .B(G140), .ZN(new_n413));
  MUX2_X1   g227(.A(new_n412), .B(new_n413), .S(KEYINPUT16), .Z(new_n414));
  XNOR2_X1  g228(.A(new_n414), .B(G146), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n213), .A2(G119), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n416), .B1(G119), .B2(new_n209), .ZN(new_n417));
  XNOR2_X1  g231(.A(KEYINPUT24), .B(G110), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NOR3_X1   g233(.A1(new_n410), .A2(new_n415), .A3(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  OR2_X1    g235(.A1(new_n414), .A2(new_n204), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT78), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n413), .B(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n204), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  OR2_X1    g240(.A1(new_n409), .A2(G110), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n417), .A2(new_n418), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n243), .A2(G221), .A3(G234), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n431), .B(KEYINPUT79), .ZN(new_n432));
  XOR2_X1   g246(.A(new_n432), .B(KEYINPUT22), .Z(new_n433));
  XNOR2_X1  g247(.A(new_n433), .B(new_n189), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n421), .A2(new_n430), .A3(new_n434), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n433), .B(G137), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n436), .B1(new_n420), .B2(new_n429), .ZN(new_n437));
  AND2_X1   g251(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(G234), .ZN(new_n439));
  OAI21_X1  g253(.A(G217), .B1(new_n303), .B2(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n440), .B(KEYINPUT75), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n441), .A2(G902), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n442), .B(KEYINPUT81), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n438), .A2(new_n443), .ZN(new_n444));
  XOR2_X1   g258(.A(new_n444), .B(KEYINPUT82), .Z(new_n445));
  NAND3_X1  g259(.A1(new_n435), .A2(new_n437), .A3(new_n304), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT25), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT25), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n435), .A2(new_n437), .A3(new_n448), .A4(new_n304), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n447), .A2(new_n441), .A3(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT80), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n447), .A2(KEYINPUT80), .A3(new_n441), .A4(new_n449), .ZN(new_n453));
  AND3_X1   g267(.A1(new_n445), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(G113), .B(G122), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(new_n316), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT19), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n413), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n458), .B1(new_n424), .B2(new_n457), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n204), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n422), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(KEYINPUT96), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT95), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n242), .A2(new_n243), .A3(G214), .ZN(new_n464));
  NOR2_X1   g278(.A1(KEYINPUT93), .A2(G143), .ZN(new_n465));
  XOR2_X1   g279(.A(new_n464), .B(new_n465), .Z(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n463), .B1(new_n467), .B2(G131), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(G131), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n466), .A2(KEYINPUT95), .A3(new_n201), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT96), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n460), .A2(new_n472), .A3(new_n422), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n462), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT18), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n466), .B1(new_n475), .B2(new_n201), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT94), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n476), .B(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n467), .A2(KEYINPUT18), .A3(G131), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n425), .B1(new_n204), .B2(new_n413), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n456), .B1(new_n474), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n467), .A2(KEYINPUT17), .A3(G131), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n415), .B(new_n483), .C1(new_n471), .C2(KEYINPUT17), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n484), .A2(new_n481), .A3(new_n456), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(G475), .A2(G902), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n488), .B(KEYINPUT97), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n487), .A2(KEYINPUT20), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n456), .B1(new_n484), .B2(new_n481), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n314), .B1(new_n485), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(G475), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT20), .ZN(new_n494));
  INV_X1    g308(.A(new_n489), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n494), .B1(new_n486), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n490), .A2(new_n493), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT13), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n498), .A2(new_n206), .A3(G128), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n206), .A2(G128), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n500), .B1(new_n405), .B2(new_n206), .ZN(new_n501));
  OAI211_X1 g315(.A(G134), .B(new_n499), .C1(new_n501), .C2(new_n498), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n502), .B1(G134), .B2(new_n501), .ZN(new_n503));
  XNOR2_X1  g317(.A(G116), .B(G122), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n504), .B(G107), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n501), .B(new_n191), .ZN(new_n506));
  INV_X1    g320(.A(G122), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(G116), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n320), .B1(new_n508), .B2(KEYINPUT14), .ZN(new_n509));
  XOR2_X1   g323(.A(new_n509), .B(new_n504), .Z(new_n510));
  OAI22_X1  g324(.A1(new_n503), .A2(new_n505), .B1(new_n506), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n313), .A2(G217), .A3(new_n243), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n511), .B(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n304), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT15), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(G478), .ZN(new_n516));
  XOR2_X1   g330(.A(new_n514), .B(new_n516), .Z(new_n517));
  NOR2_X1   g331(.A1(new_n497), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT98), .B(G952), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n519), .A2(G953), .ZN(new_n520));
  NAND2_X1  g334(.A1(G234), .A2(G237), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  XOR2_X1   g336(.A(KEYINPUT21), .B(G898), .Z(new_n523));
  NAND3_X1  g337(.A1(new_n303), .A2(G953), .A3(new_n521), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n518), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n229), .A2(new_n230), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT5), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n229), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(G113), .ZN(new_n531));
  AND2_X1   g345(.A1(new_n406), .A2(G116), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n531), .B1(new_n532), .B2(new_n528), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n527), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n367), .A2(new_n368), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n363), .A2(new_n233), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  XOR2_X1   g351(.A(G110), .B(G122), .Z(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n538), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n535), .A2(new_n540), .A3(new_n536), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n539), .A2(KEYINPUT6), .A3(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT6), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n537), .A2(new_n543), .A3(new_n538), .ZN(new_n544));
  OR2_X1    g358(.A1(new_n238), .A2(new_n411), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n545), .B1(G125), .B2(new_n224), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n243), .A2(G224), .ZN(new_n547));
  XOR2_X1   g361(.A(new_n546), .B(new_n547), .Z(new_n548));
  NAND3_X1  g362(.A1(new_n542), .A2(new_n544), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n351), .A2(new_n352), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n533), .B(KEYINPUT91), .ZN(new_n551));
  OAI22_X1  g365(.A1(new_n551), .A2(new_n529), .B1(new_n229), .B2(new_n230), .ZN(new_n552));
  OAI22_X1  g366(.A1(new_n550), .A2(new_n552), .B1(new_n341), .B2(new_n534), .ZN(new_n553));
  XOR2_X1   g367(.A(new_n538), .B(KEYINPUT8), .Z(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI22_X1  g369(.A1(new_n545), .A2(KEYINPUT92), .B1(KEYINPUT7), .B2(new_n547), .ZN(new_n556));
  XOR2_X1   g370(.A(new_n556), .B(new_n546), .Z(new_n557));
  NAND3_X1  g371(.A1(new_n541), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n558), .A2(new_n314), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n549), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(G210), .B1(G237), .B2(G902), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n549), .A2(new_n559), .A3(new_n561), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n526), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n311), .A2(new_n398), .A3(new_n454), .A4(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(G101), .ZN(G3));
  NAND2_X1  g383(.A1(new_n287), .A2(new_n288), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(KEYINPUT73), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n304), .B1(new_n290), .B2(new_n291), .ZN(new_n572));
  AOI22_X1  g386(.A1(new_n571), .A2(new_n292), .B1(G472), .B2(new_n572), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n573), .A2(new_n454), .A3(new_n394), .ZN(new_n574));
  XOR2_X1   g388(.A(new_n574), .B(KEYINPUT99), .Z(new_n575));
  AOI21_X1  g389(.A(new_n561), .B1(new_n549), .B2(new_n559), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT100), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n576), .B1(new_n577), .B2(new_n564), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n560), .A2(new_n577), .A3(new_n562), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n397), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n525), .ZN(new_n582));
  OR2_X1    g396(.A1(new_n514), .A2(G478), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n513), .B(KEYINPUT33), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n304), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n584), .B1(G478), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n497), .A2(new_n587), .ZN(new_n588));
  NOR3_X1   g402(.A1(new_n581), .A2(new_n582), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n575), .A2(new_n589), .ZN(new_n590));
  XOR2_X1   g404(.A(KEYINPUT34), .B(G104), .Z(new_n591));
  XNOR2_X1  g405(.A(new_n590), .B(new_n591), .ZN(G6));
  INV_X1    g406(.A(new_n497), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n517), .ZN(new_n594));
  NOR3_X1   g408(.A1(new_n581), .A2(new_n582), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n575), .A2(new_n595), .ZN(new_n596));
  XOR2_X1   g410(.A(KEYINPUT35), .B(G107), .Z(new_n597));
  XNOR2_X1  g411(.A(new_n596), .B(new_n597), .ZN(G9));
  NAND2_X1  g412(.A1(new_n421), .A2(new_n430), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n436), .A2(KEYINPUT36), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n599), .B(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n443), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n452), .A2(new_n453), .A3(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n398), .A2(new_n567), .A3(new_n573), .A4(new_n604), .ZN(new_n605));
  XOR2_X1   g419(.A(new_n605), .B(KEYINPUT37), .Z(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(G110), .ZN(G12));
  NOR2_X1   g421(.A1(new_n581), .A2(new_n594), .ZN(new_n608));
  AND3_X1   g422(.A1(new_n386), .A2(KEYINPUT89), .A3(new_n382), .ZN(new_n609));
  AOI21_X1  g423(.A(KEYINPUT89), .B1(new_n386), .B2(new_n382), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n393), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n315), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n522), .B1(G900), .B2(new_n524), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n311), .A2(new_n608), .A3(new_n604), .A4(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(G128), .ZN(G30));
  XNOR2_X1  g431(.A(new_n565), .B(KEYINPUT38), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(new_n613), .B(KEYINPUT39), .Z(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n394), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n619), .B1(new_n622), .B2(KEYINPUT40), .ZN(new_n623));
  INV_X1    g437(.A(new_n268), .ZN(new_n624));
  INV_X1    g438(.A(new_n306), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n624), .B1(new_n248), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(G472), .B1(new_n626), .B2(G902), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n294), .A2(new_n297), .A3(new_n627), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n623), .A2(new_n603), .A3(new_n628), .ZN(new_n629));
  OR2_X1    g443(.A1(new_n622), .A2(KEYINPUT40), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n497), .A2(new_n517), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n629), .A2(new_n397), .A3(new_n630), .A4(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G143), .ZN(G45));
  NOR2_X1   g447(.A1(new_n581), .A2(new_n588), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n311), .A2(new_n634), .A3(new_n604), .A4(new_n615), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G146), .ZN(G48));
  AND2_X1   g450(.A1(new_n311), .A2(new_n454), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n386), .A2(new_n382), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n639), .B(new_n612), .C1(new_n609), .C2(new_n610), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(KEYINPUT101), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n637), .A2(new_n589), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(KEYINPUT41), .B(G113), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G15));
  AND2_X1   g458(.A1(new_n637), .A2(new_n641), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n595), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT102), .B(G116), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G18));
  INV_X1    g462(.A(new_n526), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n640), .A2(new_n581), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n311), .A2(new_n649), .A3(new_n604), .A4(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT103), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(new_n406), .ZN(G21));
  NAND2_X1  g467(.A1(new_n564), .A2(new_n577), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n563), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n396), .B1(new_n655), .B2(new_n579), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n631), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT104), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n307), .A2(new_n659), .ZN(new_n660));
  OAI211_X1 g474(.A(new_n278), .B(KEYINPUT104), .C1(new_n306), .C2(new_n277), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n660), .A2(new_n248), .A3(new_n661), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n295), .B1(new_n662), .B2(new_n272), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n663), .B1(new_n572), .B2(G472), .ZN(new_n664));
  AND3_X1   g478(.A1(new_n664), .A2(new_n454), .A3(new_n525), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n641), .A2(new_n658), .A3(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT105), .ZN(new_n667));
  OR2_X1    g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n666), .A2(new_n667), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G122), .ZN(G24));
  INV_X1    g485(.A(KEYINPUT106), .ZN(new_n672));
  INV_X1    g486(.A(new_n613), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n588), .A2(new_n673), .ZN(new_n674));
  AOI211_X1 g488(.A(new_n663), .B(new_n603), .C1(new_n572), .C2(G472), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n650), .A2(new_n672), .A3(new_n674), .A4(new_n675), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n638), .B1(new_n385), .B2(new_n387), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n656), .A2(new_n677), .A3(new_n612), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n572), .A2(G472), .ZN(new_n679));
  INV_X1    g493(.A(new_n663), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n679), .A2(new_n604), .A3(new_n680), .A4(new_n674), .ZN(new_n681));
  OAI21_X1  g495(.A(KEYINPUT106), .B1(new_n678), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n676), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G125), .ZN(G27));
  NOR2_X1   g498(.A1(new_n296), .A2(KEYINPUT32), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(KEYINPUT108), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT108), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n687), .B1(new_n296), .B2(KEYINPUT32), .ZN(new_n688));
  OAI211_X1 g502(.A(new_n686), .B(new_n310), .C1(new_n688), .C2(new_n685), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT107), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n566), .A2(new_n690), .A3(new_n397), .ZN(new_n691));
  OAI21_X1  g505(.A(KEYINPUT107), .B1(new_n565), .B2(new_n396), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n394), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n689), .A2(new_n693), .A3(new_n454), .A4(new_n674), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(KEYINPUT42), .ZN(new_n695));
  INV_X1    g509(.A(new_n674), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n696), .A2(KEYINPUT42), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n311), .A2(new_n693), .A3(new_n454), .A4(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(new_n201), .ZN(G33));
  INV_X1    g514(.A(new_n594), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n311), .A2(new_n693), .A3(new_n454), .A4(new_n701), .ZN(new_n702));
  OR2_X1    g516(.A1(new_n702), .A2(new_n673), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G134), .ZN(G36));
  NAND2_X1  g518(.A1(new_n691), .A2(new_n692), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n593), .A2(new_n587), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(KEYINPUT43), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n573), .A2(new_n603), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n705), .B1(new_n708), .B2(KEYINPUT44), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n391), .B(KEYINPUT45), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(G469), .ZN(new_n711));
  NAND2_X1  g525(.A1(G469), .A2(G902), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n711), .A2(KEYINPUT46), .A3(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT46), .ZN(new_n714));
  OAI211_X1 g528(.A(new_n714), .B(G469), .C1(new_n710), .C2(G902), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n713), .A2(new_n388), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n612), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n717), .A2(new_n620), .ZN(new_n718));
  OAI211_X1 g532(.A(new_n709), .B(new_n718), .C1(KEYINPUT44), .C2(new_n708), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G137), .ZN(G39));
  NOR4_X1   g534(.A1(new_n311), .A2(new_n705), .A3(new_n454), .A4(new_n696), .ZN(new_n721));
  XOR2_X1   g535(.A(new_n721), .B(KEYINPUT109), .Z(new_n722));
  XOR2_X1   g536(.A(new_n717), .B(KEYINPUT47), .Z(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G140), .ZN(G42));
  AND2_X1   g539(.A1(new_n642), .A2(new_n651), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n568), .A2(new_n605), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n573), .A2(new_n454), .A3(new_n394), .A4(new_n525), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n594), .A2(new_n588), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n730), .A2(new_n566), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n728), .A2(new_n396), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g547(.A(KEYINPUT111), .B1(new_n727), .B2(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n574), .A2(new_n397), .A3(new_n525), .A4(new_n731), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT111), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n735), .A2(new_n736), .A3(new_n568), .A4(new_n605), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  AOI22_X1  g552(.A1(new_n669), .A2(new_n668), .B1(new_n645), .B2(new_n595), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n693), .A2(KEYINPUT112), .A3(new_n674), .A4(new_n675), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT112), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n394), .A2(new_n691), .A3(new_n692), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n741), .B1(new_n742), .B2(new_n681), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n695), .A2(new_n744), .A3(new_n698), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n311), .A2(new_n518), .A3(new_n604), .A4(new_n615), .ZN(new_n746));
  OAI22_X1  g560(.A1(new_n702), .A2(new_n673), .B1(new_n746), .B2(new_n705), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  AND4_X1   g562(.A1(new_n726), .A2(new_n738), .A3(new_n739), .A4(new_n748), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n614), .A2(new_n657), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n628), .A2(new_n750), .A3(new_n603), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n616), .A2(new_n635), .A3(new_n683), .A4(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n749), .A2(KEYINPUT53), .A3(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n738), .A2(new_n739), .A3(new_n748), .A4(new_n726), .ZN(new_n756));
  OR2_X1    g570(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n752), .A2(new_n753), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n752), .A2(new_n753), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  XOR2_X1   g574(.A(KEYINPUT113), .B(KEYINPUT114), .Z(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n754), .A2(new_n761), .A3(new_n757), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n756), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n755), .B1(new_n765), .B2(KEYINPUT53), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(KEYINPUT54), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT53), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n749), .A2(new_n768), .A3(new_n754), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n769), .B1(new_n765), .B2(new_n768), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT54), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n707), .A2(new_n522), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n773), .A2(new_n454), .A3(new_n664), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n774), .A2(new_n640), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n656), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(new_n396), .A3(new_n619), .ZN(new_n777));
  XOR2_X1   g591(.A(KEYINPUT116), .B(KEYINPUT50), .Z(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n628), .ZN(new_n780));
  INV_X1    g594(.A(new_n522), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n705), .A2(new_n640), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n780), .A2(new_n454), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  OR3_X1    g597(.A1(new_n783), .A2(new_n497), .A3(new_n587), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n782), .A2(new_n773), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n675), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n779), .A2(new_n784), .A3(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  OR3_X1    g603(.A1(new_n777), .A2(KEYINPUT116), .A3(KEYINPUT50), .ZN(new_n790));
  OR3_X1    g604(.A1(new_n774), .A2(KEYINPUT115), .A3(new_n705), .ZN(new_n791));
  OAI21_X1  g605(.A(KEYINPUT115), .B1(new_n774), .B2(new_n705), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n677), .B(KEYINPUT110), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n612), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n791), .B(new_n792), .C1(new_n723), .C2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n789), .A2(new_n790), .A3(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT51), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n789), .A2(new_n790), .A3(KEYINPUT51), .A4(new_n795), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n689), .A2(new_n454), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n786), .A2(new_n800), .ZN(new_n801));
  XOR2_X1   g615(.A(new_n801), .B(KEYINPUT48), .Z(new_n802));
  OAI21_X1  g616(.A(new_n520), .B1(new_n783), .B2(new_n588), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n798), .A2(new_n799), .A3(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n767), .A2(new_n772), .A3(new_n776), .A4(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(G952), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(new_n243), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  XOR2_X1   g623(.A(new_n793), .B(KEYINPUT49), .Z(new_n810));
  NOR3_X1   g624(.A1(new_n618), .A2(new_n396), .A3(new_n706), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n780), .A2(new_n454), .A3(new_n612), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n809), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT117), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n809), .A2(KEYINPUT117), .A3(new_n813), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(G75));
  NAND2_X1  g632(.A1(new_n807), .A2(G953), .ZN(new_n819));
  XOR2_X1   g633(.A(new_n819), .B(KEYINPUT119), .Z(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n770), .A2(new_n304), .A3(new_n561), .ZN(new_n822));
  OR2_X1    g636(.A1(new_n822), .A2(KEYINPUT56), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n542), .A2(new_n544), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(new_n548), .ZN(new_n825));
  XOR2_X1   g639(.A(KEYINPUT118), .B(KEYINPUT55), .Z(new_n826));
  XNOR2_X1  g640(.A(new_n825), .B(new_n826), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n823), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n823), .A2(new_n827), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n821), .B1(new_n828), .B2(new_n829), .ZN(G51));
  OR2_X1    g644(.A1(new_n765), .A2(new_n768), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT121), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n831), .A2(new_n832), .A3(KEYINPUT54), .A4(new_n769), .ZN(new_n833));
  OAI21_X1  g647(.A(KEYINPUT121), .B1(new_n770), .B2(new_n771), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n833), .A2(new_n772), .A3(new_n834), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n712), .B(KEYINPUT120), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(KEYINPUT57), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(new_n381), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n770), .A2(new_n304), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n840), .A2(G469), .A3(new_n710), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n821), .B1(new_n839), .B2(new_n841), .ZN(G54));
  NAND3_X1  g656(.A1(new_n840), .A2(KEYINPUT58), .A3(G475), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n843), .A2(KEYINPUT122), .A3(new_n486), .ZN(new_n844));
  AOI21_X1  g658(.A(KEYINPUT122), .B1(new_n843), .B2(new_n486), .ZN(new_n845));
  AND4_X1   g659(.A1(KEYINPUT58), .A2(new_n840), .A3(G475), .A4(new_n487), .ZN(new_n846));
  NOR4_X1   g660(.A1(new_n844), .A2(new_n845), .A3(new_n821), .A4(new_n846), .ZN(G60));
  NAND2_X1  g661(.A1(G478), .A2(G902), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n848), .B(KEYINPUT59), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n835), .A2(new_n585), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n767), .A2(new_n772), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n585), .B1(new_n851), .B2(new_n849), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n850), .A2(new_n821), .A3(new_n852), .ZN(G63));
  NAND2_X1  g667(.A1(G217), .A2(G902), .ZN(new_n854));
  XOR2_X1   g668(.A(new_n854), .B(KEYINPUT123), .Z(new_n855));
  XNOR2_X1  g669(.A(new_n855), .B(KEYINPUT60), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n770), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(new_n601), .ZN(new_n858));
  OR2_X1    g672(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n859));
  INV_X1    g673(.A(new_n438), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n860), .B1(new_n770), .B2(new_n856), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n858), .A2(new_n820), .A3(new_n859), .A4(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n862), .B(new_n863), .ZN(G66));
  AOI21_X1  g678(.A(new_n243), .B1(new_n523), .B2(G224), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n738), .A2(new_n739), .A3(new_n726), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n865), .B1(new_n866), .B2(new_n243), .ZN(new_n867));
  INV_X1    g681(.A(G898), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n824), .B1(new_n868), .B2(G953), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n867), .B(new_n869), .ZN(G69));
  NAND2_X1  g684(.A1(new_n258), .A2(new_n262), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(new_n459), .Z(new_n872));
  NAND2_X1  g686(.A1(new_n373), .A2(G953), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n724), .A2(new_n719), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n616), .A2(new_n635), .A3(new_n683), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n718), .A2(new_n800), .A3(new_n658), .ZN(new_n876));
  AND4_X1   g690(.A1(new_n695), .A2(new_n875), .A3(new_n876), .A4(new_n698), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n874), .A2(new_n703), .A3(new_n877), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n872), .B(new_n873), .C1(new_n878), .C2(G953), .ZN(new_n879));
  OAI21_X1  g693(.A(G900), .B1(new_n872), .B2(G227), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(G953), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n622), .A2(new_n705), .A3(new_n730), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n637), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n632), .A2(new_n875), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT62), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n884), .B(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n874), .A2(new_n883), .A3(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  OR2_X1    g702(.A1(new_n872), .A2(G953), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n879), .B(new_n881), .C1(new_n888), .C2(new_n889), .ZN(G72));
  NAND2_X1  g704(.A1(G472), .A2(G902), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n891), .B(KEYINPUT63), .Z(new_n892));
  OAI211_X1 g706(.A(new_n766), .B(new_n892), .C1(new_n624), .C2(new_n300), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT127), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n892), .B1(new_n887), .B2(new_n866), .ZN(new_n895));
  OR2_X1    g709(.A1(new_n895), .A2(KEYINPUT125), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n298), .B1(new_n895), .B2(KEYINPUT125), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n896), .A2(new_n247), .A3(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(new_n892), .ZN(new_n899));
  INV_X1    g713(.A(new_n866), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n899), .B1(new_n878), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n298), .A2(new_n248), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT126), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n820), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n894), .A2(new_n898), .A3(new_n904), .ZN(G57));
endmodule


