//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 0 1 1 1 1 1 0 1 1 0 0 1 1 1 1 1 0 1 1 1 1 1 1 0 0 0 1 0 0 0 0 0 1 1 1 0 1 1 0 1 0 1 0 0 1 0 1 0 0 1 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:18 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1268, new_n1269, new_n1270, new_n1271, new_n1273,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1353,
    new_n1354;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  XNOR2_X1  g0001(.A(new_n201), .B(KEYINPUT64), .ZN(new_n202));
  INV_X1    g0002(.A(G77), .ZN(new_n203));
  AND2_X1   g0003(.A1(new_n202), .A2(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  OAI21_X1  g0005(.A(G50), .B1(G58), .B2(G68), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G1), .A2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NAND3_X1  g0009(.A1(new_n207), .A2(G20), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  XOR2_X1   g0014(.A(KEYINPUT65), .B(G77), .Z(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(KEYINPUT66), .B(G244), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G107), .A2(G264), .ZN(new_n222));
  NAND4_X1  g0022(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n211), .B1(new_n218), .B2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n210), .B(new_n214), .C1(new_n224), .C2(KEYINPUT1), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G250), .B(G257), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT67), .ZN(new_n228));
  XOR2_X1   g0028(.A(G264), .B(G270), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n230), .B(new_n235), .ZN(G358));
  XNOR2_X1  g0036(.A(G68), .B(G77), .ZN(new_n237));
  INV_X1    g0037(.A(G58), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT68), .B(G50), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G351));
  INV_X1    g0045(.A(G1), .ZN(new_n246));
  NAND3_X1  g0046(.A1(new_n246), .A2(G13), .A3(G20), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G97), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n208), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n246), .A2(G33), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n253), .A2(new_n247), .A3(new_n254), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n250), .B1(new_n255), .B2(new_n249), .ZN(new_n256));
  INV_X1    g0056(.A(G107), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(KEYINPUT6), .A3(G97), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT82), .ZN(new_n259));
  OR2_X1    g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT6), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n249), .A2(new_n257), .ZN(new_n262));
  NOR2_X1   g0062(.A1(G97), .A2(G107), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n261), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n258), .A2(new_n259), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n260), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(G20), .A2(G33), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n266), .A2(G20), .B1(G77), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G20), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT77), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT3), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n273));
  AOI21_X1  g0073(.A(G33), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G33), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n275), .A2(KEYINPUT3), .ZN(new_n276));
  OAI211_X1 g0076(.A(KEYINPUT7), .B(new_n269), .C1(new_n274), .C2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT7), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n271), .A2(G33), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(new_n276), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n278), .B1(new_n280), .B2(G20), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n277), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n268), .B1(new_n282), .B2(new_n257), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n256), .B1(new_n283), .B2(new_n252), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT5), .B(G41), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n246), .A2(G45), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(G33), .A2(G41), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n289), .A2(G1), .A3(G13), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n288), .A2(G257), .A3(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G274), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n292), .B1(new_n209), .B2(new_n289), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n293), .A2(new_n287), .A3(new_n285), .ZN(new_n294));
  AND2_X1   g0094(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n275), .A2(KEYINPUT3), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n271), .A2(G33), .ZN(new_n297));
  AND2_X1   g0097(.A1(KEYINPUT4), .A2(G244), .ZN(new_n298));
  INV_X1    g0098(.A(G1698), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n296), .A2(new_n297), .A3(new_n298), .A4(new_n299), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n296), .A2(new_n297), .A3(G250), .A4(G1698), .ZN(new_n301));
  NAND2_X1  g0101(.A1(G33), .A2(G283), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT4), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n272), .A2(G33), .A3(new_n273), .ZN(new_n305));
  INV_X1    g0105(.A(G244), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n306), .A2(G1698), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n305), .A2(new_n296), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n303), .B1(new_n304), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n295), .B1(new_n309), .B2(new_n290), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n310), .A2(G179), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n291), .A2(new_n294), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n308), .A2(new_n304), .ZN(new_n313));
  AND3_X1   g0113(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n290), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n312), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n317), .A2(G169), .ZN(new_n318));
  NOR3_X1   g0118(.A1(new_n284), .A2(new_n311), .A3(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT83), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n310), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n317), .A2(KEYINPUT83), .ZN(new_n322));
  AND3_X1   g0122(.A1(new_n321), .A2(new_n322), .A3(G200), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n317), .A2(G190), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n284), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g0125(.A(KEYINPUT84), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n268), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n257), .B1(new_n277), .B2(new_n281), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n252), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n256), .ZN(new_n330));
  AND3_X1   g0130(.A1(new_n329), .A2(new_n324), .A3(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT84), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n321), .A2(new_n322), .A3(G200), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n319), .B1(new_n326), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT14), .ZN(new_n336));
  XOR2_X1   g0136(.A(KEYINPUT75), .B(KEYINPUT13), .Z(new_n337));
  INV_X1    g0137(.A(G41), .ZN(new_n338));
  INV_X1    g0138(.A(G45), .ZN(new_n339));
  AOI21_X1  g0139(.A(G1), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(KEYINPUT69), .B1(new_n293), .B2(new_n340), .ZN(new_n341));
  AND4_X1   g0141(.A1(KEYINPUT69), .A2(new_n340), .A3(new_n290), .A4(G274), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT73), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n246), .B1(G41), .B2(G45), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n290), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(G238), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n343), .B1(new_n290), .B2(new_n344), .ZN(new_n347));
  OAI22_X1  g0147(.A1(new_n341), .A2(new_n342), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT74), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n340), .A2(new_n290), .A3(G274), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT69), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n293), .A2(KEYINPUT69), .A3(new_n340), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n290), .A2(new_n344), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(KEYINPUT73), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n357), .A2(G238), .A3(new_n345), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n355), .A2(new_n358), .A3(KEYINPUT74), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n350), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n296), .A2(new_n297), .A3(G232), .A4(G1698), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n296), .A2(new_n297), .A3(G226), .A4(new_n299), .ZN(new_n362));
  NAND2_X1  g0162(.A1(G33), .A2(G97), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(new_n316), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n337), .B1(new_n360), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n337), .ZN(new_n367));
  INV_X1    g0167(.A(new_n365), .ZN(new_n368));
  AOI211_X1 g0168(.A(new_n367), .B(new_n368), .C1(new_n350), .C2(new_n359), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n336), .B(G169), .C1(new_n366), .C2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(KEYINPUT76), .ZN(new_n371));
  OAI21_X1  g0171(.A(G169), .B1(new_n366), .B2(new_n369), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(KEYINPUT14), .ZN(new_n373));
  AND3_X1   g0173(.A1(new_n355), .A2(new_n358), .A3(KEYINPUT74), .ZN(new_n374));
  AOI21_X1  g0174(.A(KEYINPUT74), .B1(new_n355), .B2(new_n358), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n365), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n367), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n360), .A2(new_n337), .A3(new_n365), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT76), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n379), .A2(new_n380), .A3(new_n336), .A4(G169), .ZN(new_n381));
  INV_X1    g0181(.A(new_n376), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT13), .ZN(new_n383));
  OAI211_X1 g0183(.A(G179), .B(new_n378), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n371), .A2(new_n373), .A3(new_n381), .A4(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(G68), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n248), .A2(new_n386), .ZN(new_n387));
  XNOR2_X1  g0187(.A(new_n387), .B(KEYINPUT12), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n267), .A2(G50), .B1(G20), .B2(new_n386), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n269), .A2(G33), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n389), .B1(new_n203), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n391), .A2(KEYINPUT11), .A3(new_n252), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n248), .A2(new_n252), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n393), .B(G68), .C1(G1), .C2(new_n269), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n388), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT11), .B1(new_n391), .B2(new_n252), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n385), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n378), .B1(new_n382), .B2(new_n383), .ZN(new_n400));
  INV_X1    g0200(.A(G190), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n397), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(G200), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n403), .B1(new_n377), .B2(new_n378), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n399), .A2(new_n406), .ZN(new_n407));
  XNOR2_X1  g0207(.A(KEYINPUT8), .B(G58), .ZN(new_n408));
  INV_X1    g0208(.A(G150), .ZN(new_n409));
  INV_X1    g0209(.A(new_n267), .ZN(new_n410));
  OAI22_X1  g0210(.A1(new_n408), .A2(new_n390), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OAI22_X1  g0211(.A1(new_n202), .A2(new_n269), .B1(new_n411), .B2(KEYINPUT71), .ZN(new_n412));
  AND2_X1   g0212(.A1(new_n411), .A2(KEYINPUT71), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n252), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(G50), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n415), .B1(new_n246), .B2(G20), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n393), .A2(new_n416), .B1(new_n415), .B2(new_n248), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT9), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g0220(.A(new_n420), .B(KEYINPUT72), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT70), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n280), .A2(new_n299), .ZN(new_n423));
  INV_X1    g0223(.A(G222), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n280), .A2(KEYINPUT70), .A3(G222), .A4(new_n299), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n296), .A2(new_n297), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n428), .A2(new_n299), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n429), .A2(G223), .B1(new_n215), .B2(new_n428), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n290), .B1(new_n427), .B2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(G226), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n355), .B1(new_n432), .B2(new_n356), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(G200), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n434), .A2(G190), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n418), .A2(new_n419), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(KEYINPUT10), .B1(new_n421), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT72), .ZN(new_n441));
  XNOR2_X1  g0241(.A(new_n420), .B(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT10), .ZN(new_n443));
  AND2_X1   g0243(.A1(new_n437), .A2(new_n438), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n442), .A2(new_n443), .A3(new_n436), .A4(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n440), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(G169), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n435), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(G179), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n434), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n448), .A2(new_n418), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n446), .A2(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(G223), .A2(G1698), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n453), .B1(new_n432), .B2(G1698), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n454), .A2(new_n305), .A3(new_n296), .ZN(new_n455));
  NAND2_X1  g0255(.A1(G33), .A2(G87), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(new_n316), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n290), .A2(G232), .A3(new_n344), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT79), .ZN(new_n460));
  XNOR2_X1  g0260(.A(new_n459), .B(new_n460), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n458), .A2(new_n401), .A3(new_n461), .A4(new_n355), .ZN(new_n462));
  AND3_X1   g0262(.A1(new_n458), .A2(new_n355), .A3(new_n461), .ZN(new_n463));
  OAI211_X1 g0263(.A(KEYINPUT81), .B(new_n462), .C1(new_n463), .C2(G200), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT16), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n386), .B1(new_n277), .B2(new_n281), .ZN(new_n466));
  INV_X1    g0266(.A(G159), .ZN(new_n467));
  OAI21_X1  g0267(.A(KEYINPUT78), .B1(new_n410), .B2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT78), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n267), .A2(new_n469), .A3(G159), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  XNOR2_X1  g0271(.A(G58), .B(G68), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(G20), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n465), .B1(new_n466), .B2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n474), .ZN(new_n476));
  AOI21_X1  g0276(.A(G20), .B1(new_n305), .B2(new_n296), .ZN(new_n477));
  OAI21_X1  g0277(.A(G68), .B1(new_n477), .B2(new_n278), .ZN(new_n478));
  AND2_X1   g0278(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n479));
  NOR2_X1   g0279(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n279), .B1(new_n481), .B2(G33), .ZN(new_n482));
  NOR3_X1   g0282(.A1(new_n482), .A2(KEYINPUT7), .A3(G20), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n476), .B1(new_n478), .B2(new_n483), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n475), .B(new_n252), .C1(new_n484), .C2(new_n465), .ZN(new_n485));
  OR2_X1    g0285(.A1(new_n462), .A2(KEYINPUT81), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n408), .B1(new_n246), .B2(G20), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n487), .A2(new_n393), .B1(new_n248), .B2(new_n408), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n464), .A2(new_n485), .A3(new_n486), .A4(new_n488), .ZN(new_n489));
  XNOR2_X1  g0289(.A(new_n489), .B(KEYINPUT17), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n485), .A2(new_n488), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n458), .A2(G179), .A3(new_n461), .A4(new_n355), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n492), .B1(new_n463), .B2(new_n447), .ZN(new_n493));
  AOI21_X1  g0293(.A(KEYINPUT18), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT80), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n491), .A2(KEYINPUT18), .A3(new_n493), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n491), .A2(new_n493), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT18), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n498), .A2(new_n495), .A3(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n490), .B1(new_n497), .B2(new_n501), .ZN(new_n502));
  XNOR2_X1  g0302(.A(KEYINPUT15), .B(G87), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n390), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n504), .A2(new_n505), .B1(new_n215), .B2(G20), .ZN(new_n506));
  INV_X1    g0306(.A(new_n408), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n267), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n253), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n393), .ZN(new_n510));
  OAI21_X1  g0310(.A(G77), .B1(new_n269), .B2(G1), .ZN(new_n511));
  OAI22_X1  g0311(.A1(new_n510), .A2(new_n511), .B1(new_n215), .B2(new_n247), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n355), .B1(new_n217), .B2(new_n356), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n429), .A2(G238), .B1(G107), .B2(new_n428), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(new_n232), .B2(new_n423), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n515), .B1(new_n517), .B2(new_n316), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n514), .B1(new_n518), .B2(G190), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n519), .B1(new_n403), .B2(new_n518), .ZN(new_n520));
  OR2_X1    g0320(.A1(new_n518), .A2(G169), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n518), .A2(new_n449), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n521), .A2(new_n514), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  NOR4_X1   g0324(.A1(new_n407), .A2(new_n452), .A3(new_n502), .A4(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n503), .A2(new_n248), .ZN(new_n526));
  INV_X1    g0326(.A(new_n255), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n504), .ZN(new_n528));
  XOR2_X1   g0328(.A(KEYINPUT85), .B(G87), .Z(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n263), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT19), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n531), .B1(new_n363), .B2(new_n269), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n531), .B1(new_n390), .B2(new_n249), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n482), .A2(new_n269), .A3(G68), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT86), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n482), .A2(KEYINPUT86), .A3(new_n269), .A4(G68), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n535), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n526), .B(new_n528), .C1(new_n540), .C2(new_n253), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n293), .A2(new_n287), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n290), .A2(G250), .A3(new_n286), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(G238), .A2(G1698), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n546), .B1(new_n306), .B2(G1698), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n547), .A2(new_n305), .A3(new_n296), .ZN(new_n548));
  INV_X1    g0348(.A(G116), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n548), .B1(new_n275), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n545), .B1(new_n550), .B2(new_n316), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n447), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n551), .A2(new_n449), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(G87), .ZN(new_n556));
  OAI221_X1 g0356(.A(new_n526), .B1(new_n556), .B2(new_n255), .C1(new_n540), .C2(new_n253), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n552), .A2(G200), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n551), .A2(G190), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI22_X1  g0360(.A1(new_n542), .A2(new_n555), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n290), .A2(G274), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n288), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n316), .B1(new_n287), .B2(new_n285), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n564), .B1(new_n565), .B2(G270), .ZN(new_n566));
  MUX2_X1   g0366(.A(G257), .B(G264), .S(G1698), .Z(new_n567));
  AOI22_X1  g0367(.A1(new_n482), .A2(new_n567), .B1(G303), .B2(new_n428), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n566), .B1(new_n290), .B2(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n302), .B(new_n269), .C1(G33), .C2(new_n249), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT87), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT20), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n571), .A2(new_n572), .B1(new_n549), .B2(G20), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n570), .A2(new_n573), .A3(new_n252), .ZN(new_n574));
  NAND2_X1  g0374(.A1(KEYINPUT87), .A2(KEYINPUT20), .ZN(new_n575));
  XNOR2_X1  g0375(.A(new_n574), .B(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n247), .A2(new_n549), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(new_n527), .B2(new_n549), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n569), .A2(G169), .A3(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT21), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n566), .B(G190), .C1(new_n290), .C2(new_n568), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n576), .A2(new_n578), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n482), .A2(new_n567), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n428), .A2(G303), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n290), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n288), .A2(new_n290), .ZN(new_n588));
  INV_X1    g0388(.A(G270), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n294), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n583), .B(new_n584), .C1(new_n403), .C2(new_n591), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n569), .A2(new_n579), .A3(KEYINPUT21), .A4(G169), .ZN(new_n593));
  NOR3_X1   g0393(.A1(new_n587), .A2(new_n449), .A3(new_n590), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n579), .ZN(new_n595));
  AND4_X1   g0395(.A1(new_n582), .A2(new_n592), .A3(new_n593), .A4(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n248), .A2(KEYINPUT25), .A3(new_n257), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(KEYINPUT90), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT25), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n599), .B1(new_n247), .B2(G107), .ZN(new_n600));
  OR2_X1    g0400(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n598), .A2(new_n600), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n601), .A2(new_n602), .B1(G107), .B2(new_n527), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT22), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n604), .A2(new_n556), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n305), .A2(new_n269), .A3(new_n296), .A4(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n269), .A2(G87), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n604), .B1(new_n428), .B2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT23), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(new_n269), .B2(G107), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n257), .A2(KEYINPUT23), .A3(G20), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n275), .A2(new_n549), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n610), .A2(new_n611), .B1(new_n612), .B2(new_n269), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n606), .A2(new_n608), .A3(new_n613), .ZN(new_n614));
  OR2_X1    g0414(.A1(new_n614), .A2(KEYINPUT89), .ZN(new_n615));
  XOR2_X1   g0415(.A(KEYINPUT88), .B(KEYINPUT24), .Z(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n614), .A2(KEYINPUT89), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n615), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n252), .B1(new_n618), .B2(new_n617), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n603), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  MUX2_X1   g0421(.A(G250), .B(G257), .S(G1698), .Z(new_n622));
  NAND3_X1  g0422(.A1(new_n622), .A2(new_n305), .A3(new_n296), .ZN(new_n623));
  NAND2_X1  g0423(.A1(G33), .A2(G294), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n290), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n288), .A2(G264), .A3(new_n290), .ZN(new_n626));
  NOR3_X1   g0426(.A1(new_n625), .A2(new_n626), .A3(new_n564), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n627), .A2(G169), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n628), .B1(new_n449), .B2(new_n627), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n621), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n627), .A2(new_n401), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n631), .B1(G200), .B2(new_n627), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n632), .B(new_n603), .C1(new_n619), .C2(new_n620), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n596), .A2(new_n630), .A3(new_n633), .ZN(new_n634));
  AND4_X1   g0434(.A1(new_n335), .A2(new_n525), .A3(new_n562), .A4(new_n634), .ZN(G372));
  INV_X1    g0435(.A(new_n555), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n541), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT26), .ZN(new_n639));
  OR3_X1    g0439(.A1(new_n284), .A2(new_n311), .A3(new_n318), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n639), .B1(new_n561), .B2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n557), .ZN(new_n642));
  INV_X1    g0442(.A(new_n560), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n644), .A2(new_n637), .A3(new_n319), .A4(KEYINPUT26), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n638), .B1(new_n641), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n335), .A2(new_n562), .A3(new_n633), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n621), .A2(new_n629), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n582), .A2(new_n593), .A3(new_n595), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT91), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n582), .A2(new_n593), .A3(KEYINPUT91), .A4(new_n595), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n648), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n646), .B1(new_n647), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n525), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n451), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n498), .A2(new_n499), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n496), .ZN(new_n658));
  INV_X1    g0458(.A(new_n523), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n406), .A2(new_n659), .B1(new_n385), .B2(new_n398), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n485), .A2(new_n488), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n661), .A2(KEYINPUT17), .A3(new_n486), .A4(new_n464), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT17), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n489), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n658), .B1(new_n660), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n656), .B1(new_n666), .B2(new_n446), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n655), .A2(new_n667), .ZN(G369));
  NAND3_X1  g0468(.A1(new_n246), .A2(new_n269), .A3(G13), .ZN(new_n669));
  OR2_X1    g0469(.A1(new_n669), .A2(KEYINPUT27), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(KEYINPUT27), .ZN(new_n671));
  AND3_X1   g0471(.A1(new_n670), .A2(G213), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(G343), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n673), .B(KEYINPUT92), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(new_n579), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n596), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n651), .A2(new_n652), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n677), .B1(new_n678), .B2(new_n676), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(G330), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n630), .A2(new_n633), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n621), .A2(new_n675), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n648), .A2(new_n675), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n681), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n649), .A2(new_n674), .ZN(new_n689));
  OAI22_X1  g0489(.A1(new_n682), .A2(new_n689), .B1(new_n630), .B2(new_n675), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n688), .A2(new_n691), .ZN(G399));
  INV_X1    g0492(.A(new_n212), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(G41), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(G1), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n529), .A2(new_n549), .A3(new_n263), .ZN(new_n697));
  OAI22_X1  g0497(.A1(new_n696), .A2(new_n697), .B1(new_n206), .B2(new_n695), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT28), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n654), .A2(new_n674), .ZN(new_n700));
  XNOR2_X1  g0500(.A(KEYINPUT97), .B(KEYINPUT29), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n648), .A2(new_n649), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n703), .A2(new_n335), .A3(new_n562), .A4(new_n633), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n675), .B1(new_n704), .B2(new_n646), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(KEYINPUT29), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n594), .A2(new_n317), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n625), .A2(new_n626), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n551), .A2(new_n708), .A3(KEYINPUT93), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n551), .A2(new_n708), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT93), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n707), .A2(KEYINPUT30), .A3(new_n709), .A4(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n712), .A2(new_n317), .A3(new_n594), .A4(new_n709), .ZN(new_n715));
  XNOR2_X1  g0515(.A(KEYINPUT94), .B(KEYINPUT30), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(KEYINPUT95), .B1(new_n317), .B2(new_n627), .ZN(new_n718));
  INV_X1    g0518(.A(new_n626), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n623), .A2(new_n624), .ZN(new_n720));
  OAI211_X1 g0520(.A(new_n719), .B(new_n294), .C1(new_n720), .C2(new_n290), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT95), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n310), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n718), .A2(new_n723), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n591), .A2(G179), .A3(new_n551), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n717), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n714), .B1(new_n727), .B2(KEYINPUT96), .ZN(new_n728));
  AOI22_X1  g0528(.A1(new_n715), .A2(new_n716), .B1(new_n724), .B2(new_n725), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT96), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n732), .A2(KEYINPUT31), .A3(new_n675), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n717), .A2(new_n713), .A3(new_n726), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(new_n675), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT31), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n634), .A2(new_n335), .A3(new_n562), .A4(new_n674), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n733), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  AOI22_X1  g0539(.A1(new_n702), .A2(new_n706), .B1(G330), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n699), .B1(new_n740), .B2(G1), .ZN(G364));
  AND2_X1   g0541(.A1(new_n269), .A2(G13), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n246), .B1(new_n742), .B2(G45), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(new_n694), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n681), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n746), .B1(G330), .B2(new_n679), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n693), .A2(new_n428), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G355), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n749), .B1(G116), .B2(new_n212), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n241), .A2(G45), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n482), .A2(new_n693), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n753), .B1(new_n339), .B2(new_n207), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n750), .B1(new_n751), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n209), .B1(new_n269), .B2(G169), .ZN(new_n756));
  OR2_X1    g0556(.A1(new_n756), .A2(KEYINPUT98), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(KEYINPUT98), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(G13), .A2(G33), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(G20), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n745), .B1(new_n755), .B2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n759), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n269), .A2(new_n449), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G200), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n401), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n768), .A2(G190), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n415), .A2(new_n770), .B1(new_n772), .B2(new_n386), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n767), .A2(G190), .A3(new_n403), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G190), .A2(G200), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n767), .A2(new_n775), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n280), .B1(new_n774), .B2(new_n238), .C1(new_n216), .C2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n269), .A2(G179), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(new_n775), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n467), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT32), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n778), .A2(G190), .A3(G200), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n780), .A2(new_n781), .B1(new_n529), .B2(new_n782), .ZN(new_n783));
  NOR3_X1   g0583(.A1(new_n773), .A2(new_n777), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n780), .A2(new_n781), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n401), .A2(G179), .A3(G200), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n269), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(new_n249), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n778), .A2(new_n401), .A3(G200), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n788), .B1(G107), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n784), .A2(new_n785), .A3(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(G322), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n774), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G311), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n428), .B1(new_n776), .B2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n779), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n794), .B(new_n796), .C1(G329), .C2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n769), .A2(G326), .ZN(new_n799));
  XNOR2_X1  g0599(.A(KEYINPUT33), .B(G317), .ZN(new_n800));
  INV_X1    g0600(.A(new_n782), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n771), .A2(new_n800), .B1(new_n801), .B2(G303), .ZN(new_n802));
  INV_X1    g0602(.A(new_n787), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n803), .A2(G294), .B1(new_n790), .B2(G283), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n798), .A2(new_n799), .A3(new_n802), .A4(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n766), .B1(new_n792), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n765), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n762), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n807), .B1(new_n679), .B2(new_n808), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n747), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(G396));
  OAI21_X1  g0611(.A(new_n520), .B1(new_n513), .B2(new_n674), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(new_n523), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n523), .A2(new_n675), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n700), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n816), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n654), .A2(new_n674), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n739), .A2(G330), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n745), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(new_n821), .B2(new_n820), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n766), .A2(new_n761), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n745), .B1(new_n824), .B2(G77), .ZN(new_n825));
  INV_X1    g0625(.A(G283), .ZN(new_n826));
  INV_X1    g0626(.A(G303), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n826), .A2(new_n772), .B1(new_n770), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n828), .B1(G107), .B2(new_n801), .ZN(new_n829));
  INV_X1    g0629(.A(G294), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n774), .A2(new_n830), .B1(new_n779), .B2(new_n795), .ZN(new_n831));
  INV_X1    g0631(.A(new_n776), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n280), .B(new_n831), .C1(G116), .C2(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n789), .A2(new_n556), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n788), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n829), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n774), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n837), .A2(G143), .B1(new_n832), .B2(G159), .ZN(new_n838));
  INV_X1    g0638(.A(G137), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n838), .B1(new_n770), .B2(new_n839), .C1(new_n409), .C2(new_n772), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT34), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n482), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(G132), .B2(new_n797), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n782), .A2(new_n415), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n789), .A2(new_n386), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n845), .B(new_n846), .C1(G58), .C2(new_n803), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n842), .A2(new_n844), .A3(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n840), .A2(new_n841), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n836), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n825), .B1(new_n850), .B2(new_n759), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n818), .B2(new_n761), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n823), .A2(new_n852), .ZN(G384));
  INV_X1    g0653(.A(KEYINPUT40), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n675), .A2(new_n398), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n399), .A2(new_n406), .A3(new_n855), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n398), .B(new_n675), .C1(new_n385), .C2(new_n405), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n674), .B1(new_n729), .B2(new_n713), .ZN(new_n859));
  AOI21_X1  g0659(.A(KEYINPUT101), .B1(new_n859), .B2(KEYINPUT31), .ZN(new_n860));
  AND4_X1   g0660(.A1(KEYINPUT101), .A2(new_n734), .A3(KEYINPUT31), .A4(new_n675), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n738), .B(new_n737), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n858), .A2(new_n818), .A3(new_n862), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n484), .A2(new_n465), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n252), .B1(new_n484), .B2(new_n465), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n488), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n493), .B2(new_n672), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n489), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(KEYINPUT37), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n491), .A2(new_n672), .ZN(new_n870));
  XNOR2_X1  g0670(.A(KEYINPUT100), .B(KEYINPUT37), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n498), .A2(new_n870), .A3(new_n489), .A4(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n496), .A2(new_n495), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n657), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n665), .B1(new_n875), .B2(new_n500), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n866), .A2(new_n672), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n873), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT38), .ZN(new_n879));
  INV_X1    g0679(.A(new_n877), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n502), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n879), .B1(new_n869), .B2(new_n872), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n878), .A2(new_n879), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n854), .B1(new_n863), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n498), .A2(new_n870), .A3(new_n489), .ZN(new_n885));
  INV_X1    g0685(.A(new_n871), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n872), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n870), .B1(new_n490), .B2(new_n658), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n879), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n882), .B1(new_n876), .B2(new_n877), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n854), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n816), .B1(new_n856), .B2(new_n857), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n893), .A2(new_n894), .A3(new_n862), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n884), .A2(new_n895), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n525), .A2(new_n862), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n896), .A2(new_n897), .ZN(new_n899));
  INV_X1    g0699(.A(G330), .ZN(new_n900));
  NOR3_X1   g0700(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n883), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n819), .A2(new_n815), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n902), .A2(new_n858), .A3(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT39), .ZN(new_n905));
  INV_X1    g0705(.A(new_n872), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT37), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n907), .B1(new_n867), .B2(new_n489), .ZN(new_n908));
  OAI21_X1  g0708(.A(KEYINPUT38), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n909), .B1(new_n502), .B2(new_n880), .ZN(new_n910));
  INV_X1    g0710(.A(new_n870), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n657), .A2(new_n496), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n911), .B1(new_n912), .B2(new_n665), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT38), .B1(new_n913), .B2(new_n888), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n905), .B1(new_n910), .B2(new_n914), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n502), .A2(new_n880), .B1(new_n872), .B2(new_n869), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n892), .B(KEYINPUT39), .C1(new_n916), .C2(KEYINPUT38), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n399), .A2(new_n675), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n915), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n672), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n912), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n904), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n525), .A2(new_n706), .A3(new_n702), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n667), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n922), .B(new_n924), .Z(new_n925));
  OAI22_X1  g0725(.A1(new_n901), .A2(new_n925), .B1(new_n246), .B2(new_n742), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n926), .B1(new_n925), .B2(new_n901), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n266), .A2(KEYINPUT35), .ZN(new_n928));
  NOR3_X1   g0728(.A1(new_n208), .A2(new_n269), .A3(new_n549), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n266), .B2(KEYINPUT35), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT99), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(new_n931), .B2(new_n930), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT36), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n215), .B(new_n207), .C1(new_n238), .C2(new_n386), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n415), .A2(G68), .ZN(new_n936));
  AOI211_X1 g0736(.A(new_n246), .B(G13), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  OR3_X1    g0737(.A1(new_n927), .A2(new_n934), .A3(new_n937), .ZN(G367));
  INV_X1    g0738(.A(new_n745), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n763), .B1(new_n212), .B2(new_n503), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(new_n230), .B2(new_n752), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n769), .A2(G143), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n942), .B(new_n280), .C1(new_n216), .C2(new_n789), .ZN(new_n943));
  OAI22_X1  g0743(.A1(new_n772), .A2(new_n467), .B1(new_n776), .B2(new_n415), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n943), .B1(KEYINPUT107), .B2(new_n944), .ZN(new_n945));
  OAI22_X1  g0745(.A1(new_n787), .A2(new_n386), .B1(new_n774), .B2(new_n409), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n946), .B(KEYINPUT106), .Z(new_n947));
  NAND2_X1  g0747(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  OAI22_X1  g0748(.A1(new_n782), .A2(new_n238), .B1(new_n779), .B2(new_n839), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT108), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(KEYINPUT107), .B2(new_n944), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n789), .A2(new_n249), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  OAI221_X1 g0753(.A(new_n953), .B1(new_n257), .B2(new_n787), .C1(new_n772), .C2(new_n830), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n801), .A2(G116), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT46), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n774), .A2(new_n827), .B1(new_n776), .B2(new_n826), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(G317), .B2(new_n797), .ZN(new_n958));
  XOR2_X1   g0758(.A(KEYINPUT105), .B(G311), .Z(new_n959));
  AOI21_X1  g0759(.A(new_n482), .B1(new_n769), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n956), .A2(new_n958), .A3(new_n960), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n948), .A2(new_n951), .B1(new_n954), .B2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT47), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n964), .A2(new_n759), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n962), .A2(new_n963), .ZN(new_n966));
  AOI211_X1 g0766(.A(new_n939), .B(new_n941), .C1(new_n965), .C2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n557), .A2(new_n675), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n561), .B(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n967), .B1(new_n808), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n702), .A2(new_n706), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n821), .ZN(new_n973));
  XOR2_X1   g0773(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n974));
  NOR2_X1   g0774(.A1(new_n640), .A2(new_n674), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n284), .A2(new_n674), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n975), .B1(new_n335), .B2(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n974), .B1(new_n977), .B2(new_n690), .ZN(new_n978));
  NOR3_X1   g0778(.A1(new_n323), .A2(new_n325), .A3(KEYINPUT84), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n332), .B1(new_n331), .B2(new_n333), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n640), .B(new_n976), .C1(new_n979), .C2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n975), .ZN(new_n982));
  AND4_X1   g0782(.A1(new_n690), .A2(new_n981), .A3(new_n982), .A4(new_n974), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n978), .A2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT45), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n977), .B2(new_n690), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n981), .A2(new_n982), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n987), .A2(new_n691), .A3(KEYINPUT45), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  AND3_X1   g0789(.A1(new_n984), .A2(new_n688), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n688), .B1(new_n984), .B2(new_n989), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n689), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n683), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n687), .B2(new_n993), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n995), .A2(new_n681), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n681), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n973), .B1(new_n992), .B2(new_n998), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n694), .B(KEYINPUT41), .Z(new_n1000));
  OAI21_X1  g0800(.A(KEYINPUT104), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n688), .ZN(new_n1002));
  AND2_X1   g0802(.A1(new_n986), .A2(new_n988), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n974), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n987), .B2(new_n691), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n977), .A2(new_n690), .A3(new_n974), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1002), .B1(new_n1003), .B2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n984), .A2(new_n688), .A3(new_n989), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n998), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n740), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT104), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1000), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n744), .B1(new_n1001), .B2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n987), .A2(KEYINPUT42), .A3(new_n683), .A4(new_n993), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT42), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n977), .B2(new_n994), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n640), .B1(new_n981), .B2(new_n630), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n1017), .A2(new_n1019), .B1(new_n674), .B2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n970), .A2(KEYINPUT43), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT102), .ZN(new_n1024));
  AND2_X1   g0824(.A1(new_n970), .A2(KEYINPUT43), .ZN(new_n1025));
  OR3_X1    g0825(.A1(new_n1021), .A2(new_n1022), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n688), .A2(new_n977), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1024), .A2(new_n1028), .A3(new_n1026), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n971), .B1(new_n1016), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT109), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n740), .A2(new_n998), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1036));
  AOI211_X1 g0836(.A(KEYINPUT104), .B(new_n1000), .C1(new_n1036), .C2(new_n740), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1013), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n743), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1031), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1028), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1039), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1043), .A2(KEYINPUT109), .A3(new_n971), .ZN(new_n1044));
  AND2_X1   g0844(.A1(new_n1035), .A2(new_n1044), .ZN(G387));
  NAND3_X1  g0845(.A1(new_n686), .A2(new_n685), .A3(new_n762), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n953), .B1(new_n770), .B2(new_n467), .C1(new_n408), .C2(new_n772), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n843), .B(new_n1047), .C1(G68), .C2(new_n832), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n787), .A2(new_n503), .B1(new_n774), .B2(new_n415), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT112), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n216), .A2(new_n782), .B1(new_n409), .B2(new_n779), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT111), .Z(new_n1052));
  NAND3_X1  g0852(.A1(new_n1048), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n837), .A2(G317), .B1(new_n832), .B2(G303), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n771), .A2(new_n959), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1054), .B(new_n1055), .C1(new_n793), .C2(new_n770), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT48), .ZN(new_n1057));
  OR2_X1    g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n787), .A2(new_n826), .B1(new_n782), .B2(new_n830), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1058), .A2(KEYINPUT49), .A3(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n482), .B1(G326), .B2(new_n797), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1061), .B(new_n1062), .C1(new_n549), .C2(new_n789), .ZN(new_n1063));
  AOI21_X1  g0863(.A(KEYINPUT49), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1053), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n759), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n753), .B1(new_n235), .B2(G45), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(new_n697), .B2(new_n748), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n507), .A2(new_n415), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT50), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n339), .B1(new_n386), .B2(new_n203), .ZN(new_n1071));
  NOR3_X1   g0871(.A1(new_n1070), .A2(new_n697), .A3(new_n1071), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n1068), .A2(new_n1072), .B1(G107), .B2(new_n212), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n939), .B1(new_n1073), .B2(new_n763), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1066), .B1(KEYINPUT110), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(KEYINPUT110), .B2(new_n1074), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n998), .A2(new_n744), .B1(new_n1046), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n740), .A2(new_n998), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n694), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n740), .A2(new_n998), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1077), .B1(new_n1079), .B2(new_n1080), .ZN(G393));
  NAND2_X1  g0881(.A1(new_n991), .A2(KEYINPUT113), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n1010), .B2(KEYINPUT113), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1078), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n694), .B(new_n1036), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n771), .A2(G50), .B1(new_n832), .B2(new_n507), .ZN(new_n1086));
  XOR2_X1   g0886(.A(new_n1086), .B(KEYINPUT115), .Z(new_n1087));
  AOI21_X1  g0887(.A(new_n843), .B1(G143), .B2(new_n797), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n782), .A2(new_n386), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n834), .B(new_n1089), .C1(G77), .C2(new_n803), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1087), .A2(new_n1088), .A3(new_n1090), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(G150), .A2(new_n769), .B1(new_n837), .B2(G159), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT51), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(G317), .A2(new_n769), .B1(new_n837), .B2(G311), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT52), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n428), .B1(new_n779), .B2(new_n793), .C1(new_n830), .C2(new_n776), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n772), .A2(new_n827), .B1(new_n257), .B2(new_n789), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n787), .A2(new_n549), .B1(new_n782), .B2(new_n826), .ZN(new_n1099));
  NOR4_X1   g0899(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .A4(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n759), .B1(new_n1094), .B2(new_n1100), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n763), .B1(new_n249), .B2(new_n212), .C1(new_n244), .C2(new_n753), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT114), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n939), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1101), .B(new_n1104), .C1(new_n1103), .C2(new_n1102), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n977), .B2(new_n762), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(new_n1083), .B2(new_n744), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1085), .A2(new_n1107), .ZN(G390));
  AOI21_X1  g0908(.A(new_n918), .B1(new_n891), .B2(new_n892), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n814), .B1(new_n705), .B2(new_n813), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n858), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1109), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n739), .A2(new_n858), .A3(G330), .A4(new_n818), .ZN(new_n1113));
  AND2_X1   g0913(.A1(new_n915), .A2(new_n917), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n918), .B1(new_n903), .B2(new_n858), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1112), .B(new_n1113), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n918), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n678), .A2(new_n630), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1118), .A2(new_n335), .A3(new_n562), .A4(new_n633), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n675), .B1(new_n1119), .B2(new_n646), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n814), .B1(new_n1120), .B2(new_n818), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1117), .B1(new_n1121), .B2(new_n1111), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n915), .A2(new_n917), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n705), .A2(new_n813), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n815), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n858), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n1122), .A2(new_n1123), .B1(new_n1126), .B2(new_n1109), .ZN(new_n1127));
  AND2_X1   g0927(.A1(new_n862), .A2(G330), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n894), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1116), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(KEYINPUT116), .B1(new_n1130), .B2(new_n743), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1112), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1129), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT116), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1134), .A2(new_n1135), .A3(new_n744), .A4(new_n1116), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1131), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n525), .A2(new_n1128), .ZN(new_n1138));
  AND3_X1   g0938(.A1(new_n923), .A2(new_n667), .A3(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n862), .A2(G330), .A3(new_n818), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n1111), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1141), .A2(new_n1113), .A3(new_n1110), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n738), .A2(new_n737), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n736), .B(new_n674), .C1(new_n728), .C2(new_n731), .ZN(new_n1145));
  OAI211_X1 g0945(.A(G330), .B(new_n818), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n1111), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1121), .B1(new_n1129), .B2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1139), .B1(new_n1143), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1130), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1129), .A2(new_n1147), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n903), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n1142), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1134), .A2(new_n1153), .A3(new_n1116), .A4(new_n1139), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1150), .A2(new_n1154), .A3(new_n694), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n745), .B1(new_n824), .B2(new_n507), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n428), .B1(new_n782), .B2(new_n556), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1157), .B(KEYINPUT118), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n776), .A2(new_n249), .B1(new_n779), .B2(new_n830), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(G116), .B2(new_n837), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n846), .B1(G77), .B2(new_n803), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n771), .A2(G107), .B1(new_n769), .B2(G283), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1158), .A2(new_n1160), .A3(new_n1161), .A4(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(KEYINPUT54), .B(G143), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n803), .A2(G159), .B1(new_n832), .B2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1166), .B1(new_n839), .B2(new_n772), .ZN(new_n1167));
  XOR2_X1   g0967(.A(new_n1167), .B(KEYINPUT117), .Z(new_n1168));
  NAND2_X1  g0968(.A1(new_n801), .A2(G150), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT53), .ZN(new_n1170));
  INV_X1    g0970(.A(G125), .ZN(new_n1171));
  INV_X1    g0971(.A(G132), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n280), .B1(new_n779), .B2(new_n1171), .C1(new_n774), .C2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(G128), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n770), .A2(new_n1174), .B1(new_n415), .B2(new_n789), .ZN(new_n1175));
  OR3_X1    g0975(.A1(new_n1170), .A2(new_n1173), .A3(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1163), .B1(new_n1168), .B2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1156), .B1(new_n1177), .B2(new_n759), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n1114), .B2(new_n761), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1137), .A2(new_n1155), .A3(new_n1179), .ZN(G378));
  INV_X1    g0980(.A(new_n922), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n920), .B1(new_n414), .B2(new_n417), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT55), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n452), .A2(new_n1183), .ZN(new_n1184));
  XOR2_X1   g0984(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n1185));
  INV_X1    g0985(.A(new_n1183), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n446), .A2(new_n451), .A3(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1184), .A2(new_n1185), .A3(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1185), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1186), .B1(new_n446), .B2(new_n451), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n656), .B(new_n1183), .C1(new_n440), .C2(new_n445), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1189), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  AND2_X1   g0992(.A1(new_n1188), .A2(new_n1192), .ZN(new_n1193));
  AND4_X1   g0993(.A1(G330), .A2(new_n884), .A3(new_n895), .A4(new_n1193), .ZN(new_n1194));
  AND3_X1   g0994(.A1(new_n858), .A2(new_n818), .A3(new_n862), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n900), .B1(new_n1195), .B2(new_n893), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1193), .B1(new_n1196), .B2(new_n884), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1181), .B1(new_n1194), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1193), .ZN(new_n1199));
  AOI21_X1  g0999(.A(KEYINPUT40), .B1(new_n902), .B2(new_n1195), .ZN(new_n1200));
  OAI21_X1  g1000(.A(KEYINPUT40), .B1(new_n910), .B2(new_n914), .ZN(new_n1201));
  OAI21_X1  g1001(.A(G330), .B1(new_n1201), .B2(new_n863), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1199), .B1(new_n1200), .B2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1196), .A2(new_n884), .A3(new_n1193), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1203), .A2(new_n922), .A3(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1198), .A2(KEYINPUT121), .A3(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT121), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1207), .B(new_n1181), .C1(new_n1194), .C2(new_n1197), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1206), .A2(new_n744), .A3(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1193), .A2(new_n760), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n745), .B1(new_n824), .B2(G50), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n216), .A2(new_n782), .B1(new_n826), .B2(new_n779), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(G58), .B2(new_n790), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1213), .A2(new_n338), .A3(new_n843), .ZN(new_n1214));
  XOR2_X1   g1014(.A(new_n1214), .B(KEYINPUT119), .Z(new_n1215));
  OAI22_X1  g1015(.A1(new_n774), .A2(new_n257), .B1(new_n776), .B2(new_n503), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(G68), .B2(new_n803), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n771), .A2(G97), .B1(new_n769), .B2(G116), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1215), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT58), .ZN(new_n1220));
  OR2_X1    g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(G33), .A2(G41), .ZN(new_n1223));
  AOI211_X1 g1023(.A(G50), .B(new_n1223), .C1(new_n843), .C2(new_n338), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n1171), .A2(new_n770), .B1(new_n772), .B2(new_n1172), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(G150), .B2(new_n803), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n837), .A2(G128), .B1(new_n832), .B2(G137), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1226), .B(new_n1227), .C1(new_n782), .C2(new_n1164), .ZN(new_n1228));
  OR2_X1    g1028(.A1(new_n1228), .A2(KEYINPUT59), .ZN(new_n1229));
  INV_X1    g1029(.A(G124), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n1223), .B1(new_n779), .B2(new_n1230), .C1(new_n467), .C2(new_n789), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(new_n1228), .B2(KEYINPUT59), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1224), .B1(new_n1229), .B2(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1221), .A2(new_n1222), .A3(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1211), .B1(new_n1234), .B2(new_n759), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1210), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1209), .A2(new_n1236), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1143), .A2(new_n1148), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1139), .B1(new_n1130), .B2(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1206), .A2(new_n1239), .A3(new_n1208), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT57), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1241), .B1(new_n1198), .B2(new_n1205), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n695), .B1(new_n1243), .B2(new_n1239), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1237), .B1(new_n1242), .B2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(G375));
  NAND3_X1  g1046(.A1(new_n923), .A2(new_n1138), .A3(new_n667), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1238), .A2(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1248), .A2(new_n1014), .A3(new_n1149), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1111), .A2(new_n760), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n745), .B1(new_n824), .B2(G68), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n770), .A2(new_n830), .B1(new_n203), .B2(new_n789), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(G97), .B2(new_n801), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n774), .A2(new_n826), .B1(new_n779), .B2(new_n827), .ZN(new_n1254));
  AOI211_X1 g1054(.A(new_n280), .B(new_n1254), .C1(G107), .C2(new_n832), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n504), .A2(new_n803), .B1(new_n771), .B2(G116), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1253), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n843), .B1(G58), .B2(new_n790), .ZN(new_n1258));
  OAI22_X1  g1058(.A1(new_n776), .A2(new_n409), .B1(new_n779), .B2(new_n1174), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(G137), .B2(new_n837), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n769), .A2(G132), .B1(new_n801), .B2(G159), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(G50), .A2(new_n803), .B1(new_n771), .B2(new_n1165), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1258), .A2(new_n1260), .A3(new_n1261), .A4(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1257), .A2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1251), .B1(new_n1264), .B2(new_n759), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(new_n1153), .A2(new_n744), .B1(new_n1250), .B2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1249), .A2(new_n1266), .ZN(G381));
  INV_X1    g1067(.A(G390), .ZN(new_n1268));
  INV_X1    g1068(.A(G384), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  OR4_X1    g1070(.A1(G396), .A2(new_n1270), .A3(G393), .A4(G381), .ZN(new_n1271));
  OR4_X1    g1071(.A1(G387), .A2(G375), .A3(new_n1271), .A4(G378), .ZN(G407));
  OR3_X1    g1072(.A1(G375), .A2(G343), .A3(G378), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(G407), .A2(G213), .A3(new_n1273), .ZN(G409));
  XOR2_X1   g1074(.A(KEYINPUT125), .B(KEYINPUT61), .Z(new_n1275));
  INV_X1    g1075(.A(G213), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1276), .A2(G343), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1237), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1278), .A2(G378), .A3(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n743), .B1(new_n1198), .B2(new_n1205), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1281), .B1(new_n1210), .B2(new_n1235), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1206), .A2(new_n1239), .A3(new_n1014), .A4(new_n1208), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(G378), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1277), .B1(new_n1280), .B2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1277), .A2(G2897), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1149), .A2(KEYINPUT60), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(new_n1248), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1152), .A2(KEYINPUT60), .A3(new_n1247), .A4(new_n1142), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(new_n694), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1291), .A2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(G384), .B1(new_n1295), .B2(new_n1266), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1293), .B1(new_n1248), .B2(new_n1290), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1266), .ZN(new_n1298));
  NOR3_X1   g1098(.A1(new_n1297), .A2(new_n1269), .A3(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1289), .B1(new_n1296), .B2(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1295), .A2(G384), .A3(new_n1266), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1269), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1301), .A2(new_n1302), .A3(new_n1288), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1300), .A2(new_n1303), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1275), .B1(new_n1287), .B2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT126), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  OAI211_X1 g1107(.A(KEYINPUT126), .B(new_n1275), .C1(new_n1287), .C2(new_n1304), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1296), .A2(new_n1299), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1287), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(KEYINPUT62), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT62), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1287), .A2(new_n1312), .A3(new_n1309), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1307), .A2(new_n1308), .A3(new_n1311), .A4(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1035), .A2(new_n1044), .A3(new_n1268), .ZN(new_n1315));
  OAI211_X1 g1115(.A(G390), .B(new_n971), .C1(new_n1016), .C2(new_n1032), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT123), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  XNOR2_X1  g1119(.A(G393), .B(new_n810), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1320), .B1(new_n1316), .B2(KEYINPUT123), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1315), .A2(new_n1319), .A3(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(G390), .B1(new_n1043), .B2(new_n971), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1320), .B1(new_n1323), .B2(new_n1317), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1322), .A2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1314), .A2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT124), .ZN(new_n1328));
  OAI21_X1  g1128(.A(KEYINPUT122), .B1(new_n1287), .B2(new_n1304), .ZN(new_n1329));
  AND2_X1   g1129(.A1(new_n1300), .A2(new_n1303), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT122), .ZN(new_n1331));
  AOI21_X1  g1131(.A(G378), .B1(new_n1283), .B2(new_n1282), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1332), .B1(new_n1245), .B2(G378), .ZN(new_n1333));
  OAI211_X1 g1133(.A(new_n1330), .B(new_n1331), .C1(new_n1333), .C2(new_n1277), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1329), .A2(new_n1334), .ZN(new_n1335));
  AOI21_X1  g1135(.A(KEYINPUT63), .B1(new_n1287), .B2(new_n1309), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1280), .A2(new_n1286), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1277), .ZN(new_n1339));
  AND3_X1   g1139(.A1(new_n1301), .A2(new_n1302), .A3(KEYINPUT63), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1338), .A2(new_n1339), .A3(new_n1340), .ZN(new_n1341));
  AOI21_X1  g1141(.A(KEYINPUT61), .B1(new_n1322), .B2(new_n1324), .ZN(new_n1342));
  AND2_X1   g1142(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1343));
  AND4_X1   g1143(.A1(new_n1328), .A2(new_n1335), .A3(new_n1337), .A4(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1345));
  NOR2_X1   g1145(.A1(new_n1345), .A2(new_n1336), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1328), .B1(new_n1346), .B2(new_n1335), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1327), .B1(new_n1344), .B2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1348), .A2(KEYINPUT127), .ZN(new_n1349));
  INV_X1    g1149(.A(KEYINPUT127), .ZN(new_n1350));
  OAI211_X1 g1150(.A(new_n1327), .B(new_n1350), .C1(new_n1344), .C2(new_n1347), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1349), .A2(new_n1351), .ZN(G405));
  XNOR2_X1  g1152(.A(new_n1245), .B(new_n1285), .ZN(new_n1353));
  XNOR2_X1  g1153(.A(new_n1353), .B(new_n1309), .ZN(new_n1354));
  XNOR2_X1  g1154(.A(new_n1354), .B(new_n1325), .ZN(G402));
endmodule


