//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 1 1 1 1 1 1 1 1 1 1 1 0 0 1 1 0 0 0 0 1 1 1 0 1 0 1 1 0 0 0 1 1 1 1 1 1 0 0 1 0 0 0 0 1 1 0 0 1 0 1 1 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:35 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n449, new_n451, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n556, new_n557,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n571, new_n574, new_n575,
    new_n576, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1144;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g020(.A(KEYINPUT65), .B(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n448));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  INV_X1    g025(.A(new_n449), .ZN(new_n451));
  NAND2_X1  g026(.A1(new_n451), .A2(G567), .ZN(G234));
  NAND2_X1  g027(.A1(new_n451), .A2(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT68), .ZN(new_n455));
  XNOR2_X1  g030(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n455), .B(new_n456), .ZN(new_n457));
  NAND4_X1  g032(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n457), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  NAND2_X1  g035(.A1(new_n457), .A2(G2106), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(new_n462));
  OR2_X1    g037(.A1(new_n462), .A2(KEYINPUT69), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n458), .A2(G567), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n462), .A2(KEYINPUT69), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(G319));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n468), .A2(G101), .A3(G2104), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  AND2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(KEYINPUT70), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT70), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n472), .B(new_n477), .C1(new_n474), .C2(new_n473), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n470), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g054(.A(G125), .B1(new_n473), .B2(new_n474), .ZN(new_n480));
  NAND2_X1  g055(.A1(G113), .A2(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n479), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G160));
  OR2_X1    g060(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n486));
  NAND2_X1  g061(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n487));
  AOI21_X1  g062(.A(G2105), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G136), .ZN(new_n489));
  XNOR2_X1  g064(.A(new_n489), .B(KEYINPUT71), .ZN(new_n490));
  XNOR2_X1  g065(.A(KEYINPUT3), .B(G2104), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n491), .A2(G124), .A3(G2105), .ZN(new_n492));
  XNOR2_X1  g067(.A(new_n492), .B(KEYINPUT72), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n468), .A2(G112), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n490), .B(new_n493), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT73), .ZN(new_n497));
  XNOR2_X1  g072(.A(new_n496), .B(new_n497), .ZN(G162));
  OR2_X1    g073(.A1(G102), .A2(G2105), .ZN(new_n499));
  OAI21_X1  g074(.A(G2105), .B1(KEYINPUT74), .B2(G114), .ZN(new_n500));
  AND2_X1   g075(.A1(KEYINPUT74), .A2(G114), .ZN(new_n501));
  OAI211_X1 g076(.A(G2104), .B(new_n499), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  OAI211_X1 g077(.A(G126), .B(G2105), .C1(new_n473), .C2(new_n474), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT75), .ZN(new_n505));
  OAI211_X1 g080(.A(G138), .B(new_n468), .C1(new_n473), .C2(new_n474), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT4), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT4), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n491), .A2(new_n508), .A3(G138), .A4(new_n468), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT75), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n502), .A2(new_n503), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n505), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(G164));
  INV_X1    g089(.A(G62), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT76), .A2(KEYINPUT5), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(KEYINPUT76), .A2(KEYINPUT5), .A3(G543), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n515), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(G75), .A2(G543), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  OAI21_X1  g097(.A(G651), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n518), .A2(new_n519), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT6), .B(G651), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n524), .A2(G88), .A3(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n525), .A2(G50), .A3(G543), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n523), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(G166));
  NAND3_X1  g104(.A1(new_n524), .A2(G63), .A3(G651), .ZN(new_n530));
  XOR2_X1   g105(.A(new_n530), .B(KEYINPUT77), .Z(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n525), .A2(G543), .ZN(new_n534));
  INV_X1    g109(.A(G51), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n524), .A2(new_n525), .ZN(new_n536));
  INV_X1    g111(.A(G89), .ZN(new_n537));
  OAI221_X1 g112(.A(new_n533), .B1(new_n534), .B2(new_n535), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n531), .A2(new_n538), .ZN(G168));
  AOI22_X1  g114(.A1(new_n524), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  INV_X1    g115(.A(G651), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(G90), .ZN(new_n543));
  INV_X1    g118(.A(G52), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n536), .A2(new_n543), .B1(new_n534), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n542), .A2(new_n545), .ZN(G171));
  AOI22_X1  g121(.A1(new_n524), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(new_n541), .ZN(new_n548));
  AND2_X1   g123(.A1(new_n524), .A2(new_n525), .ZN(new_n549));
  XNOR2_X1  g124(.A(KEYINPUT78), .B(G81), .ZN(new_n550));
  AND2_X1   g125(.A1(new_n525), .A2(G543), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n549), .A2(new_n550), .B1(new_n551), .B2(G43), .ZN(new_n552));
  AND2_X1   g127(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  NAND4_X1  g129(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(G188));
  INV_X1    g133(.A(G65), .ZN(new_n559));
  AND2_X1   g134(.A1(new_n518), .A2(new_n519), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT79), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n524), .A2(KEYINPUT79), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n559), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AND2_X1   g139(.A1(G78), .A2(G543), .ZN(new_n565));
  OAI21_X1  g140(.A(G651), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n525), .A2(G53), .A3(G543), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT9), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n549), .A2(G91), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n566), .A2(new_n568), .A3(new_n569), .ZN(G299));
  XNOR2_X1  g145(.A(G171), .B(KEYINPUT80), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(G301));
  OR2_X1    g147(.A1(new_n531), .A2(new_n538), .ZN(G286));
  NAND2_X1  g148(.A1(new_n528), .A2(KEYINPUT81), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT81), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n523), .A2(new_n575), .A3(new_n526), .A4(new_n527), .ZN(new_n576));
  AND2_X1   g151(.A1(new_n574), .A2(new_n576), .ZN(G303));
  AOI22_X1  g152(.A1(new_n549), .A2(G87), .B1(new_n551), .B2(G49), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n524), .B2(G74), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(G288));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  INV_X1    g156(.A(G61), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n560), .B2(new_n582), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n583), .A2(G651), .B1(new_n549), .B2(G86), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n525), .A2(G48), .A3(G543), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT82), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n585), .B(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n584), .A2(new_n587), .ZN(G305));
  AOI22_X1  g163(.A1(new_n524), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n589), .A2(new_n541), .ZN(new_n590));
  INV_X1    g165(.A(G85), .ZN(new_n591));
  INV_X1    g166(.A(G47), .ZN(new_n592));
  OAI22_X1  g167(.A1(new_n536), .A2(new_n591), .B1(new_n534), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(G290));
  INV_X1    g170(.A(G66), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n596), .B1(new_n562), .B2(new_n563), .ZN(new_n597));
  AND2_X1   g172(.A1(G79), .A2(G543), .ZN(new_n598));
  OAI21_X1  g173(.A(G651), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n549), .A2(KEYINPUT10), .A3(G92), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT10), .ZN(new_n601));
  INV_X1    g176(.A(G92), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n536), .B2(new_n602), .ZN(new_n603));
  OR2_X1    g178(.A1(new_n534), .A2(KEYINPUT83), .ZN(new_n604));
  INV_X1    g179(.A(G54), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n605), .B1(new_n534), .B2(KEYINPUT83), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n600), .A2(new_n603), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n599), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n608), .A2(G868), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n609), .B1(G868), .B2(new_n571), .ZN(G284));
  AOI21_X1  g185(.A(new_n609), .B1(G868), .B2(new_n571), .ZN(G321));
  MUX2_X1   g186(.A(G299), .B(G286), .S(G868), .Z(G297));
  XNOR2_X1  g187(.A(G297), .B(KEYINPUT84), .ZN(G280));
  INV_X1    g188(.A(new_n608), .ZN(new_n614));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(G860), .ZN(G148));
  NAND2_X1  g191(.A1(new_n614), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(G868), .ZN(new_n618));
  OR2_X1    g193(.A1(new_n618), .A2(KEYINPUT85), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(KEYINPUT85), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n619), .B(new_n620), .C1(G868), .C2(new_n553), .ZN(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g197(.A1(new_n491), .A2(G2105), .ZN(new_n623));
  INV_X1    g198(.A(G123), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n468), .A2(G111), .ZN(new_n625));
  OAI21_X1  g200(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n626));
  OAI22_X1  g201(.A1(new_n623), .A2(new_n624), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n627), .B1(G135), .B2(new_n488), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT86), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n629), .A2(G2096), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(G2096), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n468), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT12), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT13), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2100), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n630), .A2(new_n631), .A3(new_n635), .ZN(G156));
  XNOR2_X1  g211(.A(KEYINPUT87), .B(KEYINPUT14), .ZN(new_n637));
  XOR2_X1   g212(.A(KEYINPUT15), .B(G2435), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2438), .ZN(new_n639));
  XOR2_X1   g214(.A(G2427), .B(G2430), .Z(new_n640));
  AOI21_X1  g215(.A(new_n637), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(new_n639), .B2(new_n640), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2451), .B(G2454), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(G1341), .B(G1348), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n642), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n647), .A2(new_n648), .ZN(new_n650));
  AND3_X1   g225(.A1(new_n649), .A2(G14), .A3(new_n650), .ZN(G401));
  XOR2_X1   g226(.A(G2072), .B(G2078), .Z(new_n652));
  INV_X1    g227(.A(KEYINPUT89), .ZN(new_n653));
  AND2_X1   g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  NOR3_X1   g231(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n657), .B1(new_n653), .B2(new_n652), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n652), .A2(KEYINPUT17), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n652), .A2(KEYINPUT17), .ZN(new_n660));
  OAI211_X1 g235(.A(new_n659), .B(new_n660), .C1(new_n655), .C2(new_n656), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n655), .A2(new_n656), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n658), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n662), .A2(new_n652), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT88), .B(KEYINPUT18), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n664), .A2(new_n665), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n663), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2096), .B(G2100), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(G227));
  XOR2_X1   g245(.A(G1971), .B(G1976), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT19), .ZN(new_n672));
  XOR2_X1   g247(.A(G1956), .B(G2474), .Z(new_n673));
  XOR2_X1   g248(.A(G1961), .B(G1966), .Z(new_n674));
  AND2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT20), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n673), .A2(new_n674), .ZN(new_n678));
  NOR3_X1   g253(.A1(new_n672), .A2(new_n675), .A3(new_n678), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n679), .B1(new_n672), .B2(new_n678), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1981), .B(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(G229));
  INV_X1    g262(.A(G29), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(G35), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(KEYINPUT98), .Z(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(G162), .B2(new_n688), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT29), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G2090), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT99), .ZN(new_n694));
  MUX2_X1   g269(.A(G21), .B(G286), .S(G16), .Z(new_n695));
  NAND2_X1  g270(.A1(new_n553), .A2(G16), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(G16), .B2(G19), .ZN(new_n697));
  INV_X1    g272(.A(G1341), .ZN(new_n698));
  AOI22_X1  g273(.A1(new_n695), .A2(G1966), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(G2084), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n688), .B1(KEYINPUT24), .B2(G34), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(KEYINPUT24), .B2(G34), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(new_n484), .B2(G29), .ZN(new_n703));
  OAI221_X1 g278(.A(new_n699), .B1(G1966), .B2(new_n695), .C1(new_n700), .C2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n688), .A2(G32), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n468), .A2(G105), .A3(G2104), .ZN(new_n706));
  NAND3_X1  g281(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT26), .Z(new_n708));
  NAND2_X1  g283(.A1(new_n488), .A2(G141), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n491), .A2(G129), .A3(G2105), .ZN(new_n710));
  AND4_X1   g285(.A1(new_n706), .A2(new_n708), .A3(new_n709), .A4(new_n710), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n705), .B1(new_n711), .B2(new_n688), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT27), .B(G1996), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT94), .ZN(new_n716));
  OAI22_X1  g291(.A1(new_n697), .A2(new_n698), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n488), .A2(G140), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n468), .A2(G116), .ZN(new_n719));
  OAI21_X1  g294(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n720));
  INV_X1    g295(.A(G128), .ZN(new_n721));
  OAI221_X1 g296(.A(new_n718), .B1(new_n719), .B2(new_n720), .C1(new_n721), .C2(new_n623), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G29), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n688), .A2(G26), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT28), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G2067), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(new_n715), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n728), .B1(KEYINPUT94), .B2(new_n729), .ZN(new_n730));
  NOR3_X1   g305(.A1(new_n704), .A2(new_n717), .A3(new_n730), .ZN(new_n731));
  MUX2_X1   g306(.A(G4), .B(new_n608), .S(G16), .Z(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT92), .Z(new_n733));
  XOR2_X1   g308(.A(KEYINPUT91), .B(G1348), .Z(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n733), .A2(new_n735), .ZN(new_n737));
  INV_X1    g312(.A(G5), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n738), .A2(G16), .ZN(new_n739));
  INV_X1    g314(.A(G171), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n739), .B1(new_n740), .B2(G16), .ZN(new_n741));
  INV_X1    g316(.A(G1961), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT95), .Z(new_n744));
  NAND4_X1  g319(.A1(new_n731), .A2(new_n736), .A3(new_n737), .A4(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT100), .B(KEYINPUT23), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT101), .ZN(new_n747));
  INV_X1    g322(.A(G20), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n748), .A2(G16), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n747), .B(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G299), .B2(G16), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G1956), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT25), .ZN(new_n753));
  NAND2_X1  g328(.A1(G103), .A2(G2104), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n753), .B1(new_n754), .B2(G2105), .ZN(new_n755));
  NAND4_X1  g330(.A1(new_n468), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n488), .A2(G139), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n491), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n757), .B1(new_n468), .B2(new_n758), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT93), .ZN(new_n760));
  MUX2_X1   g335(.A(G33), .B(new_n760), .S(G29), .Z(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(G2072), .Z(new_n762));
  INV_X1    g337(.A(G28), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n763), .A2(KEYINPUT30), .ZN(new_n764));
  AOI21_X1  g339(.A(G29), .B1(new_n763), .B2(KEYINPUT30), .ZN(new_n765));
  OR2_X1    g340(.A1(KEYINPUT31), .A2(G11), .ZN(new_n766));
  NAND2_X1  g341(.A1(KEYINPUT31), .A2(G11), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n764), .A2(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n629), .B2(new_n688), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n712), .B2(new_n714), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n741), .A2(new_n742), .B1(new_n700), .B2(new_n703), .ZN(new_n771));
  AND4_X1   g346(.A1(new_n752), .A2(new_n762), .A3(new_n770), .A4(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n688), .A2(G27), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT96), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G164), .B2(new_n688), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G2078), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT97), .ZN(new_n777));
  OAI211_X1 g352(.A(new_n772), .B(new_n777), .C1(G2090), .C2(new_n692), .ZN(new_n778));
  NOR3_X1   g353(.A1(new_n694), .A2(new_n745), .A3(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT102), .ZN(new_n780));
  MUX2_X1   g355(.A(G23), .B(G288), .S(G16), .Z(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT33), .B(G1976), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT90), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  MUX2_X1   g360(.A(G22), .B(new_n528), .S(G16), .Z(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(G1971), .Z(new_n787));
  NAND3_X1  g362(.A1(new_n584), .A2(new_n587), .A3(G16), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G6), .B2(G16), .ZN(new_n789));
  XOR2_X1   g364(.A(KEYINPUT32), .B(G1981), .Z(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n789), .A2(new_n790), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n787), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  OR3_X1    g368(.A1(new_n785), .A2(KEYINPUT34), .A3(new_n793), .ZN(new_n794));
  OAI21_X1  g369(.A(KEYINPUT34), .B1(new_n785), .B2(new_n793), .ZN(new_n795));
  MUX2_X1   g370(.A(G24), .B(G290), .S(G16), .Z(new_n796));
  AND2_X1   g371(.A1(new_n796), .A2(G1986), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n796), .A2(G1986), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n488), .A2(G131), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n468), .A2(G107), .ZN(new_n800));
  OAI21_X1  g375(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n801));
  INV_X1    g376(.A(G119), .ZN(new_n802));
  OAI221_X1 g377(.A(new_n799), .B1(new_n800), .B2(new_n801), .C1(new_n802), .C2(new_n623), .ZN(new_n803));
  MUX2_X1   g378(.A(G25), .B(new_n803), .S(G29), .Z(new_n804));
  XOR2_X1   g379(.A(KEYINPUT35), .B(G1991), .Z(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n804), .B(new_n806), .ZN(new_n807));
  NOR3_X1   g382(.A1(new_n797), .A2(new_n798), .A3(new_n807), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n794), .A2(new_n795), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n809), .A2(KEYINPUT36), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT36), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n794), .A2(new_n811), .A3(new_n795), .A4(new_n808), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  AND3_X1   g388(.A1(new_n779), .A2(new_n780), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n780), .B1(new_n779), .B2(new_n813), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n814), .A2(new_n815), .ZN(G311));
  NAND2_X1  g391(.A1(new_n779), .A2(new_n813), .ZN(G150));
  NOR2_X1   g392(.A1(new_n608), .A2(new_n615), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n524), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n821), .A2(new_n541), .ZN(new_n822));
  INV_X1    g397(.A(G93), .ZN(new_n823));
  INV_X1    g398(.A(G55), .ZN(new_n824));
  OAI22_X1  g399(.A1(new_n536), .A2(new_n823), .B1(new_n534), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n553), .B(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n820), .B(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT39), .ZN(new_n830));
  AOI21_X1  g405(.A(G860), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(new_n830), .B2(new_n829), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n827), .A2(G860), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT37), .Z(new_n834));
  NAND2_X1  g409(.A1(new_n832), .A2(new_n834), .ZN(G145));
  XNOR2_X1  g410(.A(new_n629), .B(KEYINPUT104), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(G160), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(G162), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n504), .B1(new_n507), .B2(new_n509), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n722), .B(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(new_n711), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(new_n759), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n842), .B1(new_n760), .B2(new_n841), .ZN(new_n843));
  INV_X1    g418(.A(G130), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n468), .A2(G118), .ZN(new_n845));
  OAI21_X1  g420(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n846));
  OAI22_X1  g421(.A1(new_n623), .A2(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n847), .B1(G142), .B2(new_n488), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n848), .B(new_n633), .Z(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n803), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n843), .B(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(G37), .B1(new_n838), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(new_n838), .B2(new_n851), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g429(.A(G305), .B(new_n594), .ZN(new_n855));
  XNOR2_X1  g430(.A(G288), .B(G166), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n857), .A2(KEYINPUT42), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT106), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT42), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n857), .B(KEYINPUT105), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n859), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(G299), .B(new_n608), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT41), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n865), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n828), .B(new_n617), .ZN(new_n869));
  MUX2_X1   g444(.A(new_n864), .B(new_n868), .S(new_n869), .Z(new_n870));
  XNOR2_X1  g445(.A(new_n863), .B(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(G868), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n872), .B1(G868), .B2(new_n826), .ZN(G295));
  OAI21_X1  g448(.A(new_n872), .B1(G868), .B2(new_n826), .ZN(G331));
  NOR2_X1   g449(.A1(G168), .A2(G171), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n875), .B1(G168), .B2(new_n571), .ZN(new_n876));
  INV_X1    g451(.A(new_n828), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n876), .A2(new_n877), .ZN(new_n879));
  NAND4_X1  g454(.A1(new_n878), .A2(new_n866), .A3(new_n867), .A4(new_n879), .ZN(new_n880));
  AND2_X1   g455(.A1(new_n878), .A2(new_n879), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n880), .B1(new_n881), .B2(new_n864), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(new_n862), .ZN(new_n883));
  INV_X1    g458(.A(G37), .ZN(new_n884));
  OAI211_X1 g459(.A(new_n861), .B(new_n880), .C1(new_n864), .C2(new_n881), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(KEYINPUT43), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT43), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n883), .A2(new_n888), .A3(new_n885), .A4(new_n884), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT107), .ZN(new_n891));
  AOI21_X1  g466(.A(KEYINPUT44), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT44), .ZN(new_n893));
  AOI211_X1 g468(.A(KEYINPUT107), .B(new_n893), .C1(new_n887), .C2(new_n889), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n892), .A2(new_n894), .ZN(G397));
  INV_X1    g470(.A(G1384), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n513), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT45), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(G40), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n900), .B1(new_n482), .B2(G2105), .ZN(new_n901));
  AND3_X1   g476(.A1(new_n479), .A2(new_n901), .A3(KEYINPUT109), .ZN(new_n902));
  AOI21_X1  g477(.A(KEYINPUT109), .B1(new_n479), .B2(new_n901), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(G2078), .ZN(new_n905));
  AND2_X1   g480(.A1(new_n502), .A2(new_n503), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n510), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n907), .A2(KEYINPUT45), .A3(new_n896), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n899), .A2(new_n904), .A3(new_n905), .A4(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT53), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n897), .A2(KEYINPUT50), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(new_n904), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT50), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n907), .A2(new_n914), .A3(new_n896), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(KEYINPUT112), .ZN(new_n916));
  AOI21_X1  g491(.A(G1384), .B1(new_n510), .B2(new_n906), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT112), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n917), .A2(new_n918), .A3(new_n914), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n742), .B1(new_n913), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n513), .A2(KEYINPUT45), .A3(new_n896), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n898), .B1(new_n839), .B2(G1384), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT109), .ZN(new_n924));
  INV_X1    g499(.A(new_n478), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n477), .B1(new_n491), .B2(new_n472), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n469), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n481), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n928), .B1(new_n491), .B2(G125), .ZN(new_n929));
  OAI21_X1  g504(.A(G40), .B1(new_n929), .B2(new_n468), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n924), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n479), .A2(new_n901), .A3(KEYINPUT109), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n922), .A2(new_n923), .A3(new_n931), .A4(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n905), .A2(KEYINPUT53), .ZN(new_n934));
  OR2_X1    g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n911), .A2(new_n921), .A3(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT122), .ZN(new_n937));
  AND3_X1   g512(.A1(new_n936), .A2(new_n937), .A3(new_n571), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n937), .B1(new_n936), .B2(new_n571), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n907), .A2(new_n896), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT108), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT45), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n943), .B1(new_n942), .B2(new_n941), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n479), .A2(new_n901), .ZN(new_n945));
  AOI211_X1 g520(.A(new_n934), .B(new_n945), .C1(KEYINPUT45), .C2(new_n917), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n911), .A2(new_n921), .A3(G301), .A4(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n948), .B(KEYINPUT123), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT54), .B1(new_n940), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT51), .ZN(new_n951));
  NAND2_X1  g526(.A1(G286), .A2(G8), .ZN(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n951), .B1(new_n953), .B2(KEYINPUT121), .ZN(new_n954));
  INV_X1    g529(.A(G1966), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n933), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(KEYINPUT115), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT115), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n933), .A2(new_n958), .A3(new_n955), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n912), .A2(new_n904), .A3(new_n916), .A4(new_n919), .ZN(new_n960));
  OAI211_X1 g535(.A(new_n957), .B(new_n959), .C1(G2084), .C2(new_n960), .ZN(new_n961));
  OAI211_X1 g536(.A(G8), .B(new_n954), .C1(new_n961), .C2(G286), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n959), .B1(new_n960), .B2(G2084), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n958), .B1(new_n933), .B2(new_n955), .ZN(new_n964));
  OAI21_X1  g539(.A(G8), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n965), .A2(KEYINPUT121), .A3(new_n951), .A4(new_n952), .ZN(new_n966));
  OAI211_X1 g541(.A(G8), .B(G286), .C1(new_n963), .C2(new_n964), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT120), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT120), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n961), .A2(new_n969), .A3(G8), .A4(G286), .ZN(new_n970));
  AOI22_X1  g545(.A1(new_n962), .A2(new_n966), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n904), .A2(new_n917), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n578), .A2(G1976), .A3(new_n579), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n972), .A2(G8), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT52), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT49), .ZN(new_n976));
  INV_X1    g551(.A(G1981), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n584), .A2(new_n587), .A3(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n977), .B1(new_n584), .B2(new_n587), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n976), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n980), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n982), .A2(KEYINPUT49), .A3(new_n978), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n981), .A2(new_n983), .A3(G8), .A4(new_n972), .ZN(new_n984));
  INV_X1    g559(.A(G1976), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT52), .B1(G288), .B2(new_n985), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n972), .A2(G8), .A3(new_n973), .A4(new_n986), .ZN(new_n987));
  AND3_X1   g562(.A1(new_n975), .A2(new_n984), .A3(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n574), .A2(G8), .A3(new_n576), .ZN(new_n989));
  NAND2_X1  g564(.A1(KEYINPUT113), .A2(KEYINPUT55), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT114), .ZN(new_n992));
  XNOR2_X1  g567(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n574), .A2(new_n576), .A3(G8), .A4(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n991), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n992), .B1(new_n991), .B2(new_n994), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n908), .A2(new_n931), .A3(new_n932), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT45), .B1(new_n513), .B2(new_n896), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n513), .A2(new_n914), .A3(new_n896), .ZN(new_n1002));
  OAI21_X1  g577(.A(KEYINPUT50), .B1(new_n839), .B2(G1384), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n1002), .A2(new_n1003), .A3(new_n931), .A4(new_n932), .ZN(new_n1004));
  OAI22_X1  g579(.A1(new_n1001), .A2(G1971), .B1(new_n1004), .B2(G2090), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(G8), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n998), .A2(new_n1006), .ZN(new_n1007));
  OAI22_X1  g582(.A1(new_n960), .A2(G2090), .B1(new_n1001), .B2(G1971), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n1008), .B(G8), .C1(new_n996), .C2(new_n997), .ZN(new_n1009));
  AND3_X1   g584(.A1(new_n988), .A2(new_n1007), .A3(new_n1009), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n911), .A2(new_n921), .A3(new_n947), .ZN(new_n1011));
  OAI221_X1 g586(.A(KEYINPUT54), .B1(new_n936), .B2(new_n571), .C1(new_n1011), .C2(new_n740), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  NOR3_X1   g588(.A1(new_n950), .A2(new_n971), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT61), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT117), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n568), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT57), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  XOR2_X1   g594(.A(G299), .B(new_n1019), .Z(new_n1020));
  XOR2_X1   g595(.A(KEYINPUT56), .B(G2072), .Z(new_n1021));
  NOR3_X1   g596(.A1(new_n999), .A2(new_n1000), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT118), .ZN(new_n1023));
  INV_X1    g598(.A(G1956), .ZN(new_n1024));
  AOI22_X1  g599(.A1(new_n1022), .A2(new_n1023), .B1(new_n1024), .B2(new_n1004), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1021), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n899), .A2(new_n904), .A3(new_n908), .A4(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT118), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1020), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1004), .A2(new_n1024), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1030), .B1(new_n1027), .B2(KEYINPUT118), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1023), .B1(new_n1001), .B2(new_n1026), .ZN(new_n1032));
  XNOR2_X1  g607(.A(G299), .B(new_n1019), .ZN(new_n1033));
  NOR3_X1   g608(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1015), .B1(new_n1029), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n931), .A2(new_n932), .ZN(new_n1036));
  NOR3_X1   g611(.A1(new_n1036), .A2(G2067), .A3(new_n941), .ZN(new_n1037));
  INV_X1    g612(.A(G1348), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1037), .B1(new_n960), .B2(new_n1038), .ZN(new_n1039));
  OR2_X1    g614(.A1(new_n1039), .A2(KEYINPUT60), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n960), .A2(new_n1038), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1037), .ZN(new_n1042));
  AND4_X1   g617(.A1(KEYINPUT60), .A2(new_n1041), .A3(new_n608), .A4(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n608), .B1(new_n1039), .B2(KEYINPUT60), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1040), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1036), .A2(new_n941), .ZN(new_n1046));
  XNOR2_X1  g621(.A(KEYINPUT58), .B(G1341), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NOR3_X1   g623(.A1(new_n999), .A2(G1996), .A3(new_n1000), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n553), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n1050), .B(KEYINPUT59), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1033), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1025), .A2(new_n1020), .A3(new_n1028), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1052), .A2(new_n1053), .A3(KEYINPUT61), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1035), .A2(new_n1045), .A3(new_n1051), .A4(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1039), .A2(new_n608), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1029), .B1(new_n1053), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT119), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1055), .A2(KEYINPUT119), .A3(new_n1057), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1014), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n988), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n972), .A2(G8), .ZN(new_n1064));
  NOR2_X1   g639(.A1(G288), .A2(G1976), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n979), .B1(new_n984), .B2(new_n1065), .ZN(new_n1066));
  OAI22_X1  g641(.A1(new_n1063), .A2(new_n1009), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n961), .A2(G8), .A3(G168), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1010), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n988), .A2(new_n1007), .A3(new_n1009), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT116), .B1(new_n1072), .B2(new_n1069), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT63), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1071), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1008), .A2(G8), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1074), .B1(new_n1076), .B2(new_n998), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1070), .A2(new_n1077), .A3(new_n1009), .A4(new_n988), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1067), .B1(new_n1075), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT124), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n940), .A2(new_n1072), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT62), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1081), .B1(new_n971), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n966), .A2(new_n962), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n968), .A2(new_n970), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1084), .A2(new_n1082), .A3(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1080), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(KEYINPUT62), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n971), .A2(new_n1082), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1089), .A2(new_n1090), .A3(KEYINPUT124), .A4(new_n1081), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1062), .A2(new_n1079), .A3(new_n1087), .A4(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n944), .A2(new_n1036), .ZN(new_n1093));
  INV_X1    g668(.A(G1996), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(KEYINPUT110), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT110), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1093), .A2(new_n1097), .A3(new_n1094), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1099), .A2(KEYINPUT111), .A3(new_n711), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT111), .B1(new_n1099), .B2(new_n711), .ZN(new_n1101));
  OR2_X1    g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g677(.A(new_n722), .B(new_n727), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1103), .B1(new_n1094), .B2(new_n711), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1093), .A2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n803), .A2(new_n806), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n803), .A2(new_n806), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1093), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1102), .A2(new_n1105), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(G1986), .ZN(new_n1110));
  XNOR2_X1  g685(.A(new_n594), .B(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1109), .B1(new_n1093), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1092), .A2(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT125), .B(KEYINPUT47), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT46), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1099), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1096), .A2(KEYINPUT46), .A3(new_n1098), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1103), .A2(new_n711), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1093), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1114), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1120), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1114), .ZN(new_n1123));
  AOI211_X1 g698(.A(new_n1122), .B(new_n1123), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1124));
  OAI21_X1  g699(.A(KEYINPUT126), .B1(new_n1121), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1117), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT46), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1120), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n1123), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT126), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1118), .A2(new_n1120), .A3(new_n1114), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1129), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1125), .A2(new_n1132), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1105), .B(new_n1106), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1134), .B1(G2067), .B2(new_n722), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(new_n1093), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1093), .A2(new_n1110), .A3(new_n594), .ZN(new_n1137));
  XNOR2_X1  g712(.A(new_n1137), .B(KEYINPUT127), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n1138), .B(KEYINPUT48), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1102), .A2(new_n1139), .A3(new_n1105), .A4(new_n1108), .ZN(new_n1140));
  AND3_X1   g715(.A1(new_n1133), .A2(new_n1136), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1113), .A2(new_n1141), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g717(.A1(G229), .A2(new_n466), .A3(G401), .A4(G227), .ZN(new_n1144));
  NAND3_X1  g718(.A1(new_n890), .A2(new_n853), .A3(new_n1144), .ZN(G225));
  INV_X1    g719(.A(G225), .ZN(G308));
endmodule


