

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774;

  OR2_X1 U373 ( .A1(n709), .A2(n590), .ZN(n365) );
  NOR2_X1 U374 ( .A1(n696), .A2(n697), .ZN(n585) );
  XNOR2_X1 U375 ( .A(n608), .B(KEYINPUT38), .ZN(n693) );
  XNOR2_X1 U376 ( .A(n764), .B(n371), .ZN(n443) );
  NAND2_X1 U377 ( .A1(n353), .A2(n410), .ZN(n409) );
  NAND2_X1 U378 ( .A1(n413), .A2(n414), .ZN(n353) );
  XNOR2_X2 U379 ( .A(n466), .B(n465), .ZN(n608) );
  AND2_X2 U380 ( .A1(n671), .A2(n672), .ZN(n673) );
  XNOR2_X1 U381 ( .A(n479), .B(KEYINPUT20), .ZN(n485) );
  NOR2_X2 U382 ( .A1(n608), .A2(n553), .ZN(n563) );
  NOR2_X2 U383 ( .A1(n368), .A2(n560), .ZN(n561) );
  XNOR2_X2 U384 ( .A(n502), .B(n501), .ZN(n649) );
  XNOR2_X1 U385 ( .A(n581), .B(n580), .ZN(n641) );
  INV_X1 U386 ( .A(n684), .ZN(n630) );
  NAND2_X1 U387 ( .A1(n357), .A2(n647), .ZN(n679) );
  NOR2_X1 U388 ( .A1(n670), .A2(n426), .ZN(n357) );
  XNOR2_X1 U389 ( .A(n366), .B(KEYINPUT40), .ZN(n405) );
  XNOR2_X1 U390 ( .A(n361), .B(n360), .ZN(n359) );
  OR2_X1 U391 ( .A1(n708), .A2(n632), .ZN(n361) );
  NOR2_X1 U392 ( .A1(n632), .A2(n688), .ZN(n631) );
  XNOR2_X1 U393 ( .A(n355), .B(n575), .ZN(n708) );
  XNOR2_X1 U394 ( .A(G140), .B(G137), .ZN(n539) );
  NOR2_X1 U395 ( .A1(n677), .A2(n676), .ZN(n408) );
  NAND2_X1 U396 ( .A1(n405), .A2(n388), .ZN(n387) );
  INV_X1 U397 ( .A(n367), .ZN(n716) );
  NAND2_X1 U398 ( .A1(n359), .A2(n579), .ZN(n581) );
  XNOR2_X1 U399 ( .A(n365), .B(KEYINPUT42), .ZN(n388) );
  NAND2_X1 U400 ( .A1(n717), .A2(n358), .ZN(n534) );
  NOR2_X1 U401 ( .A1(n574), .A2(n419), .ZN(n418) );
  XNOR2_X1 U402 ( .A(n552), .B(n551), .ZN(n368) );
  INV_X1 U403 ( .A(n628), .ZN(n354) );
  XNOR2_X1 U404 ( .A(n546), .B(G469), .ZN(n591) );
  XNOR2_X1 U405 ( .A(n540), .B(n539), .ZN(n764) );
  INV_X1 U406 ( .A(n644), .ZN(n362) );
  XNOR2_X1 U407 ( .A(n476), .B(G125), .ZN(n763) );
  INV_X1 U408 ( .A(KEYINPUT34), .ZN(n360) );
  NAND2_X1 U409 ( .A1(n630), .A2(n356), .ZN(n355) );
  NOR2_X1 U410 ( .A1(n571), .A2(n354), .ZN(n356) );
  AND2_X1 U411 ( .A1(n679), .A2(G472), .ZN(n389) );
  NAND2_X1 U412 ( .A1(n571), .A2(n619), .ZN(n611) );
  INV_X1 U413 ( .A(n571), .ZN(n358) );
  XNOR2_X1 U414 ( .A(n586), .B(KEYINPUT6), .ZN(n571) );
  NOR2_X1 U415 ( .A1(n670), .A2(KEYINPUT85), .ZN(n373) );
  NOR2_X1 U416 ( .A1(n670), .A2(n362), .ZN(n424) );
  AND2_X1 U417 ( .A1(n670), .A2(n363), .ZN(n675) );
  INV_X1 U418 ( .A(n674), .ZN(n363) );
  OR2_X1 U419 ( .A1(n670), .A2(G953), .ZN(n759) );
  XNOR2_X2 U420 ( .A(n436), .B(n364), .ZN(n670) );
  INV_X1 U421 ( .A(n375), .ZN(n364) );
  NAND2_X1 U422 ( .A1(n584), .A2(n583), .ZN(n366) );
  XNOR2_X2 U423 ( .A(n421), .B(KEYINPUT39), .ZN(n584) );
  OR2_X1 U424 ( .A1(n635), .A2(n368), .ZN(n367) );
  AND2_X1 U425 ( .A1(n648), .A2(n679), .ZN(n746) );
  XNOR2_X1 U426 ( .A(n387), .B(n404), .ZN(n369) );
  BUF_X1 U427 ( .A(n599), .Z(n370) );
  XNOR2_X1 U428 ( .A(n387), .B(n404), .ZN(n432) );
  BUF_X1 U429 ( .A(n554), .Z(n586) );
  XNOR2_X1 U430 ( .A(n504), .B(n503), .ZN(n554) );
  XOR2_X1 U431 ( .A(G472), .B(KEYINPUT75), .Z(n503) );
  NAND2_X1 U432 ( .A1(n649), .A2(n531), .ZN(n504) );
  XNOR2_X1 U433 ( .A(n384), .B(n453), .ZN(n456) );
  XOR2_X1 U434 ( .A(KEYINPUT80), .B(KEYINPUT18), .Z(n453) );
  NAND2_X1 U435 ( .A1(n765), .A2(G224), .ZN(n384) );
  AND2_X1 U436 ( .A1(n445), .A2(n610), .ZN(n444) );
  XNOR2_X1 U437 ( .A(n519), .B(n518), .ZN(n577) );
  XNOR2_X1 U438 ( .A(n517), .B(n516), .ZN(n518) );
  XOR2_X1 U439 ( .A(G110), .B(G107), .Z(n750) );
  AND2_X1 U440 ( .A1(n773), .A2(n724), .ZN(n622) );
  INV_X1 U441 ( .A(KEYINPUT76), .ZN(n399) );
  INV_X1 U442 ( .A(KEYINPUT46), .ZN(n404) );
  AND2_X1 U443 ( .A1(n622), .A2(KEYINPUT66), .ZN(n414) );
  INV_X1 U444 ( .A(n640), .ZN(n415) );
  XNOR2_X1 U445 ( .A(G113), .B(KEYINPUT3), .ZN(n461) );
  XNOR2_X1 U446 ( .A(G128), .B(KEYINPUT95), .ZN(n474) );
  NOR2_X1 U447 ( .A1(n493), .A2(n557), .ZN(n587) );
  INV_X1 U448 ( .A(n696), .ZN(n420) );
  XNOR2_X1 U449 ( .A(n440), .B(n569), .ZN(n574) );
  OR2_X1 U450 ( .A1(n577), .A2(n562), .ZN(n595) );
  XNOR2_X1 U451 ( .A(G137), .B(G146), .ZN(n499) );
  XNOR2_X1 U452 ( .A(n515), .B(n514), .ZN(n656) );
  XNOR2_X1 U453 ( .A(n513), .B(n512), .ZN(n514) );
  XOR2_X1 U454 ( .A(G140), .B(G131), .Z(n506) );
  XNOR2_X1 U455 ( .A(n463), .B(n752), .ZN(n663) );
  INV_X1 U456 ( .A(n553), .ZN(n692) );
  XNOR2_X1 U457 ( .A(n495), .B(n462), .ZN(n752) );
  XNOR2_X1 U458 ( .A(n505), .B(KEYINPUT16), .ZN(n462) );
  XNOR2_X1 U459 ( .A(n397), .B(n394), .ZN(n748) );
  XNOR2_X1 U460 ( .A(n396), .B(n395), .ZN(n394) );
  XNOR2_X1 U461 ( .A(n763), .B(n477), .ZN(n395) );
  NAND2_X1 U462 ( .A1(n423), .A2(KEYINPUT85), .ZN(n422) );
  NOR2_X1 U463 ( .A1(n725), .A2(n698), .ZN(n598) );
  NAND2_X1 U464 ( .A1(n447), .A2(n446), .ZN(n445) );
  INV_X1 U465 ( .A(KEYINPUT89), .ZN(n446) );
  INV_X1 U466 ( .A(n736), .ZN(n447) );
  AND2_X1 U467 ( .A1(n736), .A2(KEYINPUT89), .ZN(n448) );
  XOR2_X1 U468 ( .A(KEYINPUT77), .B(KEYINPUT5), .Z(n496) );
  NAND2_X1 U469 ( .A1(n412), .A2(n376), .ZN(n410) );
  XOR2_X1 U470 ( .A(KEYINPUT12), .B(KEYINPUT103), .Z(n510) );
  XNOR2_X1 U471 ( .A(G134), .B(G131), .ZN(n494) );
  XOR2_X1 U472 ( .A(G146), .B(G125), .Z(n454) );
  NAND2_X1 U473 ( .A1(G234), .A2(G237), .ZN(n488) );
  OR2_X1 U474 ( .A1(G237), .A2(G902), .ZN(n467) );
  NAND2_X1 U475 ( .A1(n554), .A2(n692), .ZN(n556) );
  XNOR2_X1 U476 ( .A(n461), .B(n460), .ZN(n438) );
  XNOR2_X1 U477 ( .A(n372), .B(n459), .ZN(n439) );
  INV_X1 U478 ( .A(KEYINPUT70), .ZN(n460) );
  XNOR2_X1 U479 ( .A(G122), .B(G104), .ZN(n505) );
  INV_X1 U480 ( .A(G953), .ZN(n755) );
  XNOR2_X1 U481 ( .A(KEYINPUT10), .B(G146), .ZN(n476) );
  XNOR2_X1 U482 ( .A(KEYINPUT97), .B(KEYINPUT23), .ZN(n477) );
  XNOR2_X1 U483 ( .A(n473), .B(n478), .ZN(n396) );
  XNOR2_X1 U484 ( .A(G119), .B(G110), .ZN(n472) );
  XNOR2_X1 U485 ( .A(G116), .B(G134), .ZN(n521) );
  XOR2_X1 U486 ( .A(G107), .B(G122), .Z(n522) );
  XNOR2_X1 U487 ( .A(KEYINPUT7), .B(KEYINPUT105), .ZN(n523) );
  XOR2_X1 U488 ( .A(KEYINPUT9), .B(KEYINPUT106), .Z(n524) );
  XNOR2_X1 U489 ( .A(G146), .B(G104), .ZN(n541) );
  XNOR2_X1 U490 ( .A(KEYINPUT72), .B(KEYINPUT73), .ZN(n451) );
  BUF_X1 U491 ( .A(n574), .Z(n632) );
  XNOR2_X1 U492 ( .A(n589), .B(n383), .ZN(n594) );
  XNOR2_X1 U493 ( .A(n588), .B(KEYINPUT28), .ZN(n383) );
  AND2_X1 U494 ( .A1(n587), .A2(n586), .ZN(n589) );
  INV_X1 U495 ( .A(KEYINPUT22), .ZN(n417) );
  INV_X1 U496 ( .A(KEYINPUT64), .ZN(n452) );
  XNOR2_X1 U497 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U498 ( .A(n663), .B(n662), .ZN(n664) );
  OR2_X1 U499 ( .A1(n765), .A2(G952), .ZN(n737) );
  XNOR2_X1 U500 ( .A(n602), .B(KEYINPUT110), .ZN(n774) );
  XNOR2_X1 U501 ( .A(n747), .B(n748), .ZN(n386) );
  NOR2_X1 U502 ( .A1(n391), .A2(n532), .ZN(n390) );
  XNOR2_X1 U503 ( .A(n742), .B(n741), .ZN(n385) );
  XOR2_X1 U504 ( .A(n545), .B(n544), .Z(n371) );
  XOR2_X1 U505 ( .A(G116), .B(G101), .Z(n372) );
  AND2_X1 U506 ( .A1(n643), .A2(n642), .ZN(n374) );
  INV_X1 U507 ( .A(G902), .ZN(n531) );
  XOR2_X1 U508 ( .A(KEYINPUT87), .B(KEYINPUT45), .Z(n375) );
  AND2_X1 U509 ( .A1(n621), .A2(KEYINPUT74), .ZN(n376) );
  INV_X1 U510 ( .A(n388), .ZN(n377) );
  XNOR2_X1 U511 ( .A(n469), .B(KEYINPUT83), .ZN(n470) );
  XOR2_X1 U512 ( .A(KEYINPUT8), .B(KEYINPUT69), .Z(n469) );
  XNOR2_X1 U513 ( .A(n400), .B(n399), .ZN(n398) );
  NOR2_X1 U514 ( .A1(n604), .A2(n434), .ZN(n433) );
  XNOR2_X1 U515 ( .A(n546), .B(G469), .ZN(n378) );
  NAND2_X1 U516 ( .A1(n443), .A2(n531), .ZN(n546) );
  NAND2_X1 U517 ( .A1(n420), .A2(n570), .ZN(n419) );
  AND2_X1 U518 ( .A1(n570), .A2(n550), .ZN(n628) );
  NAND2_X1 U519 ( .A1(n540), .A2(n495), .ZN(n381) );
  NAND2_X1 U520 ( .A1(n379), .A2(n380), .ZN(n382) );
  NAND2_X1 U521 ( .A1(n381), .A2(n382), .ZN(n502) );
  INV_X1 U522 ( .A(n540), .ZN(n379) );
  INV_X1 U523 ( .A(n495), .ZN(n380) );
  XNOR2_X1 U524 ( .A(n439), .B(n438), .ZN(n495) );
  XNOR2_X1 U525 ( .A(n418), .B(n417), .ZN(n616) );
  INV_X1 U526 ( .A(KEYINPUT48), .ZN(n434) );
  NOR2_X1 U527 ( .A1(n385), .A2(n749), .ZN(G54) );
  NOR2_X1 U528 ( .A1(n386), .A2(n749), .ZN(G66) );
  NAND2_X1 U529 ( .A1(n416), .A2(n415), .ZN(n413) );
  XNOR2_X2 U530 ( .A(n547), .B(KEYINPUT1), .ZN(n684) );
  NAND2_X1 U531 ( .A1(n648), .A2(n389), .ZN(n651) );
  NAND2_X1 U532 ( .A1(n648), .A2(n390), .ZN(n743) );
  INV_X1 U533 ( .A(n679), .ZN(n391) );
  NAND2_X1 U534 ( .A1(n648), .A2(n392), .ZN(n658) );
  AND2_X1 U535 ( .A1(n679), .A2(G475), .ZN(n392) );
  NAND2_X1 U536 ( .A1(n648), .A2(n393), .ZN(n665) );
  AND2_X1 U537 ( .A1(n679), .A2(G210), .ZN(n393) );
  NOR2_X1 U538 ( .A1(n748), .A2(G902), .ZN(n484) );
  AND2_X1 U539 ( .A1(n527), .A2(G221), .ZN(n397) );
  INV_X1 U540 ( .A(n405), .ZN(n654) );
  NAND2_X1 U541 ( .A1(n398), .A2(n603), .ZN(n604) );
  NAND2_X1 U542 ( .A1(n401), .A2(n774), .ZN(n400) );
  XNOR2_X1 U543 ( .A(n598), .B(KEYINPUT47), .ZN(n401) );
  NAND2_X1 U544 ( .A1(n402), .A2(n644), .ZN(n425) );
  NAND2_X1 U545 ( .A1(n403), .A2(n426), .ZN(n402) );
  NAND2_X1 U546 ( .A1(n671), .A2(n373), .ZN(n403) );
  XNOR2_X2 U547 ( .A(n646), .B(KEYINPUT86), .ZN(n671) );
  NAND2_X1 U548 ( .A1(n406), .A2(n713), .ZN(n715) );
  NAND2_X1 U549 ( .A1(n407), .A2(n679), .ZN(n406) );
  XNOR2_X1 U550 ( .A(n408), .B(n678), .ZN(n407) );
  NAND2_X1 U551 ( .A1(n409), .A2(n374), .ZN(n436) );
  INV_X1 U552 ( .A(n622), .ZN(n412) );
  INV_X1 U553 ( .A(n641), .ZN(n416) );
  INV_X1 U554 ( .A(n584), .ZN(n582) );
  NAND2_X1 U555 ( .A1(n599), .A2(n693), .ZN(n421) );
  XNOR2_X1 U556 ( .A(n561), .B(KEYINPUT78), .ZN(n599) );
  NAND2_X2 U557 ( .A1(n425), .A2(n422), .ZN(n648) );
  NAND2_X1 U558 ( .A1(n671), .A2(n424), .ZN(n423) );
  INV_X1 U559 ( .A(KEYINPUT2), .ZN(n426) );
  NAND2_X1 U560 ( .A1(n429), .A2(n428), .ZN(n450) );
  XNOR2_X2 U561 ( .A(n427), .B(n494), .ZN(n540) );
  XNOR2_X1 U562 ( .A(n427), .B(n545), .ZN(n458) );
  XNOR2_X2 U563 ( .A(n520), .B(KEYINPUT4), .ZN(n427) );
  NAND2_X1 U564 ( .A1(n369), .A2(n433), .ZN(n428) );
  NAND2_X1 U565 ( .A1(n430), .A2(n434), .ZN(n429) );
  NAND2_X1 U566 ( .A1(n432), .A2(n431), .ZN(n430) );
  INV_X1 U567 ( .A(n604), .ZN(n431) );
  NAND2_X1 U568 ( .A1(n450), .A2(n448), .ZN(n435) );
  NAND2_X1 U569 ( .A1(n435), .A2(n444), .ZN(n437) );
  NOR2_X2 U570 ( .A1(n437), .A2(n449), .ZN(n646) );
  NAND2_X1 U571 ( .A1(n592), .A2(n568), .ZN(n440) );
  XNOR2_X1 U572 ( .A(n563), .B(n441), .ZN(n592) );
  INV_X1 U573 ( .A(KEYINPUT19), .ZN(n441) );
  XNOR2_X2 U574 ( .A(n442), .B(G143), .ZN(n520) );
  XNOR2_X2 U575 ( .A(G128), .B(KEYINPUT65), .ZN(n442) );
  XNOR2_X1 U576 ( .A(n443), .B(n740), .ZN(n741) );
  NOR2_X1 U577 ( .A1(n450), .A2(KEYINPUT89), .ZN(n449) );
  INV_X1 U578 ( .A(n550), .ZN(n619) );
  INV_X1 U579 ( .A(KEYINPUT30), .ZN(n555) );
  INV_X1 U580 ( .A(KEYINPUT81), .ZN(n678) );
  XNOR2_X1 U581 ( .A(n750), .B(n451), .ZN(n545) );
  XNOR2_X2 U582 ( .A(n452), .B(G953), .ZN(n765) );
  XOR2_X1 U583 ( .A(KEYINPUT17), .B(n454), .Z(n455) );
  XNOR2_X1 U584 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U585 ( .A(n458), .B(n457), .ZN(n463) );
  XNOR2_X1 U586 ( .A(KEYINPUT71), .B(G119), .ZN(n459) );
  XNOR2_X1 U587 ( .A(G902), .B(KEYINPUT92), .ZN(n464) );
  XNOR2_X1 U588 ( .A(n464), .B(KEYINPUT15), .ZN(n645) );
  NAND2_X1 U589 ( .A1(n663), .A2(n645), .ZN(n466) );
  NAND2_X1 U590 ( .A1(G210), .A2(n467), .ZN(n465) );
  NAND2_X1 U591 ( .A1(G214), .A2(n467), .ZN(n468) );
  XNOR2_X1 U592 ( .A(KEYINPUT93), .B(n468), .ZN(n553) );
  NAND2_X1 U593 ( .A1(G234), .A2(n765), .ZN(n471) );
  XNOR2_X1 U594 ( .A(n471), .B(n470), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n472), .B(n539), .ZN(n473) );
  XOR2_X1 U596 ( .A(KEYINPUT96), .B(KEYINPUT24), .Z(n475) );
  XNOR2_X1 U597 ( .A(n475), .B(n474), .ZN(n478) );
  XOR2_X1 U598 ( .A(KEYINPUT98), .B(KEYINPUT79), .Z(n481) );
  NAND2_X1 U599 ( .A1(G234), .A2(n645), .ZN(n479) );
  NAND2_X1 U600 ( .A1(n485), .A2(G217), .ZN(n480) );
  XNOR2_X1 U601 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U602 ( .A(KEYINPUT25), .B(n482), .ZN(n483) );
  XNOR2_X1 U603 ( .A(n484), .B(n483), .ZN(n550) );
  XOR2_X1 U604 ( .A(KEYINPUT99), .B(KEYINPUT21), .Z(n487) );
  NAND2_X1 U605 ( .A1(n485), .A2(G221), .ZN(n486) );
  XOR2_X1 U606 ( .A(n487), .B(n486), .Z(n681) );
  NAND2_X1 U607 ( .A1(n619), .A2(n681), .ZN(n493) );
  XNOR2_X1 U608 ( .A(n488), .B(KEYINPUT14), .ZN(n491) );
  NAND2_X1 U609 ( .A1(n491), .A2(G902), .ZN(n489) );
  XOR2_X1 U610 ( .A(KEYINPUT94), .B(n489), .Z(n564) );
  NOR2_X1 U611 ( .A1(n765), .A2(G900), .ZN(n490) );
  AND2_X1 U612 ( .A1(n564), .A2(n490), .ZN(n492) );
  AND2_X1 U613 ( .A1(G952), .A2(n491), .ZN(n705) );
  AND2_X1 U614 ( .A1(n705), .A2(n755), .ZN(n565) );
  NOR2_X1 U615 ( .A1(n492), .A2(n565), .ZN(n557) );
  INV_X1 U616 ( .A(n587), .ZN(n535) );
  NOR2_X1 U617 ( .A1(G953), .A2(G237), .ZN(n508) );
  NAND2_X1 U618 ( .A1(n508), .A2(G210), .ZN(n497) );
  XNOR2_X1 U619 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U620 ( .A(n498), .B(KEYINPUT102), .Z(n500) );
  XNOR2_X1 U621 ( .A(n500), .B(n499), .ZN(n501) );
  XOR2_X1 U622 ( .A(n505), .B(n763), .Z(n507) );
  XNOR2_X1 U623 ( .A(n507), .B(n506), .ZN(n515) );
  NAND2_X1 U624 ( .A1(G214), .A2(n508), .ZN(n509) );
  XNOR2_X1 U625 ( .A(n510), .B(n509), .ZN(n511) );
  XOR2_X1 U626 ( .A(n511), .B(KEYINPUT11), .Z(n513) );
  XNOR2_X1 U627 ( .A(G113), .B(G143), .ZN(n512) );
  NOR2_X1 U628 ( .A1(G902), .A2(n656), .ZN(n519) );
  XNOR2_X1 U629 ( .A(KEYINPUT104), .B(KEYINPUT13), .ZN(n517) );
  INV_X1 U630 ( .A(G475), .ZN(n516) );
  XNOR2_X1 U631 ( .A(n522), .B(n521), .ZN(n526) );
  XNOR2_X1 U632 ( .A(n524), .B(n523), .ZN(n525) );
  XOR2_X1 U633 ( .A(n526), .B(n525), .Z(n529) );
  NAND2_X1 U634 ( .A1(G217), .A2(n527), .ZN(n528) );
  XNOR2_X1 U635 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U636 ( .A(n520), .B(n530), .ZN(n744) );
  NAND2_X1 U637 ( .A1(n744), .A2(n531), .ZN(n533) );
  INV_X1 U638 ( .A(G478), .ZN(n532) );
  XNOR2_X1 U639 ( .A(n533), .B(n532), .ZN(n576) );
  INV_X1 U640 ( .A(n576), .ZN(n562) );
  XNOR2_X1 U641 ( .A(n595), .B(KEYINPUT109), .ZN(n717) );
  NOR2_X1 U642 ( .A1(n535), .A2(n534), .ZN(n605) );
  NAND2_X1 U643 ( .A1(n563), .A2(n605), .ZN(n538) );
  XNOR2_X1 U644 ( .A(KEYINPUT91), .B(KEYINPUT112), .ZN(n536) );
  XNOR2_X1 U645 ( .A(n536), .B(KEYINPUT36), .ZN(n537) );
  XNOR2_X1 U646 ( .A(n538), .B(n537), .ZN(n548) );
  NAND2_X1 U647 ( .A1(n765), .A2(G227), .ZN(n543) );
  XNOR2_X1 U648 ( .A(n541), .B(G101), .ZN(n542) );
  XNOR2_X1 U649 ( .A(n543), .B(n542), .ZN(n544) );
  INV_X1 U650 ( .A(n378), .ZN(n547) );
  NAND2_X1 U651 ( .A1(n548), .A2(n630), .ZN(n603) );
  XOR2_X1 U652 ( .A(G125), .B(KEYINPUT37), .Z(n549) );
  XNOR2_X1 U653 ( .A(n603), .B(n549), .ZN(G27) );
  XNOR2_X1 U654 ( .A(n681), .B(KEYINPUT100), .ZN(n570) );
  NAND2_X1 U655 ( .A1(n591), .A2(n628), .ZN(n552) );
  INV_X1 U656 ( .A(KEYINPUT101), .ZN(n551) );
  XNOR2_X1 U657 ( .A(n556), .B(n555), .ZN(n559) );
  INV_X1 U658 ( .A(n557), .ZN(n558) );
  NAND2_X1 U659 ( .A1(n559), .A2(n558), .ZN(n560) );
  AND2_X1 U660 ( .A1(n562), .A2(n577), .ZN(n596) );
  INV_X1 U661 ( .A(n596), .ZN(n734) );
  OR2_X1 U662 ( .A1(n582), .A2(n734), .ZN(n610) );
  XNOR2_X1 U663 ( .A(n610), .B(G134), .ZN(G36) );
  NAND2_X1 U664 ( .A1(n577), .A2(n576), .ZN(n696) );
  NOR2_X1 U665 ( .A1(G898), .A2(n755), .ZN(n753) );
  NAND2_X1 U666 ( .A1(n564), .A2(n753), .ZN(n567) );
  INV_X1 U667 ( .A(n565), .ZN(n566) );
  NAND2_X1 U668 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U669 ( .A(KEYINPUT68), .B(KEYINPUT0), .ZN(n569) );
  INV_X1 U670 ( .A(n616), .ZN(n613) );
  INV_X1 U671 ( .A(n619), .ZN(n680) );
  NAND2_X1 U672 ( .A1(n571), .A2(n680), .ZN(n572) );
  NOR2_X1 U673 ( .A1(n572), .A2(n630), .ZN(n573) );
  NAND2_X1 U674 ( .A1(n613), .A2(n573), .ZN(n627) );
  XNOR2_X1 U675 ( .A(n627), .B(G101), .ZN(G3) );
  INV_X1 U676 ( .A(KEYINPUT33), .ZN(n575) );
  OR2_X1 U677 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U678 ( .A(n578), .B(KEYINPUT108), .ZN(n600) );
  INV_X1 U679 ( .A(n600), .ZN(n579) );
  XNOR2_X1 U680 ( .A(KEYINPUT88), .B(KEYINPUT35), .ZN(n580) );
  XOR2_X1 U681 ( .A(n641), .B(G122), .Z(G24) );
  INV_X1 U682 ( .A(n595), .ZN(n583) );
  NAND2_X1 U683 ( .A1(n693), .A2(n692), .ZN(n697) );
  XNOR2_X1 U684 ( .A(n585), .B(KEYINPUT41), .ZN(n709) );
  INV_X1 U685 ( .A(KEYINPUT111), .ZN(n588) );
  NAND2_X1 U686 ( .A1(n594), .A2(n378), .ZN(n590) );
  AND2_X1 U687 ( .A1(n378), .A2(n592), .ZN(n593) );
  NAND2_X1 U688 ( .A1(n594), .A2(n593), .ZN(n725) );
  NOR2_X1 U689 ( .A1(n583), .A2(n596), .ZN(n597) );
  XOR2_X1 U690 ( .A(n597), .B(KEYINPUT107), .Z(n698) );
  NOR2_X1 U691 ( .A1(n600), .A2(n608), .ZN(n601) );
  NAND2_X1 U692 ( .A1(n370), .A2(n601), .ZN(n602) );
  AND2_X1 U693 ( .A1(n605), .A2(n692), .ZN(n606) );
  NAND2_X1 U694 ( .A1(n606), .A2(n684), .ZN(n607) );
  XNOR2_X1 U695 ( .A(n607), .B(KEYINPUT43), .ZN(n609) );
  NAND2_X1 U696 ( .A1(n609), .A2(n608), .ZN(n736) );
  NOR2_X1 U697 ( .A1(n611), .A2(n684), .ZN(n612) );
  NAND2_X1 U698 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U699 ( .A(n614), .B(KEYINPUT32), .ZN(n773) );
  INV_X1 U700 ( .A(n586), .ZN(n633) );
  NAND2_X1 U701 ( .A1(n684), .A2(n633), .ZN(n615) );
  NOR2_X1 U702 ( .A1(n616), .A2(n615), .ZN(n618) );
  INV_X1 U703 ( .A(KEYINPUT67), .ZN(n617) );
  XNOR2_X1 U704 ( .A(n618), .B(n617), .ZN(n620) );
  NAND2_X1 U705 ( .A1(n620), .A2(n619), .ZN(n724) );
  INV_X1 U706 ( .A(KEYINPUT44), .ZN(n623) );
  NAND2_X1 U707 ( .A1(n623), .A2(KEYINPUT74), .ZN(n640) );
  NAND2_X1 U708 ( .A1(KEYINPUT66), .A2(KEYINPUT44), .ZN(n621) );
  NAND2_X1 U709 ( .A1(n623), .A2(KEYINPUT66), .ZN(n625) );
  NAND2_X1 U710 ( .A1(KEYINPUT74), .A2(KEYINPUT44), .ZN(n624) );
  NAND2_X1 U711 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U712 ( .A1(n627), .A2(n626), .ZN(n639) );
  NOR2_X1 U713 ( .A1(n633), .A2(n354), .ZN(n629) );
  NAND2_X1 U714 ( .A1(n630), .A2(n629), .ZN(n688) );
  XNOR2_X1 U715 ( .A(n631), .B(KEYINPUT31), .ZN(n733) );
  INV_X1 U716 ( .A(n733), .ZN(n636) );
  INV_X1 U717 ( .A(n632), .ZN(n634) );
  NAND2_X1 U718 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U719 ( .A1(n636), .A2(n716), .ZN(n637) );
  NOR2_X1 U720 ( .A1(n637), .A2(n698), .ZN(n638) );
  NOR2_X1 U721 ( .A1(n639), .A2(n638), .ZN(n643) );
  NAND2_X1 U722 ( .A1(n641), .A2(n640), .ZN(n642) );
  INV_X1 U723 ( .A(n645), .ZN(n644) );
  BUF_X1 U724 ( .A(n646), .Z(n647) );
  XNOR2_X1 U725 ( .A(n649), .B(KEYINPUT62), .ZN(n650) );
  XNOR2_X1 U726 ( .A(n651), .B(n650), .ZN(n652) );
  NAND2_X1 U727 ( .A1(n652), .A2(n737), .ZN(n653) );
  XNOR2_X1 U728 ( .A(n653), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U729 ( .A(n654), .B(G131), .Z(G33) );
  XOR2_X1 U730 ( .A(KEYINPUT123), .B(KEYINPUT59), .Z(n655) );
  XNOR2_X1 U731 ( .A(n658), .B(n657), .ZN(n659) );
  NAND2_X1 U732 ( .A1(n659), .A2(n737), .ZN(n661) );
  XOR2_X1 U733 ( .A(KEYINPUT124), .B(KEYINPUT60), .Z(n660) );
  XNOR2_X1 U734 ( .A(n661), .B(n660), .ZN(G60) );
  XOR2_X1 U735 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n662) );
  XNOR2_X1 U736 ( .A(n665), .B(n664), .ZN(n666) );
  NAND2_X1 U737 ( .A1(n666), .A2(n737), .ZN(n669) );
  XNOR2_X1 U738 ( .A(KEYINPUT120), .B(KEYINPUT56), .ZN(n667) );
  XOR2_X1 U739 ( .A(n667), .B(KEYINPUT90), .Z(n668) );
  XNOR2_X1 U740 ( .A(n669), .B(n668), .ZN(G51) );
  NAND2_X1 U741 ( .A1(n670), .A2(KEYINPUT84), .ZN(n672) );
  XNOR2_X1 U742 ( .A(KEYINPUT2), .B(KEYINPUT82), .ZN(n674) );
  NOR2_X1 U743 ( .A1(n673), .A2(n674), .ZN(n677) );
  NOR2_X1 U744 ( .A1(n675), .A2(KEYINPUT84), .ZN(n676) );
  NOR2_X1 U745 ( .A1(n681), .A2(n680), .ZN(n682) );
  XOR2_X1 U746 ( .A(KEYINPUT49), .B(n682), .Z(n683) );
  NOR2_X1 U747 ( .A1(n586), .A2(n683), .ZN(n687) );
  NAND2_X1 U748 ( .A1(n684), .A2(n354), .ZN(n685) );
  XNOR2_X1 U749 ( .A(n685), .B(KEYINPUT50), .ZN(n686) );
  NAND2_X1 U750 ( .A1(n687), .A2(n686), .ZN(n689) );
  NAND2_X1 U751 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U752 ( .A(KEYINPUT51), .B(n690), .ZN(n691) );
  NOR2_X1 U753 ( .A1(n691), .A2(n709), .ZN(n703) );
  NOR2_X1 U754 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U755 ( .A(KEYINPUT117), .B(n694), .Z(n695) );
  NOR2_X1 U756 ( .A1(n696), .A2(n695), .ZN(n700) );
  NOR2_X1 U757 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U758 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U759 ( .A1(n701), .A2(n708), .ZN(n702) );
  NOR2_X1 U760 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U761 ( .A(KEYINPUT52), .B(n704), .Z(n706) );
  NAND2_X1 U762 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U763 ( .A(n707), .B(KEYINPUT118), .ZN(n712) );
  NOR2_X1 U764 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U765 ( .A1(n710), .A2(G953), .ZN(n711) );
  AND2_X1 U766 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U767 ( .A(KEYINPUT119), .B(KEYINPUT53), .ZN(n714) );
  XNOR2_X1 U768 ( .A(n715), .B(n714), .ZN(G75) );
  INV_X1 U769 ( .A(n717), .ZN(n731) );
  NOR2_X1 U770 ( .A1(n367), .A2(n731), .ZN(n719) );
  XNOR2_X1 U771 ( .A(G104), .B(KEYINPUT113), .ZN(n718) );
  XNOR2_X1 U772 ( .A(n719), .B(n718), .ZN(G6) );
  XOR2_X1 U773 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n721) );
  XNOR2_X1 U774 ( .A(G107), .B(KEYINPUT114), .ZN(n720) );
  XNOR2_X1 U775 ( .A(n721), .B(n720), .ZN(n723) );
  NOR2_X1 U776 ( .A1(n367), .A2(n734), .ZN(n722) );
  XOR2_X1 U777 ( .A(n723), .B(n722), .Z(G9) );
  XNOR2_X1 U778 ( .A(G110), .B(n724), .ZN(G12) );
  NOR2_X1 U779 ( .A1(n734), .A2(n725), .ZN(n727) );
  XNOR2_X1 U780 ( .A(G128), .B(KEYINPUT29), .ZN(n726) );
  XNOR2_X1 U781 ( .A(n727), .B(n726), .ZN(G30) );
  NOR2_X1 U782 ( .A1(n731), .A2(n725), .ZN(n729) );
  XNOR2_X1 U783 ( .A(KEYINPUT115), .B(KEYINPUT116), .ZN(n728) );
  XNOR2_X1 U784 ( .A(n729), .B(n728), .ZN(n730) );
  XNOR2_X1 U785 ( .A(G146), .B(n730), .ZN(G48) );
  NOR2_X1 U786 ( .A1(n731), .A2(n733), .ZN(n732) );
  XOR2_X1 U787 ( .A(G113), .B(n732), .Z(G15) );
  NOR2_X1 U788 ( .A1(n734), .A2(n733), .ZN(n735) );
  XOR2_X1 U789 ( .A(G116), .B(n735), .Z(G18) );
  XNOR2_X1 U790 ( .A(G140), .B(n736), .ZN(G42) );
  INV_X1 U791 ( .A(n737), .ZN(n749) );
  NAND2_X1 U792 ( .A1(n746), .A2(G469), .ZN(n742) );
  XOR2_X1 U793 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(n739) );
  XNOR2_X1 U794 ( .A(KEYINPUT122), .B(KEYINPUT121), .ZN(n738) );
  XNOR2_X1 U795 ( .A(n739), .B(n738), .ZN(n740) );
  XOR2_X1 U796 ( .A(n744), .B(n743), .Z(n745) );
  NOR2_X1 U797 ( .A1(n749), .A2(n745), .ZN(G63) );
  NAND2_X1 U798 ( .A1(n746), .A2(G217), .ZN(n747) );
  XOR2_X1 U799 ( .A(n750), .B(KEYINPUT125), .Z(n751) );
  XNOR2_X1 U800 ( .A(n752), .B(n751), .ZN(n754) );
  NOR2_X1 U801 ( .A1(n754), .A2(n753), .ZN(n762) );
  NAND2_X1 U802 ( .A1(G953), .A2(G224), .ZN(n756) );
  XNOR2_X1 U803 ( .A(KEYINPUT61), .B(n756), .ZN(n757) );
  NAND2_X1 U804 ( .A1(n757), .A2(G898), .ZN(n758) );
  NAND2_X1 U805 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U806 ( .A(n760), .B(KEYINPUT126), .ZN(n761) );
  XNOR2_X1 U807 ( .A(n762), .B(n761), .ZN(G69) );
  XOR2_X1 U808 ( .A(n764), .B(n763), .Z(n767) );
  XNOR2_X1 U809 ( .A(n671), .B(n767), .ZN(n766) );
  NAND2_X1 U810 ( .A1(n766), .A2(n765), .ZN(n771) );
  XOR2_X1 U811 ( .A(G227), .B(n767), .Z(n768) );
  NAND2_X1 U812 ( .A1(n768), .A2(G900), .ZN(n769) );
  NAND2_X1 U813 ( .A1(n769), .A2(G953), .ZN(n770) );
  NAND2_X1 U814 ( .A1(n771), .A2(n770), .ZN(n772) );
  XOR2_X1 U815 ( .A(KEYINPUT127), .B(n772), .Z(G72) );
  XNOR2_X1 U816 ( .A(G119), .B(n773), .ZN(G21) );
  XNOR2_X1 U817 ( .A(G143), .B(n774), .ZN(G45) );
  XOR2_X1 U818 ( .A(n377), .B(G137), .Z(G39) );
endmodule

