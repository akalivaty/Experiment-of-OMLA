//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 1 1 1 0 0 0 1 0 1 0 1 1 0 1 1 1 1 1 0 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 1 1 0 1 1 1 1 0 1 0 1 0 1 0 0 1 1 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n803, new_n804, new_n805, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n853,
    new_n854, new_n855, new_n857, new_n858, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n871, new_n872, new_n874, new_n875, new_n876, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n909, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT31), .B(G50gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  OR2_X1    g003(.A1(new_n204), .A2(KEYINPUT81), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(KEYINPUT81), .ZN(new_n206));
  XOR2_X1   g005(.A(G155gat), .B(G162gat), .Z(new_n207));
  XNOR2_X1  g006(.A(G141gat), .B(G148gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n207), .B1(KEYINPUT2), .B2(new_n208), .ZN(new_n209));
  XOR2_X1   g008(.A(G141gat), .B(G148gat), .Z(new_n210));
  XNOR2_X1  g009(.A(G155gat), .B(G162gat), .ZN(new_n211));
  INV_X1    g010(.A(G155gat), .ZN(new_n212));
  INV_X1    g011(.A(G162gat), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT2), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n210), .A2(new_n211), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n209), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G197gat), .B(G204gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT22), .ZN(new_n218));
  INV_X1    g017(.A(G211gat), .ZN(new_n219));
  INV_X1    g018(.A(G218gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n217), .A2(new_n221), .ZN(new_n222));
  XOR2_X1   g021(.A(G211gat), .B(G218gat), .Z(new_n223));
  XNOR2_X1  g022(.A(new_n222), .B(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT29), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT80), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n226), .B(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n216), .B1(new_n228), .B2(KEYINPUT3), .ZN(new_n229));
  NAND2_X1  g028(.A1(G228gat), .A2(G233gat), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n216), .A2(KEYINPUT3), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n231), .B(KEYINPUT74), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n232), .A2(new_n225), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n229), .B(new_n230), .C1(new_n224), .C2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(G22gat), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n224), .B1(new_n232), .B2(new_n225), .ZN(new_n236));
  INV_X1    g035(.A(new_n216), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n237), .B1(new_n226), .B2(new_n238), .ZN(new_n239));
  OAI211_X1 g038(.A(G228gat), .B(G233gat), .C1(new_n236), .C2(new_n239), .ZN(new_n240));
  AND3_X1   g039(.A1(new_n234), .A2(new_n235), .A3(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n235), .B1(new_n234), .B2(new_n240), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n205), .B(new_n206), .C1(new_n241), .C2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n234), .A2(new_n240), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(G22gat), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n234), .A2(new_n235), .A3(new_n240), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n245), .A2(KEYINPUT81), .A3(new_n246), .A4(new_n204), .ZN(new_n247));
  AND2_X1   g046(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(G113gat), .B(G120gat), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n249), .A2(KEYINPUT1), .ZN(new_n250));
  XNOR2_X1  g049(.A(G127gat), .B(G134gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n251), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n253), .B1(KEYINPUT1), .B2(new_n249), .ZN(new_n254));
  AND2_X1   g053(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n255), .B1(KEYINPUT3), .B2(new_n216), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n232), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n255), .A2(new_n237), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(KEYINPUT4), .ZN(new_n259));
  NAND2_X1  g058(.A1(G225gat), .A2(G233gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n260), .B(KEYINPUT75), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n257), .A2(new_n259), .A3(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(KEYINPUT77), .B(KEYINPUT5), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT76), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n263), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(G1gat), .B(G29gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n269), .B(KEYINPUT0), .ZN(new_n270));
  XNOR2_X1  g069(.A(G57gat), .B(G85gat), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n270), .B(new_n271), .Z(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n257), .A2(new_n259), .A3(new_n262), .A4(new_n266), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n255), .B(new_n216), .ZN(new_n275));
  OR3_X1    g074(.A1(new_n275), .A2(new_n262), .A3(new_n264), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n268), .A2(new_n273), .A3(new_n274), .A4(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT6), .ZN(new_n278));
  OR2_X1    g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n274), .A2(new_n276), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n273), .B1(new_n281), .B2(new_n268), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n277), .A2(new_n278), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n279), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT35), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n248), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT71), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT67), .ZN(new_n288));
  NOR2_X1   g087(.A1(G169gat), .A2(G176gat), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT23), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n289), .B(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(G169gat), .A2(G176gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n292), .B(KEYINPUT64), .ZN(new_n293));
  AND2_X1   g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  AND2_X1   g093(.A1(new_n294), .A2(KEYINPUT25), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT65), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n296), .B(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n299));
  XOR2_X1   g098(.A(KEYINPUT66), .B(G183gat), .Z(new_n300));
  OAI211_X1 g099(.A(new_n298), .B(new_n299), .C1(G190gat), .C2(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n288), .B1(new_n295), .B2(new_n301), .ZN(new_n302));
  NAND4_X1  g101(.A1(new_n301), .A2(new_n288), .A3(KEYINPUT25), .A4(new_n294), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n299), .B1(G183gat), .B2(G190gat), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n291), .B(new_n293), .C1(new_n296), .C2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT25), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  OR2_X1    g107(.A1(new_n302), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT27), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(G183gat), .ZN(new_n311));
  XOR2_X1   g110(.A(new_n311), .B(KEYINPUT68), .Z(new_n312));
  NOR2_X1   g111(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n313));
  OAI211_X1 g112(.A(new_n312), .B(new_n313), .C1(new_n310), .C2(new_n300), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n289), .B(KEYINPUT26), .ZN(new_n315));
  AOI22_X1  g114(.A1(new_n315), .A2(new_n293), .B1(G183gat), .B2(G190gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(KEYINPUT27), .B(G183gat), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT69), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n317), .B(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(G190gat), .ZN(new_n320));
  AND2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT28), .ZN(new_n322));
  OAI211_X1 g121(.A(new_n314), .B(new_n316), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n309), .A2(KEYINPUT70), .A3(new_n255), .A4(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(G227gat), .A2(G233gat), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT70), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n323), .B1(new_n302), .B2(new_n308), .ZN(new_n327));
  INV_X1    g126(.A(new_n255), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n255), .B(new_n323), .C1(new_n302), .C2(new_n308), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n324), .B(new_n325), .C1(new_n329), .C2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT34), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n287), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n332), .A2(KEYINPUT71), .A3(KEYINPUT34), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n330), .A2(new_n326), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n327), .A2(new_n328), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(KEYINPUT70), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n337), .B1(new_n339), .B2(new_n330), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n340), .A2(new_n334), .A3(new_n325), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n335), .A2(new_n336), .A3(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n324), .B1(new_n329), .B2(new_n331), .ZN(new_n343));
  INV_X1    g142(.A(new_n325), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT33), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT32), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n346), .B1(new_n343), .B2(new_n344), .ZN(new_n347));
  XOR2_X1   g146(.A(G15gat), .B(G43gat), .Z(new_n348));
  XNOR2_X1  g147(.A(G71gat), .B(G99gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n348), .B(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NOR3_X1   g150(.A1(new_n345), .A2(new_n347), .A3(new_n351), .ZN(new_n352));
  AOI221_X4 g151(.A(new_n346), .B1(KEYINPUT33), .B2(new_n350), .C1(new_n343), .C2(new_n344), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n342), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n343), .A2(new_n344), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT32), .ZN(new_n356));
  INV_X1    g155(.A(new_n355), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n356), .B(new_n350), .C1(new_n357), .C2(KEYINPUT33), .ZN(new_n358));
  AND2_X1   g157(.A1(new_n341), .A2(new_n336), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n347), .B1(new_n345), .B2(new_n351), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n358), .A2(new_n359), .A3(new_n335), .A4(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n354), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(G226gat), .A2(G233gat), .ZN(new_n363));
  XOR2_X1   g162(.A(new_n363), .B(KEYINPUT72), .Z(new_n364));
  AOI21_X1  g163(.A(new_n364), .B1(new_n327), .B2(new_n225), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n327), .A2(new_n364), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT73), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT73), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n327), .A2(new_n369), .A3(new_n364), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n366), .A2(new_n368), .A3(new_n224), .A4(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n224), .ZN(new_n372));
  INV_X1    g171(.A(new_n367), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n372), .B1(new_n373), .B2(new_n365), .ZN(new_n374));
  AND2_X1   g173(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT30), .ZN(new_n376));
  XNOR2_X1  g175(.A(G8gat), .B(G36gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(G64gat), .B(G92gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n377), .B(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n375), .A2(new_n376), .A3(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n371), .A2(new_n374), .A3(new_n380), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT30), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n380), .B1(new_n371), .B2(new_n374), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n381), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NOR3_X1   g185(.A1(new_n286), .A2(new_n362), .A3(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n354), .A2(new_n361), .A3(new_n248), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(KEYINPUT83), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT78), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n390), .B1(new_n283), .B2(new_n282), .ZN(new_n391));
  INV_X1    g190(.A(new_n268), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n272), .B1(new_n392), .B2(new_n280), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n393), .A2(KEYINPUT78), .A3(new_n277), .A4(new_n278), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n391), .A2(new_n394), .A3(new_n279), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT79), .B1(new_n395), .B2(new_n385), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n395), .A2(new_n385), .A3(KEYINPUT79), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT83), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n354), .A2(new_n361), .A3(new_n248), .A4(new_n399), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n389), .A2(new_n397), .A3(new_n398), .A4(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n387), .B1(new_n401), .B2(KEYINPUT35), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n243), .A2(new_n247), .ZN(new_n403));
  AND3_X1   g202(.A1(new_n395), .A2(new_n385), .A3(KEYINPUT79), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n403), .B1(new_n404), .B2(new_n396), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n284), .B1(new_n375), .B2(new_n380), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT37), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n380), .B1(new_n375), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n371), .A2(new_n374), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT37), .ZN(new_n410));
  AND3_X1   g209(.A1(new_n408), .A2(KEYINPUT38), .A3(new_n410), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n373), .A2(new_n365), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT82), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n412), .A2(new_n413), .A3(new_n224), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n366), .A2(new_n368), .A3(new_n370), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n414), .B1(new_n415), .B2(new_n224), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n413), .B1(new_n412), .B2(new_n224), .ZN(new_n417));
  OAI21_X1  g216(.A(KEYINPUT37), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT38), .B1(new_n418), .B2(new_n408), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n406), .B1(new_n411), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT40), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n262), .B1(new_n257), .B2(new_n259), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n275), .A2(new_n262), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT39), .ZN(new_n424));
  OR2_X1    g223(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(new_n272), .ZN(new_n426));
  INV_X1    g225(.A(new_n422), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n427), .A2(KEYINPUT39), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n421), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(new_n277), .ZN(new_n430));
  NOR3_X1   g229(.A1(new_n426), .A2(new_n421), .A3(new_n428), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n403), .B1(new_n386), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n420), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT36), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n362), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n354), .A2(new_n361), .A3(KEYINPUT36), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AND3_X1   g237(.A1(new_n405), .A2(new_n434), .A3(new_n438), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n402), .A2(new_n439), .ZN(new_n440));
  OR2_X1    g239(.A1(G57gat), .A2(G64gat), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT93), .ZN(new_n442));
  NAND2_X1  g241(.A1(G57gat), .A2(G64gat), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  AND2_X1   g243(.A1(G57gat), .A2(G64gat), .ZN(new_n445));
  NOR2_X1   g244(.A1(G57gat), .A2(G64gat), .ZN(new_n446));
  OAI21_X1  g245(.A(KEYINPUT93), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OR2_X1    g246(.A1(G71gat), .A2(G78gat), .ZN(new_n448));
  NAND2_X1  g247(.A1(G71gat), .A2(G78gat), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n444), .A2(new_n447), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n452), .B(KEYINPUT92), .ZN(new_n453));
  OAI21_X1  g252(.A(KEYINPUT94), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n445), .A2(new_n446), .ZN(new_n455));
  AOI22_X1  g254(.A1(new_n455), .A2(new_n442), .B1(new_n449), .B2(new_n448), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT94), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT9), .ZN(new_n458));
  AND3_X1   g257(.A1(new_n449), .A2(KEYINPUT92), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT92), .B1(new_n449), .B2(new_n458), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n456), .A2(new_n457), .A3(new_n461), .A4(new_n447), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n454), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n450), .B1(new_n461), .B2(new_n455), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  XOR2_X1   g265(.A(KEYINPUT95), .B(KEYINPUT21), .Z(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AND2_X1   g267(.A1(G231gat), .A2(G233gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n468), .B(new_n469), .ZN(new_n470));
  XOR2_X1   g269(.A(KEYINPUT96), .B(KEYINPUT19), .Z(new_n471));
  XNOR2_X1  g270(.A(new_n470), .B(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(G127gat), .B(G155gat), .ZN(new_n473));
  XOR2_X1   g272(.A(new_n473), .B(KEYINPUT20), .Z(new_n474));
  XNOR2_X1  g273(.A(new_n472), .B(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(G15gat), .B(G22gat), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT16), .ZN(new_n477));
  OR2_X1    g276(.A1(new_n477), .A2(G1gat), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  OR2_X1    g278(.A1(new_n479), .A2(KEYINPUT88), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n476), .A2(G1gat), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n481), .A2(G8gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n479), .A2(KEYINPUT88), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n480), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT89), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n480), .A2(new_n482), .A3(new_n483), .A4(KEYINPUT89), .ZN(new_n487));
  INV_X1    g286(.A(new_n479), .ZN(new_n488));
  OAI21_X1  g287(.A(G8gat), .B1(new_n488), .B2(new_n481), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n486), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n490), .B(KEYINPUT91), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n463), .A2(KEYINPUT97), .A3(new_n465), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT97), .B1(new_n463), .B2(new_n465), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n491), .B1(KEYINPUT21), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n475), .A2(new_n495), .ZN(new_n496));
  OR2_X1    g295(.A1(new_n472), .A2(new_n474), .ZN(new_n497));
  INV_X1    g296(.A(new_n495), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n472), .A2(new_n474), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  XOR2_X1   g300(.A(G183gat), .B(G211gat), .Z(new_n502));
  NOR2_X1   g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n502), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n504), .B1(new_n496), .B2(new_n500), .ZN(new_n505));
  XOR2_X1   g304(.A(G134gat), .B(G162gat), .Z(new_n506));
  XNOR2_X1  g305(.A(G43gat), .B(G50gat), .ZN(new_n507));
  NOR2_X1   g306(.A1(G29gat), .A2(G36gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n508), .B(KEYINPUT14), .ZN(new_n509));
  AND2_X1   g308(.A1(G29gat), .A2(G36gat), .ZN(new_n510));
  OAI211_X1 g309(.A(KEYINPUT15), .B(new_n507), .C1(new_n509), .C2(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n509), .B(KEYINPUT87), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n510), .B1(new_n507), .B2(KEYINPUT15), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n513), .B1(KEYINPUT15), .B2(new_n507), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n511), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(KEYINPUT17), .ZN(new_n516));
  XNOR2_X1  g315(.A(G99gat), .B(G106gat), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(G99gat), .A2(G106gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT8), .ZN(new_n520));
  NAND2_X1  g319(.A1(G85gat), .A2(G92gat), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT7), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n520), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  AND2_X1   g324(.A1(KEYINPUT98), .A2(G92gat), .ZN(new_n526));
  NOR2_X1   g325(.A1(KEYINPUT98), .A2(G92gat), .ZN(new_n527));
  NOR3_X1   g326(.A1(new_n526), .A2(new_n527), .A3(G85gat), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n518), .B1(new_n525), .B2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT99), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OAI211_X1 g330(.A(KEYINPUT99), .B(new_n518), .C1(new_n525), .C2(new_n528), .ZN(new_n532));
  INV_X1    g331(.A(new_n527), .ZN(new_n533));
  INV_X1    g332(.A(G85gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(KEYINPUT98), .A2(G92gat), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  AOI22_X1  g335(.A1(new_n522), .A2(new_n521), .B1(new_n519), .B2(KEYINPUT8), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n536), .A2(new_n537), .A3(new_n517), .A4(new_n524), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n531), .A2(new_n532), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n516), .A2(new_n539), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n531), .A2(new_n532), .A3(new_n538), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n515), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n540), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G190gat), .B(G218gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(KEYINPUT100), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n540), .A2(new_n546), .A3(new_n542), .A4(new_n543), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n548), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n550), .B1(new_n548), .B2(new_n551), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n506), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n554), .ZN(new_n556));
  INV_X1    g355(.A(new_n506), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n556), .A2(new_n552), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  NOR3_X1   g358(.A1(new_n503), .A2(new_n505), .A3(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(G230gat), .A2(G233gat), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  AND2_X1   g362(.A1(new_n529), .A2(new_n538), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n463), .A2(new_n465), .A3(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT10), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n464), .B1(new_n454), .B2(new_n462), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n565), .B(new_n566), .C1(new_n567), .C2(new_n541), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT101), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n466), .A2(new_n539), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n571), .A2(KEYINPUT101), .A3(new_n566), .A4(new_n565), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n531), .A2(KEYINPUT10), .A3(new_n532), .A4(new_n538), .ZN(new_n574));
  NOR3_X1   g373(.A1(new_n492), .A2(new_n493), .A3(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(KEYINPUT102), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n575), .B1(new_n570), .B2(new_n572), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT102), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n563), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G120gat), .B(G148gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(G176gat), .B(G204gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n562), .B1(new_n571), .B2(new_n565), .ZN(new_n586));
  XOR2_X1   g385(.A(new_n586), .B(KEYINPUT103), .Z(new_n587));
  OR3_X1    g386(.A1(new_n582), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n579), .A2(new_n563), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n585), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT104), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n590), .A2(new_n591), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n588), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n491), .A2(new_n515), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n490), .B(KEYINPUT90), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(new_n516), .ZN(new_n597));
  NAND2_X1  g396(.A1(G229gat), .A2(G233gat), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n595), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT18), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(new_n598), .B(KEYINPUT13), .Z(new_n602));
  INV_X1    g401(.A(new_n595), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n491), .A2(new_n515), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n595), .A2(new_n597), .A3(KEYINPUT18), .A4(new_n598), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n601), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(G113gat), .B(G141gat), .Z(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT85), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT86), .ZN(new_n610));
  XNOR2_X1  g409(.A(G169gat), .B(G197gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n610), .B(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(new_n614), .B(KEYINPUT12), .Z(new_n615));
  NAND2_X1  g414(.A1(new_n607), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n615), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n601), .A2(new_n617), .A3(new_n605), .A4(new_n606), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NOR4_X1   g419(.A1(new_n440), .A2(new_n561), .A3(new_n594), .A4(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n395), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g423(.A(KEYINPUT16), .B(G8gat), .Z(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(KEYINPUT105), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n621), .A2(new_n386), .A3(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n627), .A2(KEYINPUT42), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT42), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n621), .A2(new_n386), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n629), .B1(new_n630), .B2(G8gat), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n628), .B1(new_n627), .B2(new_n631), .ZN(G1325gat));
  INV_X1    g431(.A(G15gat), .ZN(new_n633));
  INV_X1    g432(.A(new_n362), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n621), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n438), .B(KEYINPUT106), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n635), .B1(new_n638), .B2(new_n633), .ZN(G1326gat));
  NAND2_X1  g438(.A1(new_n621), .A2(new_n403), .ZN(new_n640));
  XNOR2_X1  g439(.A(KEYINPUT43), .B(G22gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(G1327gat));
  OAI21_X1  g441(.A(new_n559), .B1(new_n402), .B2(new_n439), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n503), .A2(new_n505), .ZN(new_n645));
  NOR3_X1   g444(.A1(new_n645), .A2(new_n594), .A3(new_n620), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  NOR3_X1   g446(.A1(new_n647), .A2(G29gat), .A3(new_n395), .ZN(new_n648));
  OR2_X1    g447(.A1(new_n648), .A2(KEYINPUT45), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(KEYINPUT45), .ZN(new_n650));
  INV_X1    g449(.A(G29gat), .ZN(new_n651));
  AND2_X1   g450(.A1(KEYINPUT107), .A2(KEYINPUT44), .ZN(new_n652));
  NOR2_X1   g451(.A1(KEYINPUT107), .A2(KEYINPUT44), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n643), .A2(new_n654), .ZN(new_n655));
  OAI211_X1 g454(.A(new_n559), .B(new_n652), .C1(new_n402), .C2(new_n439), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AND3_X1   g456(.A1(new_n657), .A2(new_n622), .A3(new_n646), .ZN(new_n658));
  OAI211_X1 g457(.A(new_n649), .B(new_n650), .C1(new_n651), .C2(new_n658), .ZN(G1328gat));
  NOR3_X1   g458(.A1(new_n647), .A2(G36gat), .A3(new_n385), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(KEYINPUT46), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n657), .A2(new_n386), .A3(new_n646), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(G36gat), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n661), .A2(new_n663), .ZN(G1329gat));
  NAND4_X1  g463(.A1(new_n657), .A2(new_n436), .A3(new_n437), .A4(new_n646), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n665), .A2(G43gat), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n647), .A2(G43gat), .A3(new_n362), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT47), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n657), .A2(new_n636), .A3(new_n646), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n667), .B1(new_n670), .B2(G43gat), .ZN(new_n671));
  OAI22_X1  g470(.A1(new_n666), .A2(new_n669), .B1(new_n671), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g471(.A(G50gat), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n655), .A2(new_n403), .A3(new_n656), .A4(new_n646), .ZN(new_n674));
  OR2_X1    g473(.A1(new_n674), .A2(KEYINPUT108), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(KEYINPUT108), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n673), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n644), .A2(new_n673), .A3(new_n403), .A4(new_n646), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(KEYINPUT48), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n674), .A2(G50gat), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n680), .A2(new_n678), .ZN(new_n681));
  OAI22_X1  g480(.A1(new_n677), .A2(new_n679), .B1(KEYINPUT48), .B2(new_n681), .ZN(G1331gat));
  NAND3_X1  g481(.A1(new_n405), .A2(new_n434), .A3(new_n438), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n401), .A2(KEYINPUT35), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n683), .B1(new_n684), .B2(new_n387), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n685), .A2(new_n560), .A3(new_n594), .A4(new_n620), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n395), .B(KEYINPUT109), .ZN(new_n687));
  OR2_X1    g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(G57gat), .ZN(G1332gat));
  INV_X1    g488(.A(new_n686), .ZN(new_n690));
  XOR2_X1   g489(.A(KEYINPUT49), .B(G64gat), .Z(new_n691));
  NAND3_X1  g490(.A1(new_n690), .A2(new_n386), .A3(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n693), .B1(new_n686), .B2(new_n385), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT110), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(G1333gat));
  INV_X1    g496(.A(G71gat), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n698), .B1(new_n686), .B2(new_n362), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n636), .A2(G71gat), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n699), .B1(new_n686), .B2(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g501(.A1(new_n690), .A2(new_n403), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g503(.A1(new_n645), .A2(new_n619), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n685), .A2(KEYINPUT51), .A3(new_n559), .A4(new_n705), .ZN(new_n706));
  OAI211_X1 g505(.A(new_n559), .B(new_n705), .C1(new_n402), .C2(new_n439), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT51), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n622), .A2(new_n594), .A3(new_n534), .ZN(new_n711));
  XOR2_X1   g510(.A(new_n711), .B(KEYINPUT112), .Z(new_n712));
  NAND2_X1  g511(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n594), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n645), .A2(new_n714), .A3(new_n619), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n657), .A2(new_n622), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(KEYINPUT111), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(G85gat), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n716), .A2(KEYINPUT111), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n713), .B1(new_n718), .B2(new_n719), .ZN(G1336gat));
  NAND4_X1  g519(.A1(new_n655), .A2(new_n386), .A3(new_n656), .A4(new_n715), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n533), .A2(new_n535), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT113), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n714), .A2(new_n385), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n726), .A2(G92gat), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n728), .B1(new_n706), .B2(new_n709), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n723), .B1(new_n724), .B2(new_n729), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n729), .A2(new_n724), .ZN(new_n731));
  OAI21_X1  g530(.A(KEYINPUT52), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT114), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n706), .A2(new_n709), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n733), .B1(new_n734), .B2(new_n728), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT52), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n729), .A2(KEYINPUT114), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n735), .A2(new_n736), .A3(new_n723), .A4(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n732), .A2(new_n738), .ZN(G1337gat));
  AND3_X1   g538(.A1(new_n657), .A2(new_n636), .A3(new_n715), .ZN(new_n740));
  INV_X1    g539(.A(G99gat), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n634), .A2(new_n741), .A3(new_n594), .ZN(new_n742));
  OAI22_X1  g541(.A1(new_n740), .A2(new_n741), .B1(new_n734), .B2(new_n742), .ZN(G1338gat));
  NOR3_X1   g542(.A1(new_n714), .A2(G106gat), .A3(new_n248), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n710), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n655), .A2(new_n403), .A3(new_n656), .A4(new_n715), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(G106gat), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT53), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n745), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT116), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n744), .B(KEYINPUT115), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n747), .B1(new_n734), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(KEYINPUT53), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n745), .A2(new_n747), .A3(KEYINPUT116), .A4(new_n748), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n751), .A2(new_n754), .A3(new_n755), .ZN(G1339gat));
  INV_X1    g555(.A(new_n645), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT55), .ZN(new_n758));
  AOI211_X1 g557(.A(KEYINPUT102), .B(new_n575), .C1(new_n570), .C2(new_n572), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n580), .B1(new_n573), .B2(new_n576), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n562), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT117), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT54), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n763), .B1(new_n579), .B2(new_n563), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n761), .A2(new_n762), .A3(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n585), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n766), .B1(new_n589), .B2(new_n763), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n762), .B1(new_n761), .B2(new_n764), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n758), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(new_n764), .ZN(new_n771));
  OAI21_X1  g570(.A(KEYINPUT117), .B1(new_n582), .B2(new_n771), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n772), .A2(KEYINPUT55), .A3(new_n765), .A4(new_n767), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n770), .A2(new_n588), .A3(new_n619), .A4(new_n773), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n603), .A2(new_n604), .A3(new_n602), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n598), .B1(new_n595), .B2(new_n597), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n614), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n594), .A2(new_n618), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n559), .B1(new_n774), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n618), .A2(new_n777), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n780), .B1(new_n558), .B2(new_n555), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n781), .A2(new_n588), .A3(new_n773), .A4(new_n770), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n757), .B1(new_n779), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n560), .A2(new_n714), .A3(new_n620), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n403), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n362), .A2(new_n395), .A3(new_n386), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(G113gat), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n788), .A2(new_n789), .A3(new_n620), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n687), .B1(new_n784), .B2(new_n785), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n791), .A2(new_n385), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n389), .A2(new_n400), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n619), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n790), .B1(new_n795), .B2(new_n789), .ZN(G1340gat));
  INV_X1    g595(.A(G120gat), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n794), .A2(new_n797), .A3(new_n594), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n786), .A2(new_n594), .A3(new_n787), .ZN(new_n799));
  AND3_X1   g598(.A1(new_n799), .A2(KEYINPUT118), .A3(G120gat), .ZN(new_n800));
  AOI21_X1  g599(.A(KEYINPUT118), .B1(new_n799), .B2(G120gat), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n798), .B1(new_n800), .B2(new_n801), .ZN(G1341gat));
  INV_X1    g601(.A(G127gat), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n794), .A2(new_n803), .A3(new_n645), .ZN(new_n804));
  OAI21_X1  g603(.A(G127gat), .B1(new_n788), .B2(new_n757), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(G1342gat));
  INV_X1    g605(.A(G134gat), .ZN(new_n807));
  INV_X1    g606(.A(new_n559), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n808), .A2(new_n386), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n791), .A2(new_n807), .A3(new_n793), .A4(new_n809), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n810), .A2(KEYINPUT56), .ZN(new_n811));
  XOR2_X1   g610(.A(new_n811), .B(KEYINPUT119), .Z(new_n812));
  NAND2_X1  g611(.A1(new_n810), .A2(KEYINPUT56), .ZN(new_n813));
  OAI21_X1  g612(.A(G134gat), .B1(new_n788), .B2(new_n808), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(G1343gat));
  NAND3_X1  g614(.A1(new_n438), .A2(new_n622), .A3(new_n385), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n248), .B1(new_n784), .B2(new_n785), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT57), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n816), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n782), .B1(new_n779), .B2(KEYINPUT120), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT120), .ZN(new_n821));
  AOI211_X1 g620(.A(new_n821), .B(new_n559), .C1(new_n774), .C2(new_n778), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n757), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n248), .B1(new_n823), .B2(new_n785), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n619), .B(new_n819), .C1(new_n824), .C2(new_n818), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(G141gat), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT122), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n636), .A2(new_n248), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n620), .A2(G141gat), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n830), .B(KEYINPUT121), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n792), .A2(new_n829), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n826), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n828), .A2(new_n833), .A3(KEYINPUT58), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT58), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n826), .B(new_n832), .C1(new_n827), .C2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n834), .A2(new_n836), .ZN(G1344gat));
  NOR2_X1   g636(.A1(new_n714), .A2(G148gat), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n792), .A2(new_n829), .A3(new_n838), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(KEYINPUT123), .ZN(new_n840));
  XOR2_X1   g639(.A(KEYINPUT124), .B(KEYINPUT59), .Z(new_n841));
  AND2_X1   g640(.A1(new_n784), .A2(new_n785), .ZN(new_n842));
  OAI21_X1  g641(.A(KEYINPUT57), .B1(new_n842), .B2(new_n248), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n817), .A2(new_n818), .ZN(new_n844));
  AND3_X1   g643(.A1(new_n843), .A2(new_n594), .A3(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n816), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n841), .B1(new_n847), .B2(G148gat), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n594), .B(new_n819), .C1(new_n824), .C2(new_n818), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT59), .ZN(new_n850));
  AND3_X1   g649(.A1(new_n849), .A2(new_n850), .A3(G148gat), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n840), .B1(new_n848), .B2(new_n851), .ZN(G1345gat));
  OAI21_X1  g651(.A(new_n819), .B1(new_n824), .B2(new_n818), .ZN(new_n853));
  OAI21_X1  g652(.A(G155gat), .B1(new_n853), .B2(new_n757), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n792), .A2(new_n212), .A3(new_n645), .A4(new_n829), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(G1346gat));
  OAI21_X1  g655(.A(G162gat), .B1(new_n853), .B2(new_n808), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n829), .A2(new_n213), .A3(new_n791), .A4(new_n809), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(G1347gat));
  NAND2_X1  g658(.A1(new_n687), .A2(new_n386), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n860), .A2(new_n362), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n786), .A2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(G169gat), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n862), .A2(new_n863), .A3(new_n620), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n622), .B1(new_n784), .B2(new_n785), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n793), .A2(new_n386), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n619), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n864), .B1(new_n863), .B2(new_n869), .ZN(G1348gat));
  OAI21_X1  g669(.A(G176gat), .B1(new_n862), .B2(new_n714), .ZN(new_n871));
  OR2_X1    g670(.A1(new_n714), .A2(G176gat), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n871), .B1(new_n867), .B2(new_n872), .ZN(G1349gat));
  OAI21_X1  g672(.A(new_n300), .B1(new_n862), .B2(new_n757), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n645), .A2(new_n319), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n874), .B1(new_n867), .B2(new_n875), .ZN(new_n876));
  XNOR2_X1  g675(.A(new_n876), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g676(.A1(new_n868), .A2(new_n320), .A3(new_n559), .ZN(new_n878));
  OAI21_X1  g677(.A(G190gat), .B1(new_n862), .B2(new_n808), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n879), .A2(KEYINPUT61), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n879), .A2(KEYINPUT61), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n878), .B1(new_n880), .B2(new_n881), .ZN(G1351gat));
  XNOR2_X1  g681(.A(KEYINPUT126), .B(G197gat), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n829), .A2(new_n386), .A3(new_n865), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT125), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n829), .A2(KEYINPUT125), .A3(new_n865), .A4(new_n386), .ZN(new_n888));
  AOI211_X1 g687(.A(new_n620), .B(new_n884), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n636), .A2(new_n860), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n843), .A2(new_n619), .A3(new_n844), .A4(new_n890), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n891), .A2(new_n884), .ZN(new_n892));
  OAI21_X1  g691(.A(KEYINPUT127), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT127), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n891), .A2(new_n884), .ZN(new_n895));
  INV_X1    g694(.A(new_n887), .ZN(new_n896));
  INV_X1    g695(.A(new_n888), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n620), .A2(new_n884), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n894), .B(new_n895), .C1(new_n898), .C2(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n893), .A2(new_n901), .ZN(G1352gat));
  NAND2_X1  g701(.A1(new_n829), .A2(new_n865), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n903), .A2(G204gat), .A3(new_n726), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n904), .B(KEYINPUT62), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n845), .A2(new_n890), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(G204gat), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n905), .A2(new_n907), .ZN(G1353gat));
  NAND4_X1  g707(.A1(new_n843), .A2(new_n645), .A3(new_n844), .A4(new_n890), .ZN(new_n909));
  AND3_X1   g708(.A1(new_n909), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n910));
  AOI21_X1  g709(.A(KEYINPUT63), .B1(new_n909), .B2(G211gat), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n645), .A2(new_n219), .ZN(new_n912));
  OAI22_X1  g711(.A1(new_n910), .A2(new_n911), .B1(new_n898), .B2(new_n912), .ZN(G1354gat));
  NAND3_X1  g712(.A1(new_n843), .A2(new_n844), .A3(new_n890), .ZN(new_n914));
  OAI21_X1  g713(.A(G218gat), .B1(new_n914), .B2(new_n808), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n559), .A2(new_n220), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n915), .B1(new_n898), .B2(new_n916), .ZN(G1355gat));
endmodule


