

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U554 ( .A1(n695), .A2(n694), .ZN(n714) );
  XOR2_X1 U555 ( .A(n625), .B(KEYINPUT31), .Z(n518) );
  AND2_X1 U556 ( .A1(n614), .A2(G8), .ZN(n519) );
  OR2_X1 U557 ( .A1(n718), .A2(n717), .ZN(n520) );
  XNOR2_X1 U558 ( .A(KEYINPUT102), .B(KEYINPUT27), .ZN(n626) );
  XNOR2_X1 U559 ( .A(n627), .B(n626), .ZN(n629) );
  INV_X1 U560 ( .A(KEYINPUT104), .ZN(n678) );
  XNOR2_X1 U561 ( .A(n679), .B(n678), .ZN(n689) );
  NAND2_X1 U562 ( .A1(n741), .A2(n613), .ZN(n619) );
  NAND2_X1 U563 ( .A1(G8), .A2(n619), .ZN(n718) );
  INV_X1 U564 ( .A(KEYINPUT17), .ZN(n526) );
  NAND2_X1 U565 ( .A1(n719), .A2(n520), .ZN(n720) );
  XNOR2_X1 U566 ( .A(n526), .B(KEYINPUT66), .ZN(n527) );
  NOR2_X1 U567 ( .A1(G2105), .A2(n522), .ZN(n897) );
  NOR2_X1 U568 ( .A1(G651), .A2(n591), .ZN(n799) );
  NOR2_X1 U569 ( .A1(n774), .A2(n773), .ZN(n775) );
  NOR2_X1 U570 ( .A1(n560), .A2(n559), .ZN(n612) );
  NOR2_X1 U571 ( .A1(n532), .A2(n531), .ZN(G160) );
  INV_X1 U572 ( .A(G2104), .ZN(n522) );
  NAND2_X1 U573 ( .A1(G101), .A2(n897), .ZN(n521) );
  XOR2_X1 U574 ( .A(KEYINPUT23), .B(n521), .Z(n525) );
  AND2_X1 U575 ( .A1(n522), .A2(G2105), .ZN(n901) );
  NAND2_X1 U576 ( .A1(G125), .A2(n901), .ZN(n523) );
  XOR2_X1 U577 ( .A(KEYINPUT65), .B(n523), .Z(n524) );
  NAND2_X1 U578 ( .A1(n525), .A2(n524), .ZN(n532) );
  AND2_X1 U579 ( .A1(G2104), .A2(G2105), .ZN(n902) );
  NAND2_X1 U580 ( .A1(G113), .A2(n902), .ZN(n530) );
  NOR2_X1 U581 ( .A1(G2104), .A2(G2105), .ZN(n528) );
  XNOR2_X2 U582 ( .A(n528), .B(n527), .ZN(n898) );
  NAND2_X1 U583 ( .A1(G137), .A2(n898), .ZN(n529) );
  NAND2_X1 U584 ( .A1(n530), .A2(n529), .ZN(n531) );
  INV_X1 U585 ( .A(G651), .ZN(n538) );
  NOR2_X1 U586 ( .A1(G543), .A2(n538), .ZN(n533) );
  XOR2_X1 U587 ( .A(KEYINPUT1), .B(n533), .Z(n800) );
  NAND2_X1 U588 ( .A1(n800), .A2(G64), .ZN(n536) );
  XNOR2_X1 U589 ( .A(G543), .B(KEYINPUT0), .ZN(n534) );
  XNOR2_X1 U590 ( .A(n534), .B(KEYINPUT67), .ZN(n591) );
  NAND2_X1 U591 ( .A1(n799), .A2(G52), .ZN(n535) );
  NAND2_X1 U592 ( .A1(n536), .A2(n535), .ZN(n543) );
  NOR2_X1 U593 ( .A1(G543), .A2(G651), .ZN(n796) );
  NAND2_X1 U594 ( .A1(n796), .A2(G90), .ZN(n537) );
  XNOR2_X1 U595 ( .A(n537), .B(KEYINPUT70), .ZN(n540) );
  NOR2_X1 U596 ( .A1(n591), .A2(n538), .ZN(n794) );
  NAND2_X1 U597 ( .A1(G77), .A2(n794), .ZN(n539) );
  NAND2_X1 U598 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U599 ( .A(KEYINPUT9), .B(n541), .Z(n542) );
  NOR2_X1 U600 ( .A1(n543), .A2(n542), .ZN(G171) );
  INV_X1 U601 ( .A(G171), .ZN(G301) );
  AND2_X1 U602 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U603 ( .A1(n898), .A2(G135), .ZN(n544) );
  XNOR2_X1 U604 ( .A(n544), .B(KEYINPUT80), .ZN(n551) );
  NAND2_X1 U605 ( .A1(G99), .A2(n897), .ZN(n546) );
  NAND2_X1 U606 ( .A1(G111), .A2(n902), .ZN(n545) );
  NAND2_X1 U607 ( .A1(n546), .A2(n545), .ZN(n549) );
  NAND2_X1 U608 ( .A1(n901), .A2(G123), .ZN(n547) );
  XOR2_X1 U609 ( .A(KEYINPUT18), .B(n547), .Z(n548) );
  NOR2_X1 U610 ( .A1(n549), .A2(n548), .ZN(n550) );
  NAND2_X1 U611 ( .A1(n551), .A2(n550), .ZN(n927) );
  XNOR2_X1 U612 ( .A(G2096), .B(n927), .ZN(n552) );
  OR2_X1 U613 ( .A1(G2100), .A2(n552), .ZN(G156) );
  NAND2_X1 U614 ( .A1(G138), .A2(n898), .ZN(n554) );
  NAND2_X1 U615 ( .A1(G102), .A2(n897), .ZN(n553) );
  NAND2_X1 U616 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U617 ( .A(n555), .B(KEYINPUT95), .ZN(n557) );
  NAND2_X1 U618 ( .A1(G126), .A2(n901), .ZN(n556) );
  NAND2_X1 U619 ( .A1(n557), .A2(n556), .ZN(n560) );
  NAND2_X1 U620 ( .A1(n902), .A2(G114), .ZN(n558) );
  XOR2_X1 U621 ( .A(KEYINPUT94), .B(n558), .Z(n559) );
  BUF_X1 U622 ( .A(n612), .Z(G164) );
  NAND2_X1 U623 ( .A1(n796), .A2(G89), .ZN(n561) );
  XNOR2_X1 U624 ( .A(KEYINPUT4), .B(n561), .ZN(n564) );
  NAND2_X1 U625 ( .A1(n794), .A2(G76), .ZN(n562) );
  XOR2_X1 U626 ( .A(KEYINPUT77), .B(n562), .Z(n563) );
  NAND2_X1 U627 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U628 ( .A(n565), .B(KEYINPUT5), .ZN(n570) );
  NAND2_X1 U629 ( .A1(G51), .A2(n799), .ZN(n567) );
  NAND2_X1 U630 ( .A1(G63), .A2(n800), .ZN(n566) );
  NAND2_X1 U631 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U632 ( .A(KEYINPUT6), .B(n568), .Z(n569) );
  NAND2_X1 U633 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U634 ( .A(n571), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U635 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U636 ( .A1(G78), .A2(n794), .ZN(n573) );
  NAND2_X1 U637 ( .A1(G53), .A2(n799), .ZN(n572) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n576) );
  NAND2_X1 U639 ( .A1(G91), .A2(n796), .ZN(n574) );
  XNOR2_X1 U640 ( .A(KEYINPUT71), .B(n574), .ZN(n575) );
  NOR2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n578) );
  NAND2_X1 U642 ( .A1(n800), .A2(G65), .ZN(n577) );
  NAND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(G299) );
  NAND2_X1 U644 ( .A1(G62), .A2(n800), .ZN(n585) );
  NAND2_X1 U645 ( .A1(G88), .A2(n796), .ZN(n580) );
  NAND2_X1 U646 ( .A1(G50), .A2(n799), .ZN(n579) );
  NAND2_X1 U647 ( .A1(n580), .A2(n579), .ZN(n583) );
  NAND2_X1 U648 ( .A1(G75), .A2(n794), .ZN(n581) );
  XNOR2_X1 U649 ( .A(KEYINPUT87), .B(n581), .ZN(n582) );
  NOR2_X1 U650 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U651 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n586), .B(KEYINPUT88), .ZN(G303) );
  NAND2_X1 U653 ( .A1(G49), .A2(n799), .ZN(n588) );
  NAND2_X1 U654 ( .A1(G74), .A2(G651), .ZN(n587) );
  NAND2_X1 U655 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U656 ( .A1(n800), .A2(n589), .ZN(n590) );
  XOR2_X1 U657 ( .A(KEYINPUT83), .B(n590), .Z(n593) );
  NAND2_X1 U658 ( .A1(n591), .A2(G87), .ZN(n592) );
  NAND2_X1 U659 ( .A1(n593), .A2(n592), .ZN(G288) );
  NAND2_X1 U660 ( .A1(n800), .A2(G61), .ZN(n594) );
  XNOR2_X1 U661 ( .A(n594), .B(KEYINPUT84), .ZN(n596) );
  NAND2_X1 U662 ( .A1(G86), .A2(n796), .ZN(n595) );
  NAND2_X1 U663 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U664 ( .A(KEYINPUT85), .B(n597), .ZN(n603) );
  NAND2_X1 U665 ( .A1(G73), .A2(n794), .ZN(n598) );
  XOR2_X1 U666 ( .A(KEYINPUT2), .B(n598), .Z(n601) );
  NAND2_X1 U667 ( .A1(n799), .A2(G48), .ZN(n599) );
  XOR2_X1 U668 ( .A(KEYINPUT86), .B(n599), .Z(n600) );
  NOR2_X1 U669 ( .A1(n601), .A2(n600), .ZN(n602) );
  NAND2_X1 U670 ( .A1(n603), .A2(n602), .ZN(G305) );
  NAND2_X1 U671 ( .A1(G85), .A2(n796), .ZN(n605) );
  NAND2_X1 U672 ( .A1(G72), .A2(n794), .ZN(n604) );
  NAND2_X1 U673 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U674 ( .A(KEYINPUT68), .B(n606), .ZN(n609) );
  NAND2_X1 U675 ( .A1(G60), .A2(n800), .ZN(n607) );
  XNOR2_X1 U676 ( .A(KEYINPUT69), .B(n607), .ZN(n608) );
  NOR2_X1 U677 ( .A1(n609), .A2(n608), .ZN(n611) );
  NAND2_X1 U678 ( .A1(n799), .A2(G47), .ZN(n610) );
  NAND2_X1 U679 ( .A1(n611), .A2(n610), .ZN(G290) );
  INV_X1 U680 ( .A(KEYINPUT40), .ZN(n776) );
  NOR2_X1 U681 ( .A1(n612), .A2(G1384), .ZN(n741) );
  NAND2_X1 U682 ( .A1(G160), .A2(G40), .ZN(n740) );
  INV_X1 U683 ( .A(n740), .ZN(n613) );
  NOR2_X1 U684 ( .A1(G1966), .A2(n718), .ZN(n690) );
  INV_X1 U685 ( .A(n690), .ZN(n615) );
  NOR2_X1 U686 ( .A1(G2084), .A2(n619), .ZN(n688) );
  INV_X1 U687 ( .A(n688), .ZN(n614) );
  NAND2_X1 U688 ( .A1(n615), .A2(n519), .ZN(n616) );
  XNOR2_X1 U689 ( .A(n616), .B(KEYINPUT30), .ZN(n617) );
  NOR2_X1 U690 ( .A1(n617), .A2(G168), .ZN(n618) );
  XNOR2_X1 U691 ( .A(n618), .B(KEYINPUT103), .ZN(n624) );
  INV_X1 U692 ( .A(n619), .ZN(n653) );
  XOR2_X1 U693 ( .A(KEYINPUT25), .B(G2078), .Z(n982) );
  NAND2_X1 U694 ( .A1(n653), .A2(n982), .ZN(n621) );
  NAND2_X1 U695 ( .A1(G1961), .A2(n619), .ZN(n620) );
  NAND2_X1 U696 ( .A1(n621), .A2(n620), .ZN(n622) );
  XOR2_X1 U697 ( .A(KEYINPUT101), .B(n622), .Z(n674) );
  NAND2_X1 U698 ( .A1(n674), .A2(G301), .ZN(n623) );
  NAND2_X1 U699 ( .A1(n624), .A2(n623), .ZN(n625) );
  NAND2_X1 U700 ( .A1(G2072), .A2(n653), .ZN(n627) );
  AND2_X1 U701 ( .A1(n619), .A2(G1956), .ZN(n628) );
  NOR2_X1 U702 ( .A1(n629), .A2(n628), .ZN(n632) );
  INV_X1 U703 ( .A(G299), .ZN(n806) );
  NOR2_X1 U704 ( .A1(n632), .A2(n806), .ZN(n631) );
  INV_X1 U705 ( .A(KEYINPUT28), .ZN(n630) );
  XNOR2_X1 U706 ( .A(n631), .B(n630), .ZN(n672) );
  NAND2_X1 U707 ( .A1(n632), .A2(n806), .ZN(n670) );
  NAND2_X1 U708 ( .A1(n796), .A2(G81), .ZN(n633) );
  XNOR2_X1 U709 ( .A(n633), .B(KEYINPUT12), .ZN(n635) );
  NAND2_X1 U710 ( .A1(G68), .A2(n794), .ZN(n634) );
  NAND2_X1 U711 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U712 ( .A(n636), .B(KEYINPUT13), .ZN(n638) );
  NAND2_X1 U713 ( .A1(G43), .A2(n799), .ZN(n637) );
  NAND2_X1 U714 ( .A1(n638), .A2(n637), .ZN(n642) );
  NAND2_X1 U715 ( .A1(G56), .A2(n800), .ZN(n639) );
  XNOR2_X1 U716 ( .A(n639), .B(KEYINPUT73), .ZN(n640) );
  XNOR2_X1 U717 ( .A(n640), .B(KEYINPUT14), .ZN(n641) );
  NOR2_X1 U718 ( .A1(n642), .A2(n641), .ZN(n643) );
  XOR2_X1 U719 ( .A(KEYINPUT74), .B(n643), .Z(n966) );
  XNOR2_X1 U720 ( .A(KEYINPUT64), .B(KEYINPUT26), .ZN(n660) );
  NOR2_X1 U721 ( .A1(G1996), .A2(n660), .ZN(n644) );
  NOR2_X1 U722 ( .A1(n966), .A2(n644), .ZN(n657) );
  NAND2_X1 U723 ( .A1(G92), .A2(n796), .ZN(n646) );
  NAND2_X1 U724 ( .A1(G66), .A2(n800), .ZN(n645) );
  NAND2_X1 U725 ( .A1(n646), .A2(n645), .ZN(n651) );
  NAND2_X1 U726 ( .A1(G79), .A2(n794), .ZN(n648) );
  NAND2_X1 U727 ( .A1(G54), .A2(n799), .ZN(n647) );
  NAND2_X1 U728 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U729 ( .A(KEYINPUT76), .B(n649), .ZN(n650) );
  NOR2_X1 U730 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U731 ( .A(n652), .B(KEYINPUT15), .ZN(n953) );
  NAND2_X1 U732 ( .A1(G1348), .A2(n619), .ZN(n655) );
  NAND2_X1 U733 ( .A1(G2067), .A2(n653), .ZN(n654) );
  NAND2_X1 U734 ( .A1(n655), .A2(n654), .ZN(n666) );
  NAND2_X1 U735 ( .A1(n953), .A2(n666), .ZN(n656) );
  NAND2_X1 U736 ( .A1(n657), .A2(n656), .ZN(n665) );
  INV_X1 U737 ( .A(G1341), .ZN(n658) );
  NAND2_X1 U738 ( .A1(n658), .A2(n660), .ZN(n659) );
  NAND2_X1 U739 ( .A1(n659), .A2(n619), .ZN(n663) );
  INV_X1 U740 ( .A(G1996), .ZN(n762) );
  NOR2_X1 U741 ( .A1(n762), .A2(n619), .ZN(n661) );
  NAND2_X1 U742 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U743 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U744 ( .A1(n665), .A2(n664), .ZN(n668) );
  NOR2_X1 U745 ( .A1(n666), .A2(n953), .ZN(n667) );
  NOR2_X1 U746 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U747 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U748 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U749 ( .A(n673), .B(KEYINPUT29), .ZN(n676) );
  NOR2_X1 U750 ( .A1(G301), .A2(n674), .ZN(n675) );
  NOR2_X1 U751 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U752 ( .A1(n518), .A2(n677), .ZN(n679) );
  NAND2_X1 U753 ( .A1(n689), .A2(G286), .ZN(n686) );
  INV_X1 U754 ( .A(G8), .ZN(n684) );
  NOR2_X1 U755 ( .A1(G1971), .A2(n718), .ZN(n681) );
  NOR2_X1 U756 ( .A1(G2090), .A2(n619), .ZN(n680) );
  NOR2_X1 U757 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U758 ( .A1(n682), .A2(G303), .ZN(n683) );
  OR2_X1 U759 ( .A1(n684), .A2(n683), .ZN(n685) );
  AND2_X1 U760 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U761 ( .A(n687), .B(KEYINPUT32), .ZN(n695) );
  NAND2_X1 U762 ( .A1(G8), .A2(n688), .ZN(n693) );
  INV_X1 U763 ( .A(n689), .ZN(n691) );
  NOR2_X1 U764 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U765 ( .A1(n693), .A2(n692), .ZN(n694) );
  INV_X1 U766 ( .A(n714), .ZN(n697) );
  OR2_X1 U767 ( .A1(G303), .A2(G1971), .ZN(n696) );
  OR2_X1 U768 ( .A1(G1976), .A2(G288), .ZN(n699) );
  NAND2_X1 U769 ( .A1(n696), .A2(n699), .ZN(n972) );
  NOR2_X1 U770 ( .A1(n697), .A2(n972), .ZN(n698) );
  NOR2_X1 U771 ( .A1(n718), .A2(n698), .ZN(n705) );
  NAND2_X1 U772 ( .A1(G1976), .A2(G288), .ZN(n956) );
  INV_X1 U773 ( .A(KEYINPUT33), .ZN(n707) );
  OR2_X1 U774 ( .A1(n718), .A2(n699), .ZN(n700) );
  NOR2_X1 U775 ( .A1(n707), .A2(n700), .ZN(n701) );
  XNOR2_X1 U776 ( .A(n701), .B(KEYINPUT105), .ZN(n706) );
  AND2_X1 U777 ( .A1(n956), .A2(n706), .ZN(n703) );
  XNOR2_X1 U778 ( .A(G1981), .B(G305), .ZN(n962) );
  INV_X1 U779 ( .A(n962), .ZN(n702) );
  AND2_X1 U780 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U781 ( .A1(n705), .A2(n704), .ZN(n711) );
  INV_X1 U782 ( .A(n706), .ZN(n708) );
  OR2_X1 U783 ( .A1(n708), .A2(n707), .ZN(n709) );
  OR2_X1 U784 ( .A1(n962), .A2(n709), .ZN(n710) );
  NAND2_X1 U785 ( .A1(n711), .A2(n710), .ZN(n721) );
  NOR2_X1 U786 ( .A1(G2090), .A2(G303), .ZN(n712) );
  NAND2_X1 U787 ( .A1(G8), .A2(n712), .ZN(n713) );
  NAND2_X1 U788 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U789 ( .A1(n715), .A2(n718), .ZN(n719) );
  NOR2_X1 U790 ( .A1(G1981), .A2(G305), .ZN(n716) );
  XOR2_X1 U791 ( .A(n716), .B(KEYINPUT24), .Z(n717) );
  NOR2_X1 U792 ( .A1(n721), .A2(n720), .ZN(n758) );
  NAND2_X1 U793 ( .A1(G129), .A2(n901), .ZN(n723) );
  NAND2_X1 U794 ( .A1(G117), .A2(n902), .ZN(n722) );
  NAND2_X1 U795 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U796 ( .A(KEYINPUT100), .B(n724), .ZN(n729) );
  NAND2_X1 U797 ( .A1(n897), .A2(G105), .ZN(n725) );
  XNOR2_X1 U798 ( .A(n725), .B(KEYINPUT38), .ZN(n727) );
  NAND2_X1 U799 ( .A1(G141), .A2(n898), .ZN(n726) );
  NAND2_X1 U800 ( .A1(n727), .A2(n726), .ZN(n728) );
  NOR2_X1 U801 ( .A1(n729), .A2(n728), .ZN(n892) );
  NOR2_X1 U802 ( .A1(n892), .A2(n762), .ZN(n739) );
  NAND2_X1 U803 ( .A1(n902), .A2(G107), .ZN(n736) );
  NAND2_X1 U804 ( .A1(G119), .A2(n901), .ZN(n731) );
  NAND2_X1 U805 ( .A1(G131), .A2(n898), .ZN(n730) );
  NAND2_X1 U806 ( .A1(n731), .A2(n730), .ZN(n734) );
  NAND2_X1 U807 ( .A1(G95), .A2(n897), .ZN(n732) );
  XOR2_X1 U808 ( .A(KEYINPUT98), .B(n732), .Z(n733) );
  NOR2_X1 U809 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U810 ( .A1(n736), .A2(n735), .ZN(n737) );
  XOR2_X1 U811 ( .A(n737), .B(KEYINPUT99), .Z(n893) );
  AND2_X1 U812 ( .A1(G1991), .A2(n893), .ZN(n738) );
  NOR2_X1 U813 ( .A1(n739), .A2(n738), .ZN(n926) );
  NOR2_X1 U814 ( .A1(n741), .A2(n740), .ZN(n771) );
  INV_X1 U815 ( .A(n771), .ZN(n742) );
  NOR2_X1 U816 ( .A1(n926), .A2(n742), .ZN(n761) );
  INV_X1 U817 ( .A(n761), .ZN(n756) );
  XNOR2_X1 U818 ( .A(G1986), .B(G290), .ZN(n959) );
  NAND2_X1 U819 ( .A1(n959), .A2(n771), .ZN(n743) );
  XNOR2_X1 U820 ( .A(n743), .B(KEYINPUT96), .ZN(n754) );
  NAND2_X1 U821 ( .A1(G104), .A2(n897), .ZN(n745) );
  NAND2_X1 U822 ( .A1(G140), .A2(n898), .ZN(n744) );
  NAND2_X1 U823 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U824 ( .A(KEYINPUT34), .B(n746), .ZN(n752) );
  NAND2_X1 U825 ( .A1(G128), .A2(n901), .ZN(n748) );
  NAND2_X1 U826 ( .A1(G116), .A2(n902), .ZN(n747) );
  NAND2_X1 U827 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U828 ( .A(KEYINPUT97), .B(n749), .ZN(n750) );
  XNOR2_X1 U829 ( .A(KEYINPUT35), .B(n750), .ZN(n751) );
  NOR2_X1 U830 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U831 ( .A(KEYINPUT36), .B(n753), .ZN(n912) );
  XNOR2_X1 U832 ( .A(G2067), .B(KEYINPUT37), .ZN(n768) );
  NOR2_X1 U833 ( .A1(n912), .A2(n768), .ZN(n933) );
  NAND2_X1 U834 ( .A1(n771), .A2(n933), .ZN(n766) );
  AND2_X1 U835 ( .A1(n754), .A2(n766), .ZN(n755) );
  NAND2_X1 U836 ( .A1(n756), .A2(n755), .ZN(n757) );
  NOR2_X1 U837 ( .A1(n758), .A2(n757), .ZN(n774) );
  NOR2_X1 U838 ( .A1(G1986), .A2(G290), .ZN(n759) );
  NOR2_X1 U839 ( .A1(G1991), .A2(n893), .ZN(n930) );
  NOR2_X1 U840 ( .A1(n759), .A2(n930), .ZN(n760) );
  NOR2_X1 U841 ( .A1(n761), .A2(n760), .ZN(n764) );
  AND2_X1 U842 ( .A1(n892), .A2(n762), .ZN(n763) );
  XNOR2_X1 U843 ( .A(n763), .B(KEYINPUT106), .ZN(n939) );
  NOR2_X1 U844 ( .A1(n764), .A2(n939), .ZN(n765) );
  XNOR2_X1 U845 ( .A(n765), .B(KEYINPUT39), .ZN(n767) );
  NAND2_X1 U846 ( .A1(n767), .A2(n766), .ZN(n769) );
  NAND2_X1 U847 ( .A1(n912), .A2(n768), .ZN(n925) );
  NAND2_X1 U848 ( .A1(n769), .A2(n925), .ZN(n770) );
  NAND2_X1 U849 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U850 ( .A(n772), .B(KEYINPUT107), .ZN(n773) );
  XNOR2_X1 U851 ( .A(n776), .B(n775), .ZN(G329) );
  NAND2_X1 U852 ( .A1(G7), .A2(G661), .ZN(n777) );
  XNOR2_X1 U853 ( .A(n777), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U854 ( .A(G223), .ZN(n848) );
  NAND2_X1 U855 ( .A1(n848), .A2(G567), .ZN(n778) );
  XOR2_X1 U856 ( .A(KEYINPUT11), .B(n778), .Z(G234) );
  XNOR2_X1 U857 ( .A(G860), .B(KEYINPUT75), .ZN(n785) );
  OR2_X1 U858 ( .A1(n966), .A2(n785), .ZN(G153) );
  NAND2_X1 U859 ( .A1(G868), .A2(G301), .ZN(n780) );
  INV_X1 U860 ( .A(G868), .ZN(n818) );
  NAND2_X1 U861 ( .A1(n953), .A2(n818), .ZN(n779) );
  NAND2_X1 U862 ( .A1(n780), .A2(n779), .ZN(G284) );
  NOR2_X1 U863 ( .A1(G868), .A2(G299), .ZN(n781) );
  XOR2_X1 U864 ( .A(KEYINPUT79), .B(n781), .Z(n784) );
  NOR2_X1 U865 ( .A1(G286), .A2(n818), .ZN(n782) );
  XNOR2_X1 U866 ( .A(KEYINPUT78), .B(n782), .ZN(n783) );
  NOR2_X1 U867 ( .A1(n784), .A2(n783), .ZN(G297) );
  NAND2_X1 U868 ( .A1(n785), .A2(G559), .ZN(n786) );
  INV_X1 U869 ( .A(n953), .ZN(n791) );
  NAND2_X1 U870 ( .A1(n786), .A2(n791), .ZN(n787) );
  XNOR2_X1 U871 ( .A(n787), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U872 ( .A1(n966), .A2(G868), .ZN(n790) );
  NAND2_X1 U873 ( .A1(G868), .A2(n791), .ZN(n788) );
  NOR2_X1 U874 ( .A1(G559), .A2(n788), .ZN(n789) );
  NOR2_X1 U875 ( .A1(n790), .A2(n789), .ZN(G282) );
  NAND2_X1 U876 ( .A1(n791), .A2(G559), .ZN(n815) );
  XNOR2_X1 U877 ( .A(n966), .B(n815), .ZN(n792) );
  NOR2_X1 U878 ( .A1(G860), .A2(n792), .ZN(n793) );
  XNOR2_X1 U879 ( .A(n793), .B(KEYINPUT81), .ZN(n805) );
  NAND2_X1 U880 ( .A1(G80), .A2(n794), .ZN(n795) );
  XNOR2_X1 U881 ( .A(n795), .B(KEYINPUT82), .ZN(n798) );
  NAND2_X1 U882 ( .A1(n796), .A2(G93), .ZN(n797) );
  NAND2_X1 U883 ( .A1(n798), .A2(n797), .ZN(n804) );
  NAND2_X1 U884 ( .A1(G55), .A2(n799), .ZN(n802) );
  NAND2_X1 U885 ( .A1(G67), .A2(n800), .ZN(n801) );
  NAND2_X1 U886 ( .A1(n802), .A2(n801), .ZN(n803) );
  NOR2_X1 U887 ( .A1(n804), .A2(n803), .ZN(n817) );
  XOR2_X1 U888 ( .A(n805), .B(n817), .Z(G145) );
  XNOR2_X1 U889 ( .A(G288), .B(G290), .ZN(n814) );
  XNOR2_X1 U890 ( .A(n966), .B(n817), .ZN(n810) );
  XOR2_X1 U891 ( .A(KEYINPUT89), .B(KEYINPUT90), .Z(n808) );
  XNOR2_X1 U892 ( .A(n806), .B(KEYINPUT19), .ZN(n807) );
  XNOR2_X1 U893 ( .A(n808), .B(n807), .ZN(n809) );
  XNOR2_X1 U894 ( .A(n810), .B(n809), .ZN(n811) );
  XNOR2_X1 U895 ( .A(G303), .B(n811), .ZN(n812) );
  XNOR2_X1 U896 ( .A(n812), .B(G305), .ZN(n813) );
  XNOR2_X1 U897 ( .A(n814), .B(n813), .ZN(n915) );
  XOR2_X1 U898 ( .A(n915), .B(n815), .Z(n816) );
  NOR2_X1 U899 ( .A1(n818), .A2(n816), .ZN(n820) );
  AND2_X1 U900 ( .A1(n818), .A2(n817), .ZN(n819) );
  NOR2_X1 U901 ( .A1(n820), .A2(n819), .ZN(G295) );
  NAND2_X1 U902 ( .A1(G2078), .A2(G2084), .ZN(n821) );
  XNOR2_X1 U903 ( .A(n821), .B(KEYINPUT20), .ZN(n822) );
  XNOR2_X1 U904 ( .A(n822), .B(KEYINPUT91), .ZN(n823) );
  NAND2_X1 U905 ( .A1(n823), .A2(G2090), .ZN(n824) );
  XNOR2_X1 U906 ( .A(KEYINPUT21), .B(n824), .ZN(n825) );
  NAND2_X1 U907 ( .A1(n825), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U908 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U909 ( .A(KEYINPUT72), .B(G57), .Z(G237) );
  NAND2_X1 U910 ( .A1(G132), .A2(G82), .ZN(n826) );
  XNOR2_X1 U911 ( .A(n826), .B(KEYINPUT92), .ZN(n827) );
  XNOR2_X1 U912 ( .A(n827), .B(KEYINPUT22), .ZN(n828) );
  NOR2_X1 U913 ( .A1(G218), .A2(n828), .ZN(n829) );
  NAND2_X1 U914 ( .A1(G96), .A2(n829), .ZN(n853) );
  NAND2_X1 U915 ( .A1(G2106), .A2(n853), .ZN(n833) );
  NAND2_X1 U916 ( .A1(G120), .A2(G69), .ZN(n830) );
  NOR2_X1 U917 ( .A1(G237), .A2(n830), .ZN(n831) );
  NAND2_X1 U918 ( .A1(G108), .A2(n831), .ZN(n854) );
  NAND2_X1 U919 ( .A1(G567), .A2(n854), .ZN(n832) );
  NAND2_X1 U920 ( .A1(n833), .A2(n832), .ZN(n834) );
  XNOR2_X1 U921 ( .A(KEYINPUT93), .B(n834), .ZN(G319) );
  INV_X1 U922 ( .A(G319), .ZN(n836) );
  NAND2_X1 U923 ( .A1(G661), .A2(G483), .ZN(n835) );
  NOR2_X1 U924 ( .A1(n836), .A2(n835), .ZN(n852) );
  NAND2_X1 U925 ( .A1(n852), .A2(G36), .ZN(G176) );
  XNOR2_X1 U926 ( .A(G2443), .B(G2451), .ZN(n846) );
  XOR2_X1 U927 ( .A(G2446), .B(G2430), .Z(n838) );
  XNOR2_X1 U928 ( .A(KEYINPUT109), .B(G2438), .ZN(n837) );
  XNOR2_X1 U929 ( .A(n838), .B(n837), .ZN(n842) );
  XOR2_X1 U930 ( .A(G2435), .B(G2454), .Z(n840) );
  XNOR2_X1 U931 ( .A(G1341), .B(G1348), .ZN(n839) );
  XNOR2_X1 U932 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U933 ( .A(n842), .B(n841), .Z(n844) );
  XNOR2_X1 U934 ( .A(G2427), .B(KEYINPUT108), .ZN(n843) );
  XNOR2_X1 U935 ( .A(n844), .B(n843), .ZN(n845) );
  XNOR2_X1 U936 ( .A(n846), .B(n845), .ZN(n847) );
  NAND2_X1 U937 ( .A1(n847), .A2(G14), .ZN(n919) );
  XOR2_X1 U938 ( .A(KEYINPUT110), .B(n919), .Z(G401) );
  NAND2_X1 U939 ( .A1(n848), .A2(G2106), .ZN(n849) );
  XOR2_X1 U940 ( .A(KEYINPUT111), .B(n849), .Z(G217) );
  AND2_X1 U941 ( .A1(G15), .A2(G2), .ZN(n850) );
  NAND2_X1 U942 ( .A1(G661), .A2(n850), .ZN(G259) );
  NAND2_X1 U943 ( .A1(G3), .A2(G1), .ZN(n851) );
  NAND2_X1 U944 ( .A1(n852), .A2(n851), .ZN(G188) );
  XOR2_X1 U945 ( .A(G69), .B(KEYINPUT112), .Z(G235) );
  INV_X1 U947 ( .A(G132), .ZN(G219) );
  INV_X1 U948 ( .A(G120), .ZN(G236) );
  INV_X1 U949 ( .A(G108), .ZN(G238) );
  INV_X1 U950 ( .A(G82), .ZN(G220) );
  NOR2_X1 U951 ( .A1(n854), .A2(n853), .ZN(G325) );
  INV_X1 U952 ( .A(G325), .ZN(G261) );
  XOR2_X1 U953 ( .A(G2100), .B(G2096), .Z(n856) );
  XNOR2_X1 U954 ( .A(KEYINPUT42), .B(G2678), .ZN(n855) );
  XNOR2_X1 U955 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U956 ( .A(KEYINPUT43), .B(G2090), .Z(n858) );
  XNOR2_X1 U957 ( .A(G2067), .B(G2072), .ZN(n857) );
  XNOR2_X1 U958 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U959 ( .A(n860), .B(n859), .Z(n862) );
  XNOR2_X1 U960 ( .A(G2078), .B(G2084), .ZN(n861) );
  XNOR2_X1 U961 ( .A(n862), .B(n861), .ZN(G227) );
  XOR2_X1 U962 ( .A(G1976), .B(G1971), .Z(n864) );
  XNOR2_X1 U963 ( .A(G1966), .B(G1961), .ZN(n863) );
  XNOR2_X1 U964 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U965 ( .A(n865), .B(G2474), .Z(n867) );
  XNOR2_X1 U966 ( .A(G1991), .B(G1996), .ZN(n866) );
  XNOR2_X1 U967 ( .A(n867), .B(n866), .ZN(n871) );
  XOR2_X1 U968 ( .A(KEYINPUT41), .B(G1986), .Z(n869) );
  XNOR2_X1 U969 ( .A(G1956), .B(G1981), .ZN(n868) );
  XNOR2_X1 U970 ( .A(n869), .B(n868), .ZN(n870) );
  XNOR2_X1 U971 ( .A(n871), .B(n870), .ZN(G229) );
  NAND2_X1 U972 ( .A1(G100), .A2(n897), .ZN(n873) );
  NAND2_X1 U973 ( .A1(G112), .A2(n902), .ZN(n872) );
  NAND2_X1 U974 ( .A1(n873), .A2(n872), .ZN(n881) );
  NAND2_X1 U975 ( .A1(G136), .A2(n898), .ZN(n874) );
  XNOR2_X1 U976 ( .A(KEYINPUT114), .B(n874), .ZN(n878) );
  XOR2_X1 U977 ( .A(KEYINPUT113), .B(KEYINPUT44), .Z(n876) );
  NAND2_X1 U978 ( .A1(G124), .A2(n901), .ZN(n875) );
  XNOR2_X1 U979 ( .A(n876), .B(n875), .ZN(n877) );
  NAND2_X1 U980 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U981 ( .A(KEYINPUT115), .B(n879), .Z(n880) );
  NOR2_X1 U982 ( .A1(n881), .A2(n880), .ZN(G162) );
  NAND2_X1 U983 ( .A1(G106), .A2(n897), .ZN(n883) );
  NAND2_X1 U984 ( .A1(G142), .A2(n898), .ZN(n882) );
  NAND2_X1 U985 ( .A1(n883), .A2(n882), .ZN(n884) );
  XNOR2_X1 U986 ( .A(n884), .B(KEYINPUT45), .ZN(n889) );
  NAND2_X1 U987 ( .A1(G130), .A2(n901), .ZN(n886) );
  NAND2_X1 U988 ( .A1(G118), .A2(n902), .ZN(n885) );
  NAND2_X1 U989 ( .A1(n886), .A2(n885), .ZN(n887) );
  XOR2_X1 U990 ( .A(KEYINPUT116), .B(n887), .Z(n888) );
  NAND2_X1 U991 ( .A1(n889), .A2(n888), .ZN(n890) );
  XNOR2_X1 U992 ( .A(n890), .B(G164), .ZN(n891) );
  XNOR2_X1 U993 ( .A(G162), .B(n891), .ZN(n911) );
  XOR2_X1 U994 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n895) );
  XOR2_X1 U995 ( .A(n893), .B(n892), .Z(n894) );
  XNOR2_X1 U996 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U997 ( .A(n927), .B(n896), .ZN(n909) );
  NAND2_X1 U998 ( .A1(G103), .A2(n897), .ZN(n900) );
  NAND2_X1 U999 ( .A1(G139), .A2(n898), .ZN(n899) );
  NAND2_X1 U1000 ( .A1(n900), .A2(n899), .ZN(n907) );
  NAND2_X1 U1001 ( .A1(G127), .A2(n901), .ZN(n904) );
  NAND2_X1 U1002 ( .A1(G115), .A2(n902), .ZN(n903) );
  NAND2_X1 U1003 ( .A1(n904), .A2(n903), .ZN(n905) );
  XOR2_X1 U1004 ( .A(KEYINPUT47), .B(n905), .Z(n906) );
  NOR2_X1 U1005 ( .A1(n907), .A2(n906), .ZN(n934) );
  XNOR2_X1 U1006 ( .A(G160), .B(n934), .ZN(n908) );
  XNOR2_X1 U1007 ( .A(n909), .B(n908), .ZN(n910) );
  XNOR2_X1 U1008 ( .A(n911), .B(n910), .ZN(n913) );
  XOR2_X1 U1009 ( .A(n913), .B(n912), .Z(n914) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n914), .ZN(G395) );
  XNOR2_X1 U1011 ( .A(G286), .B(n953), .ZN(n916) );
  XNOR2_X1 U1012 ( .A(n916), .B(n915), .ZN(n917) );
  XNOR2_X1 U1013 ( .A(n917), .B(G301), .ZN(n918) );
  NOR2_X1 U1014 ( .A1(G37), .A2(n918), .ZN(G397) );
  NAND2_X1 U1015 ( .A1(G319), .A2(n919), .ZN(n922) );
  NOR2_X1 U1016 ( .A1(G227), .A2(G229), .ZN(n920) );
  XNOR2_X1 U1017 ( .A(KEYINPUT49), .B(n920), .ZN(n921) );
  NOR2_X1 U1018 ( .A1(n922), .A2(n921), .ZN(n924) );
  NOR2_X1 U1019 ( .A1(G395), .A2(G397), .ZN(n923) );
  NAND2_X1 U1020 ( .A1(n924), .A2(n923), .ZN(G225) );
  INV_X1 U1021 ( .A(G225), .ZN(G308) );
  INV_X1 U1022 ( .A(G96), .ZN(G221) );
  NAND2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(n947) );
  XNOR2_X1 U1024 ( .A(G160), .B(G2084), .ZN(n928) );
  NAND2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n929) );
  NOR2_X1 U1026 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1027 ( .A(KEYINPUT117), .B(n931), .ZN(n932) );
  NOR2_X1 U1028 ( .A1(n933), .A2(n932), .ZN(n945) );
  XOR2_X1 U1029 ( .A(G2072), .B(n934), .Z(n936) );
  XOR2_X1 U1030 ( .A(G164), .B(G2078), .Z(n935) );
  NOR2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1032 ( .A(KEYINPUT50), .B(n937), .Z(n943) );
  XOR2_X1 U1033 ( .A(G2090), .B(G162), .Z(n938) );
  NOR2_X1 U1034 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1035 ( .A(KEYINPUT51), .B(n940), .Z(n941) );
  XOR2_X1 U1036 ( .A(KEYINPUT118), .B(n941), .Z(n942) );
  NOR2_X1 U1037 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1038 ( .A1(n945), .A2(n944), .ZN(n946) );
  NOR2_X1 U1039 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1040 ( .A(KEYINPUT119), .B(n948), .Z(n949) );
  XNOR2_X1 U1041 ( .A(KEYINPUT52), .B(n949), .ZN(n950) );
  XOR2_X1 U1042 ( .A(KEYINPUT55), .B(KEYINPUT120), .Z(n996) );
  NAND2_X1 U1043 ( .A1(n950), .A2(n996), .ZN(n951) );
  NAND2_X1 U1044 ( .A1(n951), .A2(G29), .ZN(n978) );
  XOR2_X1 U1045 ( .A(G16), .B(KEYINPUT56), .Z(n952) );
  XNOR2_X1 U1046 ( .A(KEYINPUT123), .B(n952), .ZN(n976) );
  XNOR2_X1 U1047 ( .A(G299), .B(G1956), .ZN(n955) );
  XNOR2_X1 U1048 ( .A(n953), .B(G1348), .ZN(n954) );
  NOR2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n957) );
  NAND2_X1 U1050 ( .A1(n957), .A2(n956), .ZN(n958) );
  NOR2_X1 U1051 ( .A1(n959), .A2(n958), .ZN(n965) );
  XOR2_X1 U1052 ( .A(G1966), .B(G168), .Z(n960) );
  XNOR2_X1 U1053 ( .A(KEYINPUT124), .B(n960), .ZN(n961) );
  NOR2_X1 U1054 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1055 ( .A(KEYINPUT57), .B(n963), .Z(n964) );
  NAND2_X1 U1056 ( .A1(n965), .A2(n964), .ZN(n968) );
  XNOR2_X1 U1057 ( .A(n966), .B(G1341), .ZN(n967) );
  NOR2_X1 U1058 ( .A1(n968), .A2(n967), .ZN(n974) );
  XNOR2_X1 U1059 ( .A(G171), .B(G1961), .ZN(n970) );
  NAND2_X1 U1060 ( .A1(G1971), .A2(G303), .ZN(n969) );
  NAND2_X1 U1061 ( .A1(n970), .A2(n969), .ZN(n971) );
  NOR2_X1 U1062 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1063 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1064 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1065 ( .A1(n978), .A2(n977), .ZN(n1003) );
  XOR2_X1 U1066 ( .A(G2067), .B(G26), .Z(n979) );
  NAND2_X1 U1067 ( .A1(n979), .A2(G28), .ZN(n988) );
  XNOR2_X1 U1068 ( .A(G1996), .B(G32), .ZN(n981) );
  XNOR2_X1 U1069 ( .A(G33), .B(G2072), .ZN(n980) );
  NOR2_X1 U1070 ( .A1(n981), .A2(n980), .ZN(n986) );
  XNOR2_X1 U1071 ( .A(G1991), .B(G25), .ZN(n984) );
  XNOR2_X1 U1072 ( .A(G27), .B(n982), .ZN(n983) );
  NOR2_X1 U1073 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1074 ( .A1(n986), .A2(n985), .ZN(n987) );
  NOR2_X1 U1075 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1076 ( .A(n989), .B(KEYINPUT121), .ZN(n990) );
  XNOR2_X1 U1077 ( .A(n990), .B(KEYINPUT53), .ZN(n993) );
  XOR2_X1 U1078 ( .A(G2084), .B(KEYINPUT54), .Z(n991) );
  XNOR2_X1 U1079 ( .A(G34), .B(n991), .ZN(n992) );
  NAND2_X1 U1080 ( .A1(n993), .A2(n992), .ZN(n995) );
  XNOR2_X1 U1081 ( .A(G35), .B(G2090), .ZN(n994) );
  NOR2_X1 U1082 ( .A1(n995), .A2(n994), .ZN(n997) );
  XOR2_X1 U1083 ( .A(n997), .B(n996), .Z(n999) );
  INV_X1 U1084 ( .A(G29), .ZN(n998) );
  NAND2_X1 U1085 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1086 ( .A1(G11), .A2(n1000), .ZN(n1001) );
  XNOR2_X1 U1087 ( .A(KEYINPUT122), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1088 ( .A1(n1003), .A2(n1002), .ZN(n1028) );
  XNOR2_X1 U1089 ( .A(G1966), .B(G21), .ZN(n1005) );
  XNOR2_X1 U1090 ( .A(G5), .B(G1961), .ZN(n1004) );
  NOR2_X1 U1091 ( .A1(n1005), .A2(n1004), .ZN(n1016) );
  XNOR2_X1 U1092 ( .A(KEYINPUT59), .B(G1348), .ZN(n1006) );
  XNOR2_X1 U1093 ( .A(n1006), .B(G4), .ZN(n1013) );
  XNOR2_X1 U1094 ( .A(G1956), .B(G20), .ZN(n1011) );
  XNOR2_X1 U1095 ( .A(G1341), .B(G19), .ZN(n1008) );
  XNOR2_X1 U1096 ( .A(G1981), .B(G6), .ZN(n1007) );
  NOR2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1098 ( .A(KEYINPUT125), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XOR2_X1 U1101 ( .A(KEYINPUT60), .B(n1014), .Z(n1015) );
  NAND2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1023) );
  XNOR2_X1 U1103 ( .A(G1971), .B(G22), .ZN(n1018) );
  XNOR2_X1 U1104 ( .A(G24), .B(G1986), .ZN(n1017) );
  NOR2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1020) );
  XOR2_X1 U1106 ( .A(G1976), .B(G23), .Z(n1019) );
  NAND2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1108 ( .A(KEYINPUT58), .B(n1021), .ZN(n1022) );
  NOR2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1110 ( .A(KEYINPUT61), .B(n1024), .Z(n1025) );
  NOR2_X1 U1111 ( .A1(G16), .A2(n1025), .ZN(n1026) );
  XOR2_X1 U1112 ( .A(KEYINPUT126), .B(n1026), .Z(n1027) );
  NAND2_X1 U1113 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1114 ( .A(n1029), .B(KEYINPUT127), .ZN(n1030) );
  XNOR2_X1 U1115 ( .A(KEYINPUT62), .B(n1030), .ZN(G311) );
  INV_X1 U1116 ( .A(G311), .ZN(G150) );
  INV_X1 U1117 ( .A(G303), .ZN(G166) );
endmodule

