//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 1 1 1 1 0 1 0 1 0 0 1 1 1 1 0 0 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 1 1 0 0 1 0 1 0 1 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n832, new_n834, new_n835,
    new_n836, new_n838, new_n839, new_n840, new_n841, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951;
  INV_X1    g000(.A(KEYINPUT81), .ZN(new_n202));
  INV_X1    g001(.A(G228gat), .ZN(new_n203));
  INV_X1    g002(.A(G233gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G211gat), .ZN(new_n206));
  OR2_X1    g005(.A1(KEYINPUT74), .A2(G218gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(KEYINPUT74), .A2(G218gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT22), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(G197gat), .B(G204gat), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n206), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n212), .A2(KEYINPUT22), .A3(new_n206), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(G218gat), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n212), .ZN(new_n217));
  AOI21_X1  g016(.A(KEYINPUT22), .B1(new_n207), .B2(new_n208), .ZN(new_n218));
  OAI21_X1  g017(.A(G211gat), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G218gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n219), .A2(new_n220), .A3(new_n214), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n216), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT80), .ZN(new_n223));
  NOR2_X1   g022(.A1(G155gat), .A2(G162gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT2), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(G155gat), .A2(G162gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G148gat), .ZN(new_n229));
  OR2_X1    g028(.A1(KEYINPUT78), .A2(G141gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(KEYINPUT78), .A2(G141gat), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n229), .A2(G141gat), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n228), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  AND3_X1   g034(.A1(KEYINPUT77), .A2(G155gat), .A3(G162gat), .ZN(new_n236));
  AOI21_X1  g035(.A(KEYINPUT77), .B1(G155gat), .B2(G162gat), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n224), .ZN(new_n239));
  XNOR2_X1  g038(.A(G141gat), .B(G148gat), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT77), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n241), .A2(new_n225), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n238), .B(new_n239), .C1(new_n240), .C2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n235), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT29), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n222), .A2(new_n223), .A3(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n223), .B1(new_n222), .B2(new_n247), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n205), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n244), .B1(new_n222), .B2(KEYINPUT29), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n243), .ZN(new_n252));
  AND2_X1   g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n202), .B1(new_n250), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n222), .A2(new_n247), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  OAI22_X1  g055(.A1(new_n253), .A2(new_n256), .B1(new_n203), .B2(new_n204), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n255), .A2(KEYINPUT80), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n222), .A2(new_n223), .A3(new_n247), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n251), .A2(new_n252), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n260), .A2(KEYINPUT81), .A3(new_n205), .A4(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n254), .A2(new_n257), .A3(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G78gat), .B(G106gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n264), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n254), .A2(new_n257), .A3(new_n266), .A4(new_n262), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(KEYINPUT79), .B(KEYINPUT31), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n269), .B(G50gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(G22gat), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n265), .A2(new_n271), .A3(new_n267), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT72), .ZN(new_n276));
  XNOR2_X1  g075(.A(G113gat), .B(G120gat), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT1), .ZN(new_n279));
  XNOR2_X1  g078(.A(G127gat), .B(G134gat), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  XOR2_X1   g080(.A(G127gat), .B(G134gat), .Z(new_n282));
  OAI21_X1  g081(.A(new_n282), .B1(KEYINPUT1), .B2(new_n277), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(G190gat), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT70), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n286), .A2(G183gat), .ZN(new_n287));
  INV_X1    g086(.A(G183gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n288), .A2(KEYINPUT70), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n285), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT69), .ZN(new_n291));
  NAND2_X1  g090(.A1(G183gat), .A2(G190gat), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT68), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT24), .ZN(new_n295));
  NAND3_X1  g094(.A1(KEYINPUT68), .A2(G183gat), .A3(G190gat), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n290), .A2(new_n291), .A3(new_n297), .A4(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT25), .ZN(new_n300));
  NAND2_X1  g099(.A1(G169gat), .A2(G176gat), .ZN(new_n301));
  OR2_X1    g100(.A1(new_n301), .A2(KEYINPUT66), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(KEYINPUT66), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n300), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NOR2_X1   g103(.A1(G169gat), .A2(G176gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n305), .A2(KEYINPUT23), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT67), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g107(.A(KEYINPUT67), .B1(G169gat), .B2(G176gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n306), .B1(new_n310), .B2(KEYINPUT23), .ZN(new_n311));
  AND3_X1   g110(.A1(new_n299), .A2(new_n304), .A3(new_n311), .ZN(new_n312));
  OR2_X1    g111(.A1(new_n298), .A2(new_n291), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT65), .ZN(new_n314));
  INV_X1    g113(.A(G169gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT23), .ZN(new_n316));
  INV_X1    g115(.A(G176gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(KEYINPUT64), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT64), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G176gat), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n316), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n301), .B1(new_n305), .B2(KEYINPUT23), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n314), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT23), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n324), .A2(G169gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n319), .A2(G176gat), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n317), .A2(KEYINPUT64), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n325), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AND2_X1   g127(.A1(G169gat), .A2(G176gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n315), .A2(new_n317), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n329), .B1(new_n330), .B2(new_n324), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n328), .A2(KEYINPUT65), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n292), .A2(new_n295), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n333), .B(new_n298), .C1(G183gat), .C2(G190gat), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n323), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  AOI22_X1  g134(.A1(new_n312), .A2(new_n313), .B1(new_n300), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n288), .A2(KEYINPUT70), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n286), .A2(G183gat), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(new_n338), .A3(KEYINPUT27), .ZN(new_n339));
  OR2_X1    g138(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n340));
  AOI211_X1 g139(.A(KEYINPUT28), .B(G190gat), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT26), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n301), .B1(new_n305), .B2(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n343), .B1(new_n310), .B2(new_n342), .ZN(new_n344));
  NAND2_X1  g143(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n345));
  AOI21_X1  g144(.A(G190gat), .B1(new_n340), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT28), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n292), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NOR3_X1   g147(.A1(new_n341), .A2(new_n344), .A3(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n284), .B1(new_n336), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n335), .A2(new_n300), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n299), .A2(new_n311), .A3(new_n313), .A4(new_n304), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n349), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n353), .A2(new_n281), .A3(new_n283), .A4(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(G227gat), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n356), .A2(new_n204), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n350), .A2(new_n355), .A3(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n359), .B(KEYINPUT34), .ZN(new_n360));
  XNOR2_X1  g159(.A(G15gat), .B(G43gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n361), .B(G71gat), .ZN(new_n362));
  XOR2_X1   g161(.A(KEYINPUT71), .B(G99gat), .Z(new_n363));
  XNOR2_X1  g162(.A(new_n362), .B(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n358), .B1(new_n350), .B2(new_n355), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n364), .B1(new_n365), .B2(KEYINPUT33), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT32), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n350), .A2(new_n355), .ZN(new_n370));
  AOI221_X4 g169(.A(new_n367), .B1(KEYINPUT33), .B2(new_n364), .C1(new_n370), .C2(new_n357), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n276), .B(new_n360), .C1(new_n369), .C2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n360), .B1(new_n369), .B2(new_n371), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n370), .A2(new_n357), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(KEYINPUT32), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT33), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n375), .A2(new_n377), .A3(new_n364), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT34), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n359), .B(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n366), .A2(new_n368), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n378), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n373), .A2(new_n382), .A3(KEYINPUT72), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n275), .B1(new_n372), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT35), .ZN(new_n385));
  XOR2_X1   g184(.A(KEYINPUT76), .B(G92gat), .Z(new_n386));
  XNOR2_X1  g185(.A(G8gat), .B(G36gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n386), .B(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(KEYINPUT75), .B(G64gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n388), .B(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(G226gat), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n392), .A2(new_n204), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n349), .B1(new_n351), .B2(new_n352), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n394), .B1(new_n395), .B2(KEYINPUT29), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n393), .B1(new_n336), .B2(new_n349), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n396), .A2(new_n222), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n222), .B1(new_n396), .B2(new_n397), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n391), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n222), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n353), .A2(new_n354), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n393), .B1(new_n402), .B2(new_n246), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n395), .A2(new_n394), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n401), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n396), .A2(new_n222), .A3(new_n397), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n405), .A2(new_n406), .A3(new_n390), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n400), .A2(new_n407), .A3(KEYINPUT30), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT30), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n409), .B(new_n391), .C1(new_n398), .C2(new_n399), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n235), .A2(new_n243), .A3(new_n281), .A4(new_n283), .ZN(new_n412));
  NAND2_X1  g211(.A1(G225gat), .A2(G233gat), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(G141gat), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(G148gat), .ZN(new_n417));
  AOI22_X1  g216(.A1(new_n233), .A2(new_n417), .B1(KEYINPUT77), .B2(KEYINPUT2), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n227), .A2(new_n241), .ZN(new_n419));
  NAND3_X1  g218(.A1(KEYINPUT77), .A2(G155gat), .A3(G162gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NOR3_X1   g220(.A1(new_n418), .A2(new_n421), .A3(new_n224), .ZN(new_n422));
  INV_X1    g221(.A(new_n231), .ZN(new_n423));
  NOR2_X1   g222(.A1(KEYINPUT78), .A2(G141gat), .ZN(new_n424));
  OAI21_X1  g223(.A(G148gat), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AOI22_X1  g224(.A1(new_n425), .A2(new_n233), .B1(new_n227), .B2(new_n226), .ZN(new_n426));
  OAI21_X1  g225(.A(KEYINPUT3), .B1(new_n422), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n427), .A2(new_n284), .A3(new_n245), .ZN(new_n428));
  AND2_X1   g227(.A1(new_n412), .A2(KEYINPUT4), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n412), .A2(KEYINPUT4), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n415), .B(new_n428), .C1(new_n429), .C2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT5), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n252), .A2(new_n284), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(new_n412), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n432), .B1(new_n434), .B2(new_n414), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n414), .A2(KEYINPUT5), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n428), .B(new_n437), .C1(new_n429), .C2(new_n430), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  XNOR2_X1  g238(.A(KEYINPUT0), .B(G57gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n440), .B(G85gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(G1gat), .B(G29gat), .ZN(new_n442));
  XOR2_X1   g241(.A(new_n441), .B(new_n442), .Z(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n439), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n436), .A2(new_n443), .A3(new_n438), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT6), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT83), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n439), .A2(KEYINPUT6), .A3(new_n444), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n445), .A2(new_n446), .A3(KEYINPUT83), .A4(new_n447), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n384), .A2(new_n385), .A3(new_n411), .A4(new_n453), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n273), .A2(new_n373), .A3(new_n382), .A4(new_n274), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n448), .A2(new_n451), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n411), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(KEYINPUT35), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n273), .A2(new_n274), .ZN(new_n459));
  OAI21_X1  g258(.A(KEYINPUT37), .B1(new_n398), .B2(new_n399), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT37), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n405), .A2(new_n461), .A3(new_n406), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n391), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT38), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n400), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AOI211_X1 g264(.A(KEYINPUT38), .B(new_n391), .C1(new_n460), .C2(new_n462), .ZN(new_n466));
  NOR3_X1   g265(.A1(new_n465), .A2(new_n453), .A3(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT82), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT40), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n408), .A2(new_n445), .A3(new_n410), .A4(new_n470), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n468), .A2(new_n469), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n428), .B1(new_n429), .B2(new_n430), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(new_n414), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n474), .A2(KEYINPUT39), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n475), .A2(new_n444), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n474), .B(KEYINPUT39), .C1(new_n414), .C2(new_n434), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n472), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AND3_X1   g277(.A1(new_n476), .A2(new_n472), .A3(new_n477), .ZN(new_n479));
  NOR3_X1   g278(.A1(new_n471), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n459), .B1(new_n467), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n275), .A2(new_n456), .A3(new_n411), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT36), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n383), .A2(new_n484), .A3(new_n372), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT73), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n373), .A2(new_n382), .A3(KEYINPUT36), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n383), .A2(KEYINPUT73), .A3(new_n484), .A4(new_n372), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  AOI22_X1  g289(.A1(new_n454), .A2(new_n458), .B1(new_n483), .B2(new_n490), .ZN(new_n491));
  AND3_X1   g290(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n492));
  AND2_X1   g291(.A1(KEYINPUT93), .A2(KEYINPUT7), .ZN(new_n493));
  NOR2_X1   g292(.A1(KEYINPUT93), .A2(KEYINPUT7), .ZN(new_n494));
  OAI211_X1 g293(.A(G85gat), .B(G92gat), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  OR2_X1    g294(.A1(new_n495), .A2(KEYINPUT94), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(KEYINPUT94), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT7), .ZN(new_n498));
  NAND2_X1  g297(.A1(G85gat), .A2(G92gat), .ZN(new_n499));
  XOR2_X1   g298(.A(new_n499), .B(KEYINPUT92), .Z(new_n500));
  OAI211_X1 g299(.A(new_n496), .B(new_n497), .C1(new_n498), .C2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(G99gat), .A2(G106gat), .ZN(new_n502));
  INV_X1    g301(.A(G85gat), .ZN(new_n503));
  INV_X1    g302(.A(G92gat), .ZN(new_n504));
  AOI22_X1  g303(.A1(KEYINPUT8), .A2(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  XOR2_X1   g305(.A(G99gat), .B(G106gat), .Z(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n507), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n501), .A2(new_n509), .A3(new_n505), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(G50gat), .ZN(new_n512));
  OAI21_X1  g311(.A(KEYINPUT15), .B1(new_n512), .B2(G43gat), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n513), .B1(G43gat), .B2(new_n512), .ZN(new_n514));
  OR2_X1    g313(.A1(new_n512), .A2(G43gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(KEYINPUT85), .B(G43gat), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n515), .B1(new_n516), .B2(G50gat), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT15), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n514), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g318(.A1(G29gat), .A2(G36gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n520), .B(KEYINPUT14), .ZN(new_n521));
  OR2_X1    g320(.A1(new_n521), .A2(KEYINPUT86), .ZN(new_n522));
  NAND2_X1  g321(.A1(G29gat), .A2(G36gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(KEYINPUT86), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n519), .A2(new_n522), .A3(new_n523), .A4(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n521), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(new_n523), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(new_n514), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n492), .B1(new_n511), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n508), .A2(new_n510), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT95), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT17), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n529), .B(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n530), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  XOR2_X1   g335(.A(G190gat), .B(G218gat), .Z(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  OAI211_X1 g338(.A(new_n537), .B(new_n530), .C1(new_n533), .C2(new_n535), .ZN(new_n540));
  XNOR2_X1  g339(.A(G134gat), .B(G162gat), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n539), .A2(KEYINPUT96), .A3(new_n540), .A4(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT96), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n540), .A2(new_n546), .ZN(new_n547));
  AOI22_X1  g346(.A1(new_n547), .A2(new_n543), .B1(new_n539), .B2(new_n540), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G15gat), .B(G22gat), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT16), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n550), .B1(new_n551), .B2(G1gat), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n552), .B1(G1gat), .B2(new_n550), .ZN(new_n553));
  XOR2_X1   g352(.A(new_n553), .B(G8gat), .Z(new_n554));
  XNOR2_X1  g353(.A(G57gat), .B(G64gat), .ZN(new_n555));
  AOI21_X1  g354(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n556));
  OR2_X1    g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  XOR2_X1   g356(.A(G71gat), .B(G78gat), .Z(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  XOR2_X1   g358(.A(new_n559), .B(KEYINPUT90), .Z(new_n560));
  INV_X1    g359(.A(KEYINPUT21), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n554), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(new_n206), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n559), .A2(new_n561), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT88), .B(KEYINPUT20), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  AND2_X1   g367(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n565), .A2(new_n568), .ZN(new_n570));
  XNOR2_X1  g369(.A(G127gat), .B(G155gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(G231gat), .A2(G233gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(KEYINPUT91), .B(G183gat), .ZN(new_n574));
  XOR2_X1   g373(.A(new_n573), .B(new_n574), .Z(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NOR3_X1   g375(.A1(new_n569), .A2(new_n570), .A3(new_n576), .ZN(new_n577));
  OR2_X1    g376(.A1(new_n565), .A2(new_n568), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n565), .A2(new_n568), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n575), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n549), .B1(new_n577), .B2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n554), .ZN(new_n582));
  OR2_X1    g381(.A1(new_n535), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n529), .ZN(new_n584));
  NAND2_X1  g383(.A1(G229gat), .A2(G233gat), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT18), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n586), .A2(KEYINPUT87), .A3(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(new_n554), .B(new_n529), .Z(new_n589));
  XOR2_X1   g388(.A(new_n585), .B(KEYINPUT13), .Z(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n587), .A2(KEYINPUT87), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n583), .A2(new_n584), .A3(new_n585), .A4(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n588), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G113gat), .B(G141gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G169gat), .B(G197gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  XOR2_X1   g398(.A(new_n599), .B(KEYINPUT12), .Z(new_n600));
  NAND2_X1  g399(.A1(new_n594), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n600), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n588), .A2(new_n591), .A3(new_n593), .A4(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT99), .ZN(new_n606));
  INV_X1    g405(.A(G230gat), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n607), .A2(new_n204), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n511), .A2(new_n559), .ZN(new_n609));
  INV_X1    g408(.A(new_n559), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n531), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT10), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NOR3_X1   g413(.A1(new_n560), .A2(new_n531), .A3(new_n613), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n608), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  NOR3_X1   g416(.A1(new_n612), .A2(new_n607), .A3(new_n204), .ZN(new_n618));
  XOR2_X1   g417(.A(KEYINPUT98), .B(G204gat), .Z(new_n619));
  XNOR2_X1  g418(.A(G120gat), .B(G148gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(KEYINPUT97), .B(G176gat), .ZN(new_n622));
  XOR2_X1   g421(.A(new_n621), .B(new_n622), .Z(new_n623));
  NOR3_X1   g422(.A1(new_n617), .A2(new_n618), .A3(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n623), .ZN(new_n625));
  INV_X1    g424(.A(new_n618), .ZN(new_n626));
  AOI21_X1  g425(.A(KEYINPUT10), .B1(new_n609), .B2(new_n611), .ZN(new_n627));
  OAI22_X1  g426(.A1(new_n627), .A2(new_n615), .B1(new_n607), .B2(new_n204), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n625), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n606), .B1(new_n624), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n623), .B1(new_n617), .B2(new_n618), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n626), .A2(new_n628), .A3(new_n625), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n631), .A2(KEYINPUT99), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n605), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NOR3_X1   g435(.A1(new_n491), .A2(new_n581), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n456), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(G1gat), .ZN(G1324gat));
  INV_X1    g439(.A(new_n411), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(KEYINPUT100), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT42), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n643), .B1(new_n644), .B2(G8gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(KEYINPUT16), .B(G8gat), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n637), .A2(KEYINPUT42), .A3(new_n641), .A4(new_n647), .ZN(new_n648));
  OAI211_X1 g447(.A(new_n645), .B(new_n648), .C1(KEYINPUT42), .C2(new_n647), .ZN(G1325gat));
  NAND2_X1  g448(.A1(new_n383), .A2(new_n372), .ZN(new_n650));
  AOI21_X1  g449(.A(G15gat), .B1(new_n637), .B2(new_n650), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n637), .A2(G15gat), .ZN(new_n652));
  INV_X1    g451(.A(new_n490), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n651), .B1(new_n652), .B2(new_n653), .ZN(G1326gat));
  NAND2_X1  g453(.A1(new_n637), .A2(new_n275), .ZN(new_n655));
  XNOR2_X1  g454(.A(KEYINPUT43), .B(G22gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(G1327gat));
  OR2_X1    g456(.A1(new_n577), .A2(new_n580), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n635), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n491), .A2(new_n549), .A3(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(G29gat), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n661), .A2(new_n662), .A3(new_n638), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(KEYINPUT101), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT45), .ZN(new_n665));
  OAI21_X1  g464(.A(KEYINPUT102), .B1(new_n545), .B2(new_n548), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n547), .A2(new_n543), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n539), .A2(new_n540), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT102), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n669), .A2(new_n670), .A3(new_n544), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n666), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n491), .A2(KEYINPUT44), .A3(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n483), .A2(new_n490), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n459), .A2(new_n385), .A3(new_n650), .A4(new_n453), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n458), .B1(new_n677), .B2(new_n641), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n549), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n675), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n674), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n660), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(new_n638), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT103), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n665), .B1(new_n686), .B2(new_n662), .ZN(G1328gat));
  INV_X1    g486(.A(G36gat), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n661), .A2(new_n688), .A3(new_n641), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT46), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n688), .B1(new_n684), .B2(new_n641), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT104), .ZN(G1329gat));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n682), .A2(new_n653), .A3(new_n683), .ZN(new_n695));
  INV_X1    g494(.A(new_n516), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n549), .B1(new_n676), .B2(new_n678), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n650), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n699), .A2(new_n696), .A3(new_n700), .ZN(new_n701));
  OAI211_X1 g500(.A(KEYINPUT105), .B(new_n694), .C1(new_n697), .C2(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n701), .B1(new_n695), .B2(new_n696), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT105), .ZN(new_n704));
  OAI21_X1  g503(.A(KEYINPUT106), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT47), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n702), .A2(KEYINPUT47), .A3(new_n705), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(G1330gat));
  NAND3_X1  g509(.A1(new_n684), .A2(G50gat), .A3(new_n275), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n512), .B1(new_n699), .B2(new_n459), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g513(.A(new_n634), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n491), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n581), .A2(new_n604), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n638), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g520(.A1(new_n718), .A2(new_n411), .ZN(new_n722));
  NOR2_X1   g521(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n723));
  AND2_X1   g522(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n722), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n725), .B1(new_n722), .B2(new_n723), .ZN(G1333gat));
  NAND3_X1  g525(.A1(new_n719), .A2(G71gat), .A3(new_n653), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n718), .A2(new_n700), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n727), .B1(G71gat), .B2(new_n728), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g529(.A1(new_n719), .A2(new_n275), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g531(.A1(new_n658), .A2(new_n604), .ZN(new_n733));
  OAI211_X1 g532(.A(new_n634), .B(new_n733), .C1(new_n674), .C2(new_n681), .ZN(new_n734));
  XOR2_X1   g533(.A(new_n734), .B(KEYINPUT107), .Z(new_n735));
  AND2_X1   g534(.A1(new_n735), .A2(G85gat), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT51), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n733), .B1(new_n698), .B2(KEYINPUT108), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT108), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n491), .A2(new_n739), .A3(new_n549), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n737), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n739), .B1(new_n491), .B2(new_n549), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n698), .A2(KEYINPUT108), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n742), .A2(new_n743), .A3(KEYINPUT51), .A4(new_n733), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n741), .A2(KEYINPUT109), .A3(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT109), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n746), .B(new_n737), .C1(new_n738), .C2(new_n740), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n745), .A2(new_n638), .A3(new_n634), .A4(new_n747), .ZN(new_n748));
  AOI22_X1  g547(.A1(new_n736), .A2(new_n638), .B1(new_n503), .B2(new_n748), .ZN(G1336gat));
  AOI21_X1  g548(.A(new_n504), .B1(new_n735), .B2(new_n641), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n741), .A2(new_n744), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n634), .A2(new_n504), .A3(new_n641), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT110), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(KEYINPUT52), .B1(new_n750), .B2(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n745), .A2(new_n747), .A3(new_n753), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(KEYINPUT111), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT111), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n745), .A2(new_n758), .A3(new_n747), .A4(new_n753), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(G92gat), .B1(new_n734), .B2(new_n411), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT52), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT112), .B1(new_n760), .B2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT112), .ZN(new_n766));
  AOI211_X1 g565(.A(new_n766), .B(new_n763), .C1(new_n757), .C2(new_n759), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n755), .B1(new_n765), .B2(new_n767), .ZN(G1337gat));
  AND3_X1   g567(.A1(new_n735), .A2(G99gat), .A3(new_n653), .ZN(new_n769));
  INV_X1    g568(.A(G99gat), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n745), .A2(new_n650), .A3(new_n634), .A4(new_n747), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(G1338gat));
  XNOR2_X1  g571(.A(KEYINPUT113), .B(G106gat), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n774), .B1(new_n735), .B2(new_n275), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n459), .A2(G106gat), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n751), .A2(new_n634), .A3(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(KEYINPUT53), .B1(new_n775), .B2(new_n777), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n745), .A2(new_n634), .A3(new_n747), .A4(new_n776), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT53), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n773), .B1(new_n734), .B2(new_n459), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n778), .A2(new_n782), .ZN(G1339gat));
  NAND4_X1  g582(.A1(new_n658), .A2(new_n549), .A3(new_n605), .A4(new_n715), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n585), .B1(new_n583), .B2(new_n584), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n589), .A2(new_n590), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n599), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT114), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OAI211_X1 g588(.A(KEYINPUT114), .B(new_n599), .C1(new_n785), .C2(new_n786), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n603), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n634), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n614), .A2(new_n608), .A3(new_n616), .ZN(new_n794));
  AND3_X1   g593(.A1(new_n794), .A2(new_n628), .A3(KEYINPUT54), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n623), .B1(new_n628), .B2(KEYINPUT54), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n793), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT54), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n625), .B1(new_n617), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n794), .A2(new_n628), .A3(KEYINPUT54), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n799), .A2(KEYINPUT55), .A3(new_n800), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n604), .A2(new_n797), .A3(new_n632), .A4(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n672), .B1(new_n792), .B2(new_n802), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n791), .A2(new_n632), .A3(new_n797), .A4(new_n801), .ZN(new_n804));
  OAI21_X1  g603(.A(KEYINPUT115), .B1(new_n673), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n797), .A2(new_n632), .A3(new_n801), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n603), .A2(new_n789), .A3(new_n790), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT115), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n808), .A2(new_n809), .A3(new_n672), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n803), .B1(new_n805), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n784), .B1(new_n811), .B2(new_n658), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n812), .A2(new_n384), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n641), .A2(new_n456), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT116), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n813), .A2(KEYINPUT116), .A3(new_n814), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(G113gat), .B1(new_n819), .B2(new_n605), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n581), .A2(new_n604), .A3(new_n634), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n810), .ZN(new_n822));
  INV_X1    g621(.A(new_n803), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n821), .B1(new_n824), .B2(new_n659), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n825), .A2(new_n455), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n814), .ZN(new_n827));
  OR2_X1    g626(.A1(new_n827), .A2(G113gat), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n820), .B1(new_n605), .B2(new_n828), .ZN(G1340gat));
  NOR3_X1   g628(.A1(new_n827), .A2(G120gat), .A3(new_n715), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n817), .A2(new_n634), .A3(new_n818), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n830), .B1(new_n831), .B2(G120gat), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n832), .B(KEYINPUT117), .ZN(G1341gat));
  NAND4_X1  g632(.A1(new_n817), .A2(G127gat), .A3(new_n658), .A4(new_n818), .ZN(new_n834));
  INV_X1    g633(.A(G127gat), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n835), .B1(new_n827), .B2(new_n659), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n834), .A2(new_n836), .ZN(G1342gat));
  NOR3_X1   g636(.A1(new_n827), .A2(G134gat), .A3(new_n549), .ZN(new_n838));
  XNOR2_X1  g637(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n838), .B(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(G134gat), .B1(new_n819), .B2(new_n549), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(G1343gat));
  NOR2_X1   g641(.A1(new_n423), .A2(new_n424), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n490), .A2(new_n814), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n792), .A2(new_n802), .ZN(new_n846));
  AOI22_X1  g645(.A1(new_n805), .A2(new_n810), .B1(new_n549), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n784), .B1(new_n847), .B2(new_n658), .ZN(new_n848));
  AND3_X1   g647(.A1(new_n848), .A2(KEYINPUT57), .A3(new_n275), .ZN(new_n849));
  XOR2_X1   g648(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n850));
  AOI21_X1  g649(.A(new_n850), .B1(new_n812), .B2(new_n275), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n845), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n843), .B1(new_n852), .B2(new_n605), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n825), .A2(new_n459), .A3(new_n844), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT121), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n855), .B1(new_n605), .B2(G141gat), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n604), .A2(KEYINPUT121), .A3(new_n416), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n854), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  XOR2_X1   g657(.A(KEYINPUT122), .B(KEYINPUT58), .Z(new_n859));
  NAND3_X1  g658(.A1(new_n853), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n858), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT120), .ZN(new_n862));
  INV_X1    g661(.A(new_n850), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n863), .B1(new_n825), .B2(new_n459), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n848), .A2(KEYINPUT57), .A3(new_n275), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n862), .B1(new_n866), .B2(new_n845), .ZN(new_n867));
  AOI211_X1 g666(.A(KEYINPUT120), .B(new_n844), .C1(new_n864), .C2(new_n865), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n604), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n861), .B1(new_n869), .B2(new_n843), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT58), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n860), .B1(new_n870), .B2(new_n871), .ZN(G1344gat));
  NAND3_X1  g671(.A1(new_n854), .A2(new_n229), .A3(new_n634), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(KEYINPUT123), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n852), .A2(KEYINPUT120), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n866), .A2(new_n862), .A3(new_n845), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n715), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n877), .A2(KEYINPUT59), .A3(new_n229), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT59), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n797), .A2(new_n801), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n880), .A2(KEYINPUT124), .A3(new_n680), .A4(new_n632), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT124), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n882), .B1(new_n806), .B2(new_n549), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n881), .A2(new_n791), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n846), .A2(new_n549), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n658), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n275), .B1(new_n886), .B2(new_n821), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT57), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n812), .A2(new_n275), .A3(new_n850), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n715), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(new_n845), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n879), .B1(new_n892), .B2(G148gat), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n874), .B1(new_n878), .B2(new_n893), .ZN(G1345gat));
  AOI21_X1  g693(.A(G155gat), .B1(new_n854), .B2(new_n658), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n659), .B1(new_n875), .B2(new_n876), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n895), .B1(new_n896), .B2(G155gat), .ZN(G1346gat));
  AOI21_X1  g696(.A(G162gat), .B1(new_n854), .B2(new_n680), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n673), .B1(new_n875), .B2(new_n876), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n898), .B1(new_n899), .B2(G162gat), .ZN(G1347gat));
  NOR2_X1   g699(.A1(new_n411), .A2(new_n638), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n826), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n902), .A2(new_n315), .A3(new_n604), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n813), .A2(new_n901), .ZN(new_n904));
  OAI21_X1  g703(.A(G169gat), .B1(new_n904), .B2(new_n605), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n903), .A2(new_n905), .ZN(G1348gat));
  AOI21_X1  g705(.A(G176gat), .B1(new_n902), .B2(new_n634), .ZN(new_n907));
  INV_X1    g706(.A(new_n904), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n715), .A2(new_n326), .A3(new_n327), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(G1349gat));
  AND2_X1   g709(.A1(new_n340), .A2(new_n345), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n902), .A2(new_n658), .A3(new_n912), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n337), .B(new_n338), .C1(new_n904), .C2(new_n659), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g715(.A(G190gat), .B1(new_n904), .B2(new_n549), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT61), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n902), .A2(new_n285), .A3(new_n672), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(G1351gat));
  NAND2_X1  g719(.A1(new_n490), .A2(new_n901), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n921), .B1(new_n889), .B2(new_n890), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(G197gat), .B1(new_n923), .B2(new_n605), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n490), .A2(new_n641), .A3(new_n275), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT125), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n925), .A2(new_n926), .ZN(new_n928));
  NOR4_X1   g727(.A1(new_n825), .A2(new_n638), .A3(new_n927), .A4(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(G197gat), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n929), .A2(new_n930), .A3(new_n604), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n924), .A2(new_n931), .ZN(G1352gat));
  INV_X1    g731(.A(G204gat), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n929), .A2(new_n933), .A3(new_n634), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT62), .ZN(new_n935));
  INV_X1    g734(.A(new_n921), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n933), .B1(new_n891), .B2(new_n936), .ZN(new_n937));
  OR2_X1    g736(.A1(new_n935), .A2(new_n937), .ZN(G1353gat));
  NAND3_X1  g737(.A1(new_n929), .A2(new_n206), .A3(new_n658), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT126), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n922), .A2(new_n940), .A3(new_n658), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n940), .B1(new_n922), .B2(new_n658), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g742(.A(KEYINPUT63), .B1(new_n943), .B2(G211gat), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT63), .ZN(new_n945));
  NOR4_X1   g744(.A1(new_n941), .A2(new_n942), .A3(new_n945), .A4(new_n206), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n939), .B1(new_n944), .B2(new_n946), .ZN(G1354gat));
  AOI21_X1  g746(.A(G218gat), .B1(new_n929), .B2(new_n672), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT127), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n549), .B1(new_n923), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n209), .B1(new_n922), .B2(KEYINPUT127), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(G1355gat));
endmodule


