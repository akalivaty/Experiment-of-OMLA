//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 1 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 0 0 1 1 0 1 1 1 0 1 0 1 1 1 1 1 1 1 0 0 1 1 1 1 1 1 0 1 1 1 1 0 0 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:19 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n564, new_n565, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n583, new_n584, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n621, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1194, new_n1195;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  INV_X1    g032(.A(new_n452), .ZN(new_n458));
  AOI21_X1  g033(.A(new_n457), .B1(new_n458), .B2(G2106), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT65), .B(G2105), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n464), .A2(new_n465), .A3(G137), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n467), .A2(G101), .A3(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n466), .A2(KEYINPUT68), .A3(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g045(.A(KEYINPUT68), .B1(new_n466), .B2(new_n468), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n467), .A2(KEYINPUT65), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT65), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G125), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n477), .B1(new_n462), .B2(new_n463), .ZN(new_n478));
  NAND2_X1  g053(.A1(G113), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(KEYINPUT66), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT66), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n481), .A2(G113), .A3(G2104), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n476), .B1(new_n478), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(KEYINPUT67), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT67), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(new_n476), .C1(new_n478), .C2(new_n483), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n472), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G160));
  AND2_X1   g065(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n491));
  NOR2_X1   g066(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G136), .ZN(new_n495));
  XOR2_X1   g070(.A(new_n495), .B(KEYINPUT69), .Z(new_n496));
  OAI221_X1 g071(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n465), .C2(G112), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n493), .A2(new_n465), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G124), .ZN(new_n499));
  AND3_X1   g074(.A1(new_n496), .A2(new_n497), .A3(new_n499), .ZN(G162));
  NAND3_X1  g075(.A1(new_n473), .A2(new_n475), .A3(G138), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT4), .B1(new_n501), .B2(new_n493), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n464), .A2(new_n465), .A3(new_n503), .A4(G138), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g080(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n506));
  INV_X1    g081(.A(G114), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n506), .B1(new_n507), .B2(G2105), .ZN(new_n508));
  AND2_X1   g083(.A1(G126), .A2(G2105), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n509), .B1(new_n491), .B2(new_n492), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT70), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OAI211_X1 g087(.A(KEYINPUT70), .B(new_n509), .C1(new_n491), .C2(new_n492), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n508), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n505), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(G164));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G62), .ZN(new_n523));
  NAND2_X1  g098(.A1(G75), .A2(G543), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n517), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n525), .A2(KEYINPUT71), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(KEYINPUT71), .ZN(new_n527));
  OR2_X1    g102(.A1(KEYINPUT6), .A2(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(KEYINPUT6), .A2(G651), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n528), .A2(new_n529), .B1(new_n520), .B2(new_n521), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n519), .B1(new_n528), .B2(new_n529), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n530), .A2(G88), .B1(new_n531), .B2(G50), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n526), .A2(new_n527), .A3(new_n532), .ZN(G303));
  INV_X1    g108(.A(G303), .ZN(G166));
  NAND2_X1  g109(.A1(new_n528), .A2(new_n529), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G89), .ZN(new_n536));
  NAND2_X1  g111(.A1(G63), .A2(G651), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(new_n522), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n531), .A2(G51), .ZN(new_n540));
  NAND3_X1  g115(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT7), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n539), .A2(new_n540), .A3(new_n542), .ZN(G286));
  INV_X1    g118(.A(G286), .ZN(G168));
  AOI22_X1  g119(.A1(new_n530), .A2(G90), .B1(new_n531), .B2(G52), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  AND2_X1   g121(.A1(new_n520), .A2(new_n521), .ZN(new_n547));
  INV_X1    g122(.A(G64), .ZN(new_n548));
  INV_X1    g123(.A(G77), .ZN(new_n549));
  OAI22_X1  g124(.A1(new_n547), .A2(new_n548), .B1(new_n549), .B2(new_n519), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT72), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n517), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OAI221_X1 g127(.A(KEYINPUT72), .B1(new_n549), .B2(new_n519), .C1(new_n547), .C2(new_n548), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n546), .B1(new_n552), .B2(new_n553), .ZN(G171));
  NAND2_X1  g129(.A1(new_n531), .A2(G43), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n535), .A2(new_n522), .ZN(new_n556));
  INV_X1    g131(.A(G81), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n522), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n559), .A2(new_n517), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(G153));
  NAND4_X1  g137(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND4_X1  g140(.A1(G319), .A2(G483), .A3(G661), .A4(new_n565), .ZN(G188));
  INV_X1    g141(.A(KEYINPUT73), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(G65), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n547), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G651), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n530), .A2(G91), .ZN(new_n572));
  AND2_X1   g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n535), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G53), .ZN(new_n575));
  OAI21_X1  g150(.A(KEYINPUT9), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT9), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n531), .A2(new_n577), .A3(G53), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n567), .B1(new_n573), .B2(new_n579), .ZN(new_n580));
  AND4_X1   g155(.A1(new_n567), .A2(new_n579), .A3(new_n571), .A4(new_n572), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n580), .A2(new_n581), .ZN(G299));
  NAND2_X1  g157(.A1(new_n550), .A2(new_n551), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n583), .A2(G651), .A3(new_n553), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(new_n545), .ZN(G301));
  NAND2_X1  g160(.A1(new_n530), .A2(G87), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n522), .B2(G74), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n531), .A2(G49), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(G288));
  AOI22_X1  g164(.A1(new_n530), .A2(G86), .B1(new_n531), .B2(G48), .ZN(new_n590));
  INV_X1    g165(.A(G61), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n591), .B1(new_n520), .B2(new_n521), .ZN(new_n592));
  AND2_X1   g167(.A1(G73), .A2(G543), .ZN(new_n593));
  OAI211_X1 g168(.A(KEYINPUT74), .B(G651), .C1(new_n592), .C2(new_n593), .ZN(new_n594));
  AND2_X1   g169(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT74), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n592), .A2(new_n593), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n597), .B2(new_n517), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n595), .A2(new_n598), .ZN(G305));
  AOI22_X1  g174(.A1(new_n522), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n600), .A2(new_n517), .ZN(new_n601));
  OR2_X1    g176(.A1(new_n601), .A2(KEYINPUT75), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(KEYINPUT75), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n530), .A2(G85), .B1(new_n531), .B2(G47), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  AND3_X1   g181(.A1(new_n535), .A2(new_n522), .A3(G92), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT10), .ZN(new_n608));
  OR2_X1    g183(.A1(new_n574), .A2(KEYINPUT76), .ZN(new_n609));
  INV_X1    g184(.A(G54), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n610), .B1(new_n574), .B2(KEYINPUT76), .ZN(new_n611));
  NAND2_X1  g186(.A1(G79), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(G66), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n547), .B2(new_n613), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n609), .A2(new_n611), .B1(G651), .B2(new_n614), .ZN(new_n615));
  AND2_X1   g190(.A1(new_n608), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n606), .B1(new_n616), .B2(G868), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT77), .Z(G284));
  XOR2_X1   g193(.A(new_n617), .B(KEYINPUT78), .Z(G321));
  NAND2_X1  g194(.A1(G286), .A2(G868), .ZN(new_n620));
  INV_X1    g195(.A(G299), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(G868), .ZN(G297));
  OAI21_X1  g197(.A(new_n620), .B1(new_n621), .B2(G868), .ZN(G280));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n616), .B1(new_n624), .B2(G860), .ZN(G148));
  OR2_X1    g200(.A1(new_n558), .A2(new_n560), .ZN(new_n626));
  INV_X1    g201(.A(G868), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n608), .A2(new_n615), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n629), .A2(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n628), .B1(new_n630), .B2(new_n627), .ZN(G323));
  XNOR2_X1  g206(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g207(.A(KEYINPUT79), .B(KEYINPUT12), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n467), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT13), .B(G2100), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  AOI22_X1  g212(.A1(G123), .A2(new_n498), .B1(new_n494), .B2(G135), .ZN(new_n638));
  OAI221_X1 g213(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n465), .C2(G111), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n640), .A2(KEYINPUT80), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(KEYINPUT80), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  AND2_X1   g219(.A1(new_n644), .A2(G2096), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n644), .A2(G2096), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n637), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT81), .Z(G156));
  XOR2_X1   g223(.A(KEYINPUT82), .B(KEYINPUT14), .Z(new_n649));
  XOR2_X1   g224(.A(KEYINPUT15), .B(G2435), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2438), .ZN(new_n651));
  XOR2_X1   g226(.A(G2427), .B(G2430), .Z(new_n652));
  AOI21_X1  g227(.A(new_n649), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n653), .B1(new_n651), .B2(new_n652), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2451), .B(G2454), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT16), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1341), .B(G1348), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n654), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2443), .B(G2446), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n661), .A2(G14), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n659), .A2(new_n660), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(G401));
  XOR2_X1   g239(.A(G2067), .B(G2678), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT83), .ZN(new_n666));
  NOR2_X1   g241(.A1(G2072), .A2(G2078), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n442), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2084), .B(G2090), .ZN(new_n669));
  NOR3_X1   g244(.A1(new_n666), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT18), .ZN(new_n671));
  INV_X1    g246(.A(new_n668), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n672), .A2(KEYINPUT84), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n672), .A2(KEYINPUT84), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n666), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n668), .B(KEYINPUT17), .ZN(new_n676));
  OAI211_X1 g251(.A(new_n675), .B(new_n669), .C1(new_n666), .C2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n669), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n666), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n671), .A2(new_n677), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(G2100), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT85), .B(G2096), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(G227));
  XNOR2_X1  g258(.A(G1956), .B(G2474), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1961), .B(G1966), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G1971), .B(G1976), .Z(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT86), .B(KEYINPUT19), .ZN(new_n688));
  AND2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n687), .A2(new_n688), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n684), .A2(new_n685), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n686), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n691), .A2(KEYINPUT87), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NOR3_X1   g270(.A1(new_n689), .A2(new_n692), .A3(new_n690), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT20), .Z(new_n697));
  NAND2_X1  g272(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1991), .B(G1996), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1981), .B(G1986), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(G229));
  NOR2_X1   g279(.A1(G29), .A2(G35), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(G162), .B2(G29), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT29), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(G2090), .Z(new_n708));
  NOR2_X1   g283(.A1(G29), .A2(G33), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT95), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT25), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(G139), .B2(new_n494), .ZN(new_n713));
  AOI22_X1  g288(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n714), .A2(new_n465), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT96), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n715), .A2(new_n716), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n713), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT97), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g296(.A1(new_n713), .A2(KEYINPUT97), .A3(new_n717), .A4(new_n718), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(G29), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n710), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G2072), .ZN(new_n726));
  INV_X1    g301(.A(G16), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G20), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT23), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(new_n621), .B2(new_n727), .ZN(new_n730));
  INV_X1    g305(.A(G1956), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n708), .A2(new_n726), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n724), .A2(G32), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n498), .A2(G129), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT98), .ZN(new_n736));
  AND3_X1   g311(.A1(new_n467), .A2(G105), .A3(G2104), .ZN(new_n737));
  NAND3_X1  g312(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT26), .ZN(new_n739));
  AOI211_X1 g314(.A(new_n737), .B(new_n739), .C1(G141), .C2(new_n494), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n736), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n734), .B1(new_n741), .B2(new_n724), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT27), .Z(new_n743));
  OR2_X1    g318(.A1(new_n743), .A2(G1996), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(G1996), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n643), .A2(new_n724), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n746), .A2(KEYINPUT99), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n724), .A2(G26), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT28), .Z(new_n749));
  AOI22_X1  g324(.A1(G128), .A2(new_n498), .B1(new_n494), .B2(G140), .ZN(new_n750));
  OAI221_X1 g325(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n465), .C2(G116), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n749), .B1(new_n752), .B2(G29), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT94), .B(G2067), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n747), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(G164), .A2(new_n724), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G27), .B2(new_n724), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n746), .A2(KEYINPUT99), .B1(G2078), .B2(new_n759), .ZN(new_n760));
  NAND4_X1  g335(.A1(new_n744), .A2(new_n745), .A3(new_n756), .A4(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(G16), .A2(G19), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n561), .B2(G16), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT93), .B(G1341), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(KEYINPUT31), .A2(G11), .ZN(new_n766));
  AND2_X1   g341(.A1(KEYINPUT31), .A2(G11), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT30), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n768), .A2(G28), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n724), .B1(new_n768), .B2(G28), .ZN(new_n770));
  OAI221_X1 g345(.A(new_n765), .B1(new_n766), .B2(new_n767), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n727), .A2(G21), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G168), .B2(new_n727), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n773), .A2(G1966), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(G1966), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n774), .B(new_n775), .C1(new_n763), .C2(new_n764), .ZN(new_n776));
  INV_X1    g351(.A(G2078), .ZN(new_n777));
  AOI211_X1 g352(.A(new_n771), .B(new_n776), .C1(new_n777), .C2(new_n758), .ZN(new_n778));
  NAND2_X1  g353(.A1(G301), .A2(G16), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n727), .A2(G5), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT24), .ZN(new_n783));
  INV_X1    g358(.A(G34), .ZN(new_n784));
  AOI21_X1  g359(.A(G29), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(new_n783), .B2(new_n784), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G160), .B2(new_n724), .ZN(new_n787));
  INV_X1    g362(.A(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(G2084), .ZN(new_n789));
  AOI22_X1  g364(.A1(new_n782), .A2(G1961), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(G1961), .ZN(new_n791));
  AOI22_X1  g366(.A1(new_n781), .A2(new_n791), .B1(new_n787), .B2(G2084), .ZN(new_n792));
  NOR2_X1   g367(.A1(G4), .A2(G16), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT91), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n629), .B2(new_n727), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT92), .B(G1348), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n778), .A2(new_n790), .A3(new_n792), .A4(new_n797), .ZN(new_n798));
  NOR3_X1   g373(.A1(new_n733), .A2(new_n761), .A3(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n727), .A2(G6), .ZN(new_n801));
  INV_X1    g376(.A(G305), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n801), .B1(new_n802), .B2(new_n727), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT89), .Z(new_n804));
  XOR2_X1   g379(.A(KEYINPUT32), .B(G1981), .Z(new_n805));
  OR2_X1    g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n804), .A2(new_n805), .ZN(new_n807));
  NAND2_X1  g382(.A1(G166), .A2(G16), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G16), .B2(G22), .ZN(new_n809));
  INV_X1    g384(.A(G1971), .ZN(new_n810));
  AND2_X1   g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n809), .A2(new_n810), .ZN(new_n812));
  NOR2_X1   g387(.A1(G16), .A2(G23), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT90), .Z(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(G288), .B2(new_n727), .ZN(new_n815));
  XNOR2_X1  g390(.A(KEYINPUT33), .B(G1976), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NOR3_X1   g392(.A1(new_n811), .A2(new_n812), .A3(new_n817), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n806), .A2(new_n807), .A3(new_n818), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n819), .A2(KEYINPUT34), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(KEYINPUT34), .ZN(new_n821));
  MUX2_X1   g396(.A(G24), .B(G290), .S(G16), .Z(new_n822));
  AND2_X1   g397(.A1(new_n822), .A2(G1986), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n822), .A2(G1986), .ZN(new_n824));
  NOR2_X1   g399(.A1(G25), .A2(G29), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n498), .A2(G119), .ZN(new_n826));
  OAI221_X1 g401(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n465), .C2(G107), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n494), .A2(G131), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n825), .B1(new_n830), .B2(G29), .ZN(new_n831));
  XOR2_X1   g406(.A(KEYINPUT35), .B(G1991), .Z(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT88), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n831), .B(new_n833), .ZN(new_n834));
  NOR3_X1   g409(.A1(new_n823), .A2(new_n824), .A3(new_n834), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n820), .A2(new_n821), .A3(new_n835), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n836), .A2(KEYINPUT36), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(KEYINPUT36), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n800), .B1(new_n837), .B2(new_n838), .ZN(G311));
  NAND2_X1  g414(.A1(new_n837), .A2(new_n838), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(new_n799), .ZN(G150));
  AOI22_X1  g416(.A1(new_n530), .A2(G93), .B1(new_n531), .B2(G55), .ZN(new_n842));
  AOI22_X1  g417(.A1(new_n522), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n842), .B1(new_n517), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(G860), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(KEYINPUT37), .Z(new_n846));
  NAND3_X1  g421(.A1(new_n626), .A2(KEYINPUT100), .A3(new_n844), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n531), .A2(G55), .ZN(new_n848));
  INV_X1    g423(.A(G93), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n848), .B1(new_n556), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n843), .A2(new_n517), .ZN(new_n851));
  OAI21_X1  g426(.A(KEYINPUT100), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT100), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n842), .B(new_n853), .C1(new_n517), .C2(new_n843), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n852), .A2(new_n561), .A3(new_n854), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n847), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT38), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n629), .A2(new_n624), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n857), .B(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(KEYINPUT39), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(KEYINPUT101), .Z(new_n862));
  INV_X1    g437(.A(G860), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n863), .B1(new_n860), .B2(KEYINPUT39), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n846), .B1(new_n862), .B2(new_n864), .ZN(G145));
  NAND3_X1  g440(.A1(new_n641), .A2(KEYINPUT102), .A3(new_n642), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(KEYINPUT102), .B1(new_n641), .B2(new_n642), .ZN(new_n868));
  OAI21_X1  g443(.A(G160), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n868), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n870), .A2(new_n489), .A3(new_n866), .ZN(new_n871));
  AND3_X1   g446(.A1(new_n869), .A2(new_n871), .A3(G162), .ZN(new_n872));
  AOI21_X1  g447(.A(G162), .B1(new_n869), .B2(new_n871), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(KEYINPUT104), .B(KEYINPUT105), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  AOI22_X1  g451(.A1(G130), .A2(new_n498), .B1(new_n494), .B2(G142), .ZN(new_n877));
  OAI221_X1 g452(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n465), .C2(G118), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(new_n635), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(new_n829), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n880), .A2(new_n829), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n876), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n883), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n885), .A2(new_n881), .A3(new_n875), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT103), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n723), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n721), .A2(KEYINPUT103), .A3(new_n722), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n736), .A2(new_n740), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(new_n752), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n736), .A2(new_n740), .A3(new_n751), .A4(new_n750), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n892), .A2(new_n515), .A3(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n515), .B1(new_n892), .B2(new_n893), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n889), .B(new_n890), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n721), .A2(new_n722), .ZN(new_n898));
  INV_X1    g473(.A(new_n896), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n898), .A2(new_n899), .A3(KEYINPUT103), .A4(new_n894), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n887), .B1(new_n897), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n874), .B1(new_n901), .B2(KEYINPUT106), .ZN(new_n902));
  INV_X1    g477(.A(new_n889), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n890), .B1(new_n895), .B2(new_n896), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n900), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n887), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT106), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n897), .A2(new_n887), .A3(new_n900), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(G37), .B1(new_n902), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n907), .A2(new_n909), .A3(new_n874), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n912), .A2(KEYINPUT107), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n912), .A2(KEYINPUT107), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n911), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n915), .B(new_n916), .ZN(G395));
  NAND2_X1  g492(.A1(new_n844), .A2(new_n627), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n629), .B1(new_n580), .B2(new_n581), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n573), .A2(new_n567), .A3(new_n579), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n576), .A2(new_n578), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n571), .A2(new_n572), .ZN(new_n922));
  OAI21_X1  g497(.A(KEYINPUT73), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n616), .A2(new_n920), .A3(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n919), .A2(KEYINPUT109), .A3(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT109), .ZN(new_n926));
  NAND3_X1  g501(.A1(G299), .A2(new_n926), .A3(new_n616), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n847), .A2(new_n855), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n929), .B(new_n630), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  XOR2_X1   g506(.A(new_n931), .B(KEYINPUT110), .Z(new_n932));
  NAND3_X1  g507(.A1(new_n925), .A2(KEYINPUT41), .A3(new_n927), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT41), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n919), .A2(new_n934), .A3(new_n924), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n933), .A2(new_n930), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n932), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n802), .B(G303), .ZN(new_n938));
  INV_X1    g513(.A(G288), .ZN(new_n939));
  XNOR2_X1  g514(.A(G290), .B(new_n939), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n938), .B(new_n940), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n941), .B(KEYINPUT42), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n937), .B(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n918), .B1(new_n943), .B2(new_n627), .ZN(G295));
  OAI21_X1  g519(.A(new_n918), .B1(new_n943), .B2(new_n627), .ZN(G331));
  XOR2_X1   g520(.A(KEYINPUT111), .B(KEYINPUT43), .Z(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT112), .ZN(new_n948));
  NAND3_X1  g523(.A1(G301), .A2(new_n948), .A3(G168), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT112), .B1(G171), .B2(G286), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n584), .A2(G286), .A3(new_n545), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT113), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(G171), .A2(KEYINPUT113), .A3(G286), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n951), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(new_n929), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n951), .A2(new_n956), .A3(new_n856), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n933), .A2(new_n958), .A3(new_n935), .A4(new_n959), .ZN(new_n960));
  AND3_X1   g535(.A1(new_n951), .A2(new_n956), .A3(new_n856), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n856), .B1(new_n951), .B2(new_n956), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n927), .B(new_n925), .C1(new_n961), .C2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n960), .A2(new_n963), .A3(new_n941), .ZN(new_n964));
  INV_X1    g539(.A(G37), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n941), .B1(new_n960), .B2(new_n963), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n947), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(KEYINPUT114), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT114), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n970), .B(new_n947), .C1(new_n966), .C2(new_n967), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT44), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n964), .A2(new_n965), .ZN(new_n974));
  INV_X1    g549(.A(new_n941), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n928), .A2(new_n934), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n961), .A2(new_n962), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT115), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n919), .A2(new_n924), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT41), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n976), .A2(new_n977), .A3(new_n978), .A4(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n963), .A2(KEYINPUT115), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n958), .A2(new_n980), .A3(new_n959), .ZN(new_n983));
  AOI21_X1  g558(.A(KEYINPUT41), .B1(new_n925), .B2(new_n927), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n975), .B(new_n981), .C1(new_n982), .C2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n974), .A2(new_n986), .A3(new_n946), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT116), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n974), .A2(new_n986), .A3(KEYINPUT116), .A4(new_n946), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n972), .A2(new_n973), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT43), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n992), .B1(new_n974), .B2(new_n986), .ZN(new_n993));
  NOR3_X1   g568(.A1(new_n966), .A2(new_n967), .A3(new_n947), .ZN(new_n994));
  OAI21_X1  g569(.A(KEYINPUT44), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n991), .A2(new_n995), .ZN(G397));
  INV_X1    g571(.A(new_n471), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n488), .A2(G40), .A3(new_n997), .A4(new_n469), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT117), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n472), .A2(KEYINPUT117), .A3(G40), .A4(new_n488), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(G1384), .B1(new_n505), .B2(new_n514), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1003), .A2(KEYINPUT45), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(G1996), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n741), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(G2067), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n752), .B(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n891), .A2(G1996), .ZN(new_n1011));
  AND3_X1   g586(.A1(new_n1008), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n830), .A2(new_n832), .ZN(new_n1013));
  OR2_X1    g588(.A1(new_n830), .A2(new_n832), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(G290), .B(G1986), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1006), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT126), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT118), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1019), .B1(new_n1003), .B2(KEYINPUT45), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT45), .ZN(new_n1021));
  AOI211_X1 g596(.A(new_n1021), .B(G1384), .C1(new_n505), .C2(new_n514), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G1384), .ZN(new_n1024));
  AND2_X1   g599(.A1(new_n502), .A2(new_n504), .ZN(new_n1025));
  INV_X1    g600(.A(new_n508), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT70), .B1(new_n464), .B2(new_n509), .ZN(new_n1027));
  INV_X1    g602(.A(new_n513), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1026), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1024), .B1(new_n1025), .B2(new_n1029), .ZN(new_n1030));
  NOR3_X1   g605(.A1(new_n1030), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1002), .B(new_n777), .C1(new_n1023), .C2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n1003), .B(KEYINPUT50), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1002), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(new_n791), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1030), .A2(new_n1021), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1003), .A2(KEYINPUT45), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1038), .A2(new_n1019), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(KEYINPUT53), .A2(G40), .ZN(new_n1043));
  OR2_X1    g618(.A1(new_n777), .A2(KEYINPUT125), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n777), .A2(KEYINPUT125), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1043), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1042), .A2(new_n472), .A3(new_n484), .A4(new_n1046), .ZN(new_n1047));
  AND3_X1   g622(.A1(new_n1034), .A2(new_n1037), .A3(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1018), .B1(new_n1048), .B2(G301), .ZN(new_n1049));
  AOI22_X1  g624(.A1(new_n1032), .A2(new_n1033), .B1(new_n791), .B2(new_n1036), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(new_n1047), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1051), .A2(KEYINPUT126), .A3(G171), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1004), .A2(new_n1022), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1002), .A2(new_n1053), .A3(KEYINPUT53), .A4(new_n777), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1034), .A2(G301), .A3(new_n1037), .A4(new_n1054), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n1055), .A2(KEYINPUT54), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1049), .A2(new_n1052), .A3(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1002), .A2(new_n789), .A3(new_n1035), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1059), .B1(new_n1001), .B2(new_n1000), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1058), .B(G168), .C1(new_n1060), .C2(G1966), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(G8), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1002), .A2(new_n1053), .ZN(new_n1063));
  INV_X1    g638(.A(G1966), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(G168), .B1(new_n1065), .B2(new_n1058), .ZN(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT51), .B1(new_n1062), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT51), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1061), .A2(new_n1068), .A3(G8), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT61), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1036), .A2(new_n731), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n573), .A2(new_n579), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT57), .B1(new_n579), .B2(KEYINPUT121), .ZN(new_n1073));
  XNOR2_X1  g648(.A(new_n1072), .B(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1071), .A2(new_n1074), .ZN(new_n1075));
  XNOR2_X1  g650(.A(KEYINPUT56), .B(G2072), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1042), .A2(new_n1002), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT122), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  AOI22_X1  g654(.A1(new_n1040), .A2(new_n1041), .B1(new_n1001), .B2(new_n1000), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1080), .A2(KEYINPUT122), .A3(new_n1076), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1075), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  AOI22_X1  g657(.A1(new_n1067), .A2(new_n1069), .B1(new_n1070), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT54), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n1050), .A2(G301), .A3(new_n1047), .ZN(new_n1085));
  AOI21_X1  g660(.A(G301), .B1(new_n1050), .B2(new_n1054), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1084), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(G8), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1088), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1089));
  INV_X1    g664(.A(G1976), .ZN(new_n1090));
  NOR2_X1   g665(.A1(G288), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  XNOR2_X1  g667(.A(KEYINPUT119), .B(G1976), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT52), .B1(G288), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1089), .A2(new_n1092), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(G1981), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n595), .A2(new_n1096), .A3(new_n598), .ZN(new_n1097));
  INV_X1    g672(.A(new_n598), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n590), .A2(new_n594), .ZN(new_n1099));
  OAI21_X1  g674(.A(G1981), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  AND3_X1   g675(.A1(new_n1097), .A2(new_n1100), .A3(KEYINPUT49), .ZN(new_n1101));
  AOI21_X1  g676(.A(KEYINPUT49), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1089), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1095), .A2(new_n1104), .ZN(new_n1105));
  AOI211_X1 g680(.A(new_n1088), .B(new_n1091), .C1(new_n1002), .C2(new_n1003), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT52), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1109));
  OAI22_X1  g684(.A1(new_n1080), .A2(G1971), .B1(new_n1036), .B2(G2090), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(G8), .ZN(new_n1111));
  NAND2_X1  g686(.A1(G303), .A2(G8), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n1112), .B(KEYINPUT55), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1113), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1110), .A2(G8), .A3(new_n1115), .ZN(new_n1116));
  AND3_X1   g691(.A1(new_n1109), .A2(new_n1114), .A3(new_n1116), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1057), .A2(new_n1083), .A3(new_n1087), .A4(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1119), .A2(new_n1071), .A3(new_n1074), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n1079), .A2(new_n1081), .B1(new_n731), .B2(new_n1036), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1121), .A2(new_n1074), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1002), .A2(new_n1009), .A3(new_n1003), .ZN(new_n1123));
  INV_X1    g698(.A(G1348), .ZN(new_n1124));
  AOI22_X1  g699(.A1(new_n1123), .A2(KEYINPUT123), .B1(new_n1036), .B2(new_n1124), .ZN(new_n1125));
  OR2_X1    g700(.A1(new_n1123), .A2(KEYINPUT123), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n629), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1120), .B1(new_n1122), .B2(new_n1127), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1125), .B(new_n1126), .C1(KEYINPUT60), .C2(new_n616), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n616), .A2(KEYINPUT60), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n1129), .B(new_n1130), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1120), .B(KEYINPUT61), .C1(new_n1074), .C2(new_n1121), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1133));
  XOR2_X1   g708(.A(KEYINPUT58), .B(G1341), .Z(new_n1134));
  AOI21_X1  g709(.A(G1996), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1135));
  AOI22_X1  g710(.A1(new_n1133), .A2(new_n1134), .B1(new_n1042), .B2(new_n1135), .ZN(new_n1136));
  OR3_X1    g711(.A1(new_n1136), .A2(KEYINPUT124), .A3(new_n626), .ZN(new_n1137));
  OAI21_X1  g712(.A(KEYINPUT124), .B1(new_n1136), .B2(new_n626), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1137), .A2(KEYINPUT59), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT59), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1131), .A2(new_n1132), .A3(new_n1139), .A4(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1118), .B1(new_n1128), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(KEYINPUT62), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT62), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1067), .A2(new_n1147), .A3(new_n1069), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1146), .A2(new_n1086), .A3(new_n1117), .A4(new_n1148), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n1095), .B(new_n1104), .C1(new_n1107), .C2(new_n1106), .ZN(new_n1150));
  NOR2_X1   g725(.A1(G288), .A2(G1976), .ZN(new_n1151));
  AOI22_X1  g726(.A1(new_n1104), .A2(new_n1151), .B1(new_n1096), .B2(new_n802), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1089), .ZN(new_n1153));
  OAI22_X1  g728(.A1(new_n1150), .A2(new_n1116), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1154), .B(KEYINPUT120), .ZN(new_n1155));
  AOI211_X1 g730(.A(new_n1088), .B(G286), .C1(new_n1065), .C2(new_n1058), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1109), .A2(new_n1114), .A3(new_n1116), .A4(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT63), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  AOI22_X1  g734(.A1(new_n1106), .A2(new_n1094), .B1(new_n1089), .B2(new_n1103), .ZN(new_n1160));
  OAI21_X1  g735(.A(KEYINPUT52), .B1(new_n1153), .B2(new_n1091), .ZN(new_n1161));
  AND3_X1   g736(.A1(new_n1116), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1162), .A2(KEYINPUT63), .A3(new_n1114), .A4(new_n1156), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1159), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1149), .A2(new_n1155), .A3(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1017), .B1(new_n1144), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1010), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1006), .B1(new_n891), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT46), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1169), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1170));
  NOR3_X1   g745(.A1(new_n1005), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1168), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n1172), .B(KEYINPUT47), .ZN(new_n1173));
  XOR2_X1   g748(.A(new_n1013), .B(KEYINPUT127), .Z(new_n1174));
  INV_X1    g749(.A(new_n1012), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1174), .B1(new_n1175), .B2(new_n1006), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n752), .A2(G2067), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1006), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  OR3_X1    g753(.A1(new_n1005), .A2(G1986), .A3(G290), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT48), .ZN(new_n1180));
  OR2_X1    g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1015), .A2(new_n1006), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  AND3_X1   g759(.A1(new_n1173), .A2(new_n1178), .A3(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1166), .A2(new_n1185), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g761(.A(G319), .B1(new_n662), .B2(new_n663), .ZN(new_n1188));
  OR2_X1    g762(.A1(G227), .A2(new_n1188), .ZN(new_n1189));
  NOR2_X1   g763(.A1(G229), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g764(.A1(new_n915), .A2(new_n1190), .ZN(new_n1191));
  AND2_X1   g765(.A1(new_n989), .A2(new_n990), .ZN(new_n1192));
  AOI21_X1  g766(.A(new_n1191), .B1(new_n972), .B2(new_n1192), .ZN(G308));
  NAND2_X1  g767(.A1(new_n1192), .A2(new_n972), .ZN(new_n1194));
  INV_X1    g768(.A(new_n1191), .ZN(new_n1195));
  NAND2_X1  g769(.A1(new_n1194), .A2(new_n1195), .ZN(G225));
endmodule


