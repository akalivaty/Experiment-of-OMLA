//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 1 1 0 1 1 0 1 0 1 0 1 0 1 0 0 0 0 0 0 0 0 1 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 0 1 1 0 1 1 0 0 0 1 1 1 1 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:30 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1276, new_n1277, new_n1279,
    new_n1280, new_n1281, new_n1282, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT64), .Z(new_n209));
  XNOR2_X1  g0009(.A(KEYINPUT65), .B(G244), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(G77), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G107), .A2(G264), .ZN(new_n217));
  NAND4_X1  g0017(.A1(new_n214), .A2(new_n215), .A3(new_n216), .A4(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n209), .B1(new_n213), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT66), .ZN(new_n220));
  INV_X1    g0020(.A(KEYINPUT1), .ZN(new_n221));
  AND2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n209), .A2(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT0), .Z(new_n225));
  NOR2_X1   g0025(.A1(new_n220), .A2(new_n221), .ZN(new_n226));
  INV_X1    g0026(.A(G58), .ZN(new_n227));
  INV_X1    g0027(.A(G68), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(G50), .ZN(new_n230));
  INV_X1    g0030(.A(G20), .ZN(new_n231));
  NAND2_X1  g0031(.A1(G1), .A2(G13), .ZN(new_n232));
  NOR3_X1   g0032(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  NOR4_X1   g0033(.A1(new_n222), .A2(new_n225), .A3(new_n226), .A4(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  INV_X1    g0035(.A(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT2), .B(G226), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G358));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT67), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G68), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n232), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G13), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n255), .A2(G1), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G20), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT71), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n254), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  NOR3_X1   g0059(.A1(new_n255), .A2(new_n231), .A3(G1), .ZN(new_n260));
  OAI21_X1  g0060(.A(KEYINPUT71), .B1(new_n260), .B2(new_n253), .ZN(new_n261));
  AND2_X1   g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G1), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G20), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n262), .A2(G68), .A3(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G20), .A2(G33), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n266), .A2(G50), .B1(G20), .B2(new_n228), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n231), .A2(G33), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n267), .B1(new_n212), .B2(new_n268), .ZN(new_n269));
  AND2_X1   g0069(.A1(new_n269), .A2(new_n253), .ZN(new_n270));
  OR2_X1    g0070(.A1(new_n270), .A2(KEYINPUT11), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n260), .A2(new_n228), .ZN(new_n272));
  XNOR2_X1  g0072(.A(new_n272), .B(KEYINPUT12), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n270), .A2(KEYINPUT11), .ZN(new_n274));
  AND4_X1   g0074(.A1(new_n265), .A2(new_n271), .A3(new_n273), .A4(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT14), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT13), .ZN(new_n277));
  INV_X1    g0077(.A(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT3), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT3), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G33), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n279), .A2(new_n281), .A3(G232), .A4(G1698), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT72), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT3), .B(G33), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n285), .A2(KEYINPUT72), .A3(G232), .A4(G1698), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G1698), .ZN(new_n288));
  NAND4_X1  g0088(.A1(new_n279), .A2(new_n281), .A3(G226), .A4(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(G33), .A2(G97), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n287), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(G33), .A2(G41), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n294), .A2(G1), .A3(G13), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G41), .ZN(new_n298));
  INV_X1    g0098(.A(G45), .ZN(new_n299));
  AOI21_X1  g0099(.A(G1), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n300), .A2(new_n295), .A3(G274), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT73), .ZN(new_n302));
  INV_X1    g0102(.A(G274), .ZN(new_n303));
  AND2_X1   g0103(.A1(G1), .A2(G13), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n303), .B1(new_n304), .B2(new_n294), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT73), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n305), .A2(new_n306), .A3(new_n300), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n263), .B1(G41), .B2(G45), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n295), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n302), .A2(new_n307), .B1(G238), .B2(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n277), .B1(new_n297), .B2(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n295), .B1(new_n287), .B2(new_n292), .ZN(new_n313));
  AND3_X1   g0113(.A1(new_n305), .A2(new_n306), .A3(new_n300), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n306), .B1(new_n305), .B2(new_n300), .ZN(new_n315));
  INV_X1    g0115(.A(G238), .ZN(new_n316));
  OAI22_X1  g0116(.A1(new_n314), .A2(new_n315), .B1(new_n316), .B2(new_n309), .ZN(new_n317));
  NOR3_X1   g0117(.A1(new_n313), .A2(new_n317), .A3(KEYINPUT13), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n276), .B(G169), .C1(new_n312), .C2(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(KEYINPUT13), .B1(new_n313), .B2(new_n317), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n291), .B1(new_n284), .B2(new_n286), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n311), .B(new_n277), .C1(new_n321), .C2(new_n295), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n320), .A2(new_n322), .A3(G179), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G169), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n325), .B1(new_n320), .B2(new_n322), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n326), .A2(new_n276), .ZN(new_n327));
  OAI21_X1  g0127(.A(KEYINPUT74), .B1(new_n324), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n320), .A2(new_n322), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(G169), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(KEYINPUT14), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT74), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n331), .A2(new_n332), .A3(new_n323), .A4(new_n319), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n275), .B1(new_n328), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n329), .ZN(new_n335));
  INV_X1    g0135(.A(G200), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G190), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n275), .B1(new_n329), .B2(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n334), .A2(new_n340), .ZN(new_n341));
  XOR2_X1   g0141(.A(KEYINPUT8), .B(G58), .Z(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n264), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n254), .A2(new_n257), .ZN(new_n344));
  OAI22_X1  g0144(.A1(new_n343), .A2(new_n344), .B1(new_n257), .B2(new_n342), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT77), .ZN(new_n346));
  XNOR2_X1  g0146(.A(new_n345), .B(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT7), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n348), .B1(new_n285), .B2(G20), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n279), .A2(new_n281), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n350), .A2(KEYINPUT7), .A3(new_n231), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n349), .A2(new_n351), .A3(KEYINPUT76), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT76), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n353), .B(new_n348), .C1(new_n285), .C2(G20), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n352), .A2(G68), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(G58), .A2(G68), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n231), .B1(new_n229), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n231), .A2(new_n278), .ZN(new_n358));
  INV_X1    g0158(.A(G159), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(KEYINPUT16), .B1(new_n355), .B2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n349), .A2(new_n351), .ZN(new_n364));
  OAI21_X1  g0164(.A(KEYINPUT75), .B1(new_n357), .B2(new_n360), .ZN(new_n365));
  INV_X1    g0165(.A(new_n356), .ZN(new_n366));
  OAI21_X1  g0166(.A(G20), .B1(new_n366), .B2(new_n201), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT75), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n266), .A2(G159), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n364), .A2(G68), .B1(new_n365), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n254), .B1(new_n371), .B2(KEYINPUT16), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n347), .B1(new_n363), .B2(new_n372), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n279), .A2(new_n281), .A3(G226), .A4(G1698), .ZN(new_n374));
  INV_X1    g0174(.A(G87), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n374), .B1(new_n278), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n279), .A2(new_n281), .A3(G223), .A4(new_n288), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT79), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n285), .A2(KEYINPUT79), .A3(G223), .A4(new_n288), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n295), .B1(new_n377), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT80), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n295), .A2(G232), .A3(new_n308), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n384), .B1(new_n301), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n301), .A2(new_n385), .A3(new_n384), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(G200), .B1(new_n383), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n388), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n391), .A2(new_n386), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n376), .B1(new_n380), .B2(new_n381), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n392), .B(G190), .C1(new_n393), .C2(new_n295), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n390), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n373), .A2(new_n395), .A3(KEYINPUT17), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT17), .ZN(new_n397));
  XNOR2_X1  g0197(.A(new_n345), .B(KEYINPUT77), .ZN(new_n398));
  NOR3_X1   g0198(.A1(new_n285), .A2(new_n348), .A3(G20), .ZN(new_n399));
  AOI21_X1  g0199(.A(KEYINPUT7), .B1(new_n350), .B2(new_n231), .ZN(new_n400));
  OAI21_X1  g0200(.A(G68), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n365), .A2(new_n370), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT16), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n253), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n398), .B1(new_n405), .B2(new_n362), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n390), .A2(new_n394), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n397), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n396), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT78), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n406), .A2(new_n411), .ZN(new_n412));
  OAI211_X1 g0212(.A(KEYINPUT78), .B(new_n398), .C1(new_n405), .C2(new_n362), .ZN(new_n413));
  OAI21_X1  g0213(.A(G169), .B1(new_n383), .B2(new_n389), .ZN(new_n414));
  INV_X1    g0214(.A(G179), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n392), .B1(new_n393), .B2(new_n295), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n414), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  XNOR2_X1  g0217(.A(KEYINPUT81), .B(KEYINPUT18), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n412), .A2(new_n413), .A3(new_n417), .A4(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n412), .A2(new_n413), .A3(new_n417), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT18), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n421), .A2(KEYINPUT81), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  AND3_X1   g0223(.A1(new_n410), .A2(new_n419), .A3(new_n423), .ZN(new_n424));
  XNOR2_X1  g0224(.A(KEYINPUT8), .B(G58), .ZN(new_n425));
  INV_X1    g0225(.A(G150), .ZN(new_n426));
  OAI22_X1  g0226(.A1(new_n425), .A2(new_n268), .B1(new_n426), .B2(new_n358), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n427), .B1(G20), .B2(new_n203), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n428), .A2(new_n254), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n260), .A2(new_n253), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n430), .A2(G50), .A3(new_n264), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n431), .B1(G50), .B2(new_n257), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NOR3_X1   g0234(.A1(new_n350), .A2(KEYINPUT68), .A3(new_n288), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT68), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n436), .B1(new_n285), .B2(G1698), .ZN(new_n437));
  OAI21_X1  g0237(.A(G223), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n350), .A2(G1698), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n439), .A2(G222), .B1(G77), .B2(new_n350), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT69), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n438), .A2(KEYINPUT69), .A3(new_n440), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n443), .A2(new_n296), .A3(new_n444), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n310), .A2(G226), .B1(new_n300), .B2(new_n305), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n445), .A2(new_n415), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n445), .A2(new_n446), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n434), .B(new_n447), .C1(new_n449), .C2(G169), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n262), .A2(G77), .A3(new_n264), .ZN(new_n451));
  OAI22_X1  g0251(.A1(new_n425), .A2(new_n358), .B1(new_n231), .B2(new_n212), .ZN(new_n452));
  XNOR2_X1  g0252(.A(KEYINPUT15), .B(G87), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n453), .A2(new_n268), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n253), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n260), .A2(new_n212), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n451), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n301), .B1(new_n211), .B2(new_n309), .ZN(new_n459));
  XNOR2_X1  g0259(.A(new_n459), .B(KEYINPUT70), .ZN(new_n460));
  OAI21_X1  g0260(.A(G238), .B1(new_n435), .B2(new_n437), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n439), .A2(G232), .B1(G107), .B2(new_n350), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n295), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(G200), .B1(new_n460), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT70), .ZN(new_n465));
  XNOR2_X1  g0265(.A(new_n459), .B(new_n465), .ZN(new_n466));
  OAI21_X1  g0266(.A(KEYINPUT68), .B1(new_n350), .B2(new_n288), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n285), .A2(new_n436), .A3(G1698), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n316), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n285), .A2(new_n288), .ZN(new_n470));
  INV_X1    g0270(.A(G107), .ZN(new_n471));
  OAI22_X1  g0271(.A1(new_n470), .A2(new_n236), .B1(new_n471), .B2(new_n285), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n296), .B1(new_n469), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n466), .A2(G190), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n458), .A2(new_n464), .A3(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n325), .B1(new_n460), .B2(new_n463), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n466), .A2(new_n415), .A3(new_n473), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n476), .A2(new_n477), .A3(new_n457), .ZN(new_n478));
  AND2_X1   g0278(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n450), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n448), .A2(G200), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT9), .ZN(new_n482));
  XNOR2_X1  g0282(.A(new_n433), .B(new_n482), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n481), .B(new_n483), .C1(new_n338), .C2(new_n448), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT10), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n449), .A2(G190), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT10), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n486), .A2(new_n487), .A3(new_n481), .A4(new_n483), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n480), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n341), .A2(new_n424), .A3(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n257), .A2(G97), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n430), .B1(G1), .B2(new_n278), .ZN(new_n493));
  INV_X1    g0293(.A(G97), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n352), .A2(G107), .A3(new_n354), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n471), .A2(KEYINPUT6), .A3(G97), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n494), .A2(new_n471), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n498), .A2(new_n205), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n497), .B1(new_n499), .B2(KEYINPUT6), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n500), .A2(G20), .B1(G77), .B2(new_n266), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n496), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n495), .B1(new_n502), .B2(new_n253), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT5), .ZN(new_n504));
  OAI21_X1  g0304(.A(KEYINPUT83), .B1(new_n504), .B2(G41), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT83), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n506), .A2(new_n298), .A3(KEYINPUT5), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n504), .A2(G41), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n299), .A2(G1), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n505), .A2(new_n507), .A3(new_n508), .A4(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n295), .A2(G274), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT84), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n263), .B(G45), .C1(new_n298), .C2(KEYINPUT5), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n504), .A2(G41), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n295), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(G257), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n513), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n298), .A2(KEYINPUT5), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n509), .A2(new_n519), .A3(new_n508), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n520), .A2(KEYINPUT84), .A3(G257), .A4(new_n295), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n512), .B1(new_n518), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(G33), .A2(G283), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n279), .A2(new_n281), .A3(G250), .A4(G1698), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n279), .A2(new_n281), .A3(G244), .A4(new_n288), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT4), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n523), .B(new_n524), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n526), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(KEYINPUT82), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT82), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n525), .A2(new_n530), .A3(new_n526), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n527), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n522), .B(G190), .C1(new_n532), .C2(new_n295), .ZN(new_n533));
  AND2_X1   g0333(.A1(new_n503), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n522), .B1(new_n532), .B2(new_n295), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT85), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT85), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n522), .B(new_n537), .C1(new_n532), .C2(new_n295), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n536), .A2(G200), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n534), .A2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n503), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n535), .A2(new_n325), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n522), .B(new_n415), .C1(new_n532), .C2(new_n295), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  AOI211_X1 g0344(.A(new_n253), .B(new_n260), .C1(new_n263), .C2(G33), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(G87), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n285), .A2(new_n231), .A3(G68), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT19), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n231), .B1(new_n290), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(G87), .B2(new_n206), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n548), .B1(new_n268), .B2(new_n494), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n547), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n253), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n453), .A2(new_n260), .ZN(new_n554));
  AND3_X1   g0354(.A1(new_n546), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n279), .A2(new_n281), .A3(G244), .A4(G1698), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n279), .A2(new_n281), .A3(G238), .A4(new_n288), .ZN(new_n557));
  NAND2_X1  g0357(.A1(G33), .A2(G116), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n296), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n509), .A2(new_n303), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n561), .B(new_n295), .C1(G250), .C2(new_n509), .ZN(new_n562));
  AND2_X1   g0362(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(G190), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n560), .A2(new_n562), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(G200), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n555), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n553), .B(new_n554), .C1(new_n453), .C2(new_n493), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n565), .A2(new_n325), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n568), .B(new_n569), .C1(G179), .C2(new_n565), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n540), .A2(new_n544), .A3(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(G116), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n574), .B1(new_n263), .B2(G33), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n259), .A2(new_n261), .A3(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n256), .A2(G20), .A3(new_n574), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n252), .A2(new_n232), .B1(G20), .B2(new_n574), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n523), .B(new_n231), .C1(G33), .C2(new_n494), .ZN(new_n579));
  AOI21_X1  g0379(.A(KEYINPUT20), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n578), .A2(KEYINPUT20), .A3(new_n579), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n576), .B(new_n577), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n279), .A2(new_n281), .A3(G264), .A4(G1698), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT86), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n285), .A2(KEYINPUT86), .A3(G264), .A4(G1698), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n279), .A2(new_n281), .A3(G257), .ZN(new_n588));
  INV_X1    g0388(.A(G303), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(KEYINPUT87), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT87), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(G303), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n588), .A2(new_n288), .B1(new_n350), .B2(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n295), .B1(new_n587), .B2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(G270), .ZN(new_n596));
  OAI22_X1  g0396(.A1(new_n516), .A2(new_n596), .B1(new_n510), .B2(new_n511), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n582), .B(G169), .C1(new_n595), .C2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT21), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n597), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n279), .A2(new_n281), .A3(G257), .A4(new_n288), .ZN(new_n602));
  XNOR2_X1  g0402(.A(KEYINPUT87), .B(G303), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n602), .B1(new_n285), .B2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n604), .B1(new_n585), .B2(new_n586), .ZN(new_n605));
  OAI211_X1 g0405(.A(G190), .B(new_n601), .C1(new_n605), .C2(new_n295), .ZN(new_n606));
  INV_X1    g0406(.A(new_n582), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n587), .A2(new_n594), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n597), .B1(new_n608), .B2(new_n296), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n606), .B(new_n607), .C1(new_n336), .C2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n609), .A2(G179), .A3(new_n582), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n601), .B1(new_n605), .B2(new_n295), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n612), .A2(KEYINPUT21), .A3(G169), .A4(new_n582), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n600), .A2(new_n610), .A3(new_n611), .A4(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT24), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n279), .A2(new_n281), .A3(new_n231), .A4(G87), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(KEYINPUT22), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT22), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n285), .A2(new_n618), .A3(new_n231), .A4(G87), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n558), .A2(G20), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT23), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n622), .B1(new_n231), .B2(G107), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n471), .A2(KEYINPUT23), .A3(G20), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n621), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n615), .B1(new_n620), .B2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n620), .A2(new_n615), .A3(new_n625), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n254), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n260), .A2(KEYINPUT25), .A3(new_n471), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT25), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n631), .B1(new_n257), .B2(G107), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n545), .A2(G107), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  OAI211_X1 g0434(.A(G264), .B(new_n295), .C1(new_n514), .C2(new_n515), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n635), .B1(new_n511), .B2(new_n510), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n279), .A2(new_n281), .A3(G257), .A4(G1698), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n279), .A2(new_n281), .A3(G250), .A4(new_n288), .ZN(new_n638));
  NAND2_X1  g0438(.A1(G33), .A2(G294), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n296), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n636), .B1(new_n641), .B2(KEYINPUT88), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT88), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n640), .A2(new_n643), .A3(new_n296), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n325), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n512), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n641), .A2(new_n646), .A3(new_n635), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n647), .A2(new_n415), .ZN(new_n648));
  OAI22_X1  g0448(.A1(new_n629), .A2(new_n634), .B1(new_n645), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n641), .A2(KEYINPUT88), .ZN(new_n650));
  INV_X1    g0450(.A(new_n636), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n650), .A2(new_n338), .A3(new_n644), .A4(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n647), .A2(new_n336), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n628), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n253), .B1(new_n655), .B2(new_n626), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n654), .A2(new_n656), .A3(new_n633), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n649), .A2(new_n657), .ZN(new_n658));
  NOR4_X1   g0458(.A1(new_n490), .A2(new_n573), .A3(new_n614), .A4(new_n658), .ZN(G372));
  INV_X1    g0459(.A(new_n450), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n485), .A2(KEYINPUT92), .A3(new_n488), .ZN(new_n661));
  AOI21_X1  g0461(.A(KEYINPUT92), .B1(new_n485), .B2(new_n488), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n478), .A2(KEYINPUT91), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT91), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n476), .A2(new_n477), .A3(new_n665), .A4(new_n457), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n340), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n410), .B1(new_n334), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n417), .A2(new_n406), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n670), .B(new_n421), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n660), .B1(new_n663), .B2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n490), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT26), .ZN(new_n675));
  NOR3_X1   g0475(.A1(new_n544), .A2(new_n571), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT90), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n254), .B1(new_n496), .B2(new_n501), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n543), .B1(new_n678), .B2(new_n495), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n535), .A2(new_n325), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n677), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n541), .A2(KEYINPUT90), .A3(new_n542), .A4(new_n543), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(new_n572), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n676), .B1(new_n683), .B2(new_n675), .ZN(new_n684));
  XOR2_X1   g0484(.A(new_n570), .B(KEYINPUT89), .Z(new_n685));
  NAND3_X1  g0485(.A1(new_n600), .A2(new_n611), .A3(new_n613), .ZN(new_n686));
  INV_X1    g0486(.A(new_n645), .ZN(new_n687));
  INV_X1    g0487(.A(new_n648), .ZN(new_n688));
  AOI22_X1  g0488(.A1(new_n687), .A2(new_n688), .B1(new_n656), .B2(new_n633), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n657), .B1(new_n686), .B2(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n685), .B1(new_n573), .B2(new_n690), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n684), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n674), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n673), .A2(new_n693), .ZN(G369));
  NAND2_X1  g0494(.A1(new_n256), .A2(new_n231), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n695), .A2(KEYINPUT27), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(KEYINPUT27), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n696), .A2(G213), .A3(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(G343), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n689), .A2(new_n700), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n701), .A2(KEYINPUT93), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(KEYINPUT93), .ZN(new_n703));
  INV_X1    g0503(.A(new_n658), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n700), .B1(new_n629), .B2(new_n634), .ZN(new_n705));
  AOI22_X1  g0505(.A1(new_n702), .A2(new_n703), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n700), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n607), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n686), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n614), .B2(new_n708), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G330), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n706), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n649), .A2(new_n700), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n702), .A2(new_n703), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n704), .A2(new_n705), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n686), .A2(new_n707), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n714), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n713), .A2(new_n720), .ZN(G399));
  INV_X1    g0521(.A(new_n223), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(G41), .ZN(new_n723));
  NOR3_X1   g0523(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n723), .A2(new_n263), .A3(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n230), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n726), .B1(new_n727), .B2(new_n723), .ZN(new_n728));
  XOR2_X1   g0528(.A(new_n728), .B(KEYINPUT28), .Z(new_n729));
  INV_X1    g0529(.A(KEYINPUT29), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n544), .A2(new_n571), .A3(KEYINPUT26), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n731), .B1(new_n683), .B2(KEYINPUT26), .ZN(new_n732));
  INV_X1    g0532(.A(new_n679), .ZN(new_n733));
  AOI22_X1  g0533(.A1(new_n539), .A2(new_n534), .B1(new_n733), .B2(new_n542), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n649), .A2(new_n600), .A3(new_n611), .A4(new_n613), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n734), .A2(new_n572), .A3(new_n657), .A4(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n732), .A2(new_n736), .A3(new_n685), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n730), .B1(new_n737), .B2(new_n707), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n730), .B(new_n707), .C1(new_n684), .C2(new_n691), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n658), .A2(new_n614), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n742), .A2(new_n734), .A3(new_n572), .A4(new_n707), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT30), .ZN(new_n744));
  AND4_X1   g0544(.A1(new_n560), .A2(new_n641), .A3(new_n562), .A4(new_n635), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n745), .A2(new_n609), .A3(G179), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n744), .B1(new_n746), .B2(new_n535), .ZN(new_n747));
  INV_X1    g0547(.A(new_n535), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n595), .A2(new_n415), .A3(new_n597), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n748), .A2(KEYINPUT30), .A3(new_n749), .A4(new_n745), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n563), .A2(G179), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n751), .A2(new_n535), .A3(new_n612), .A4(new_n647), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n747), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(KEYINPUT31), .B1(new_n753), .B2(new_n700), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n753), .A2(KEYINPUT31), .A3(new_n700), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n743), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G330), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n741), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n729), .B1(new_n760), .B2(G1), .ZN(G364));
  INV_X1    g0561(.A(new_n711), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n255), .A2(G20), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n263), .B1(new_n763), .B2(G45), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n723), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n762), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n767), .B1(G330), .B2(new_n710), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G13), .A2(G33), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(G20), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n232), .B1(G20), .B2(new_n325), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n722), .A2(new_n285), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n774), .B1(G45), .B2(new_n230), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n775), .B1(G45), .B2(new_n250), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n223), .A2(new_n285), .ZN(new_n777));
  XOR2_X1   g0577(.A(G355), .B(KEYINPUT94), .Z(new_n778));
  OAI22_X1  g0578(.A1(new_n777), .A2(new_n778), .B1(G116), .B2(new_n223), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n773), .B1(new_n776), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(new_n766), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n231), .A2(new_n415), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G200), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n338), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n285), .B1(new_n785), .B2(new_n202), .ZN(new_n786));
  NOR3_X1   g0586(.A1(new_n338), .A2(G179), .A3(G200), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(new_n231), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n783), .A2(G190), .ZN(new_n790));
  AOI22_X1  g0590(.A1(G97), .A2(new_n789), .B1(new_n790), .B2(G68), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n231), .A2(G179), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n792), .A2(new_n338), .A3(G200), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G107), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n792), .A2(G190), .A3(G200), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n791), .B(new_n795), .C1(new_n375), .C2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n782), .ZN(new_n798));
  AOI21_X1  g0598(.A(G200), .B1(new_n798), .B2(KEYINPUT95), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n799), .B1(KEYINPUT95), .B2(new_n798), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(G190), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n786), .B(new_n797), .C1(G77), .C2(new_n801), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n792), .A2(new_n338), .A3(new_n336), .ZN(new_n803));
  OR2_X1    g0603(.A1(new_n803), .A2(KEYINPUT97), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(KEYINPUT97), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(new_n359), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT32), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n800), .A2(new_n338), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n809), .B(KEYINPUT96), .Z(new_n810));
  OAI211_X1 g0610(.A(new_n802), .B(new_n808), .C1(new_n227), .C2(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n350), .B1(new_n796), .B2(new_n589), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT99), .ZN(new_n813));
  AOI22_X1  g0613(.A1(G311), .A2(new_n801), .B1(new_n809), .B2(G322), .ZN(new_n814));
  XNOR2_X1  g0614(.A(KEYINPUT33), .B(G317), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  OR2_X1    g0616(.A1(new_n816), .A2(KEYINPUT100), .ZN(new_n817));
  INV_X1    g0617(.A(new_n790), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n818), .B1(KEYINPUT100), .B2(new_n816), .ZN(new_n819));
  INV_X1    g0619(.A(new_n806), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n817), .A2(new_n819), .B1(new_n820), .B2(G329), .ZN(new_n821));
  XOR2_X1   g0621(.A(KEYINPUT98), .B(G326), .Z(new_n822));
  INV_X1    g0622(.A(G294), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n785), .A2(new_n822), .B1(new_n823), .B2(new_n788), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n824), .B1(G283), .B2(new_n794), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n814), .A2(new_n821), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n811), .B1(new_n813), .B2(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n781), .B1(new_n827), .B2(new_n772), .ZN(new_n828));
  INV_X1    g0628(.A(new_n771), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n828), .B1(new_n710), .B2(new_n829), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n768), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(G396));
  NAND2_X1  g0632(.A1(new_n692), .A2(new_n707), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n664), .A2(new_n457), .A3(new_n666), .A4(new_n700), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n478), .B(new_n475), .C1(new_n458), .C2(new_n707), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n833), .A2(new_n837), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n707), .B(new_n836), .C1(new_n684), .C2(new_n691), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n766), .B1(new_n840), .B2(new_n758), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n758), .B2(new_n840), .ZN(new_n842));
  INV_X1    g0642(.A(new_n772), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n770), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n766), .B1(G77), .B2(new_n844), .ZN(new_n845));
  AOI22_X1  g0645(.A1(G116), .A2(new_n801), .B1(new_n809), .B2(G294), .ZN(new_n846));
  INV_X1    g0646(.A(G283), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n818), .A2(new_n847), .B1(new_n785), .B2(new_n589), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n793), .A2(new_n375), .B1(new_n796), .B2(new_n471), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n820), .A2(G311), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n285), .B1(new_n789), .B2(G97), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n846), .A2(new_n850), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n790), .A2(G150), .B1(new_n784), .B2(G137), .ZN(new_n854));
  INV_X1    g0654(.A(new_n801), .ZN(new_n855));
  INV_X1    g0655(.A(G143), .ZN(new_n856));
  OAI221_X1 g0656(.A(new_n854), .B1(new_n359), .B2(new_n855), .C1(new_n810), .C2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n858), .A2(KEYINPUT34), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n285), .B1(new_n788), .B2(new_n227), .ZN(new_n860));
  OAI22_X1  g0660(.A1(new_n793), .A2(new_n228), .B1(new_n796), .B2(new_n202), .ZN(new_n861));
  AOI211_X1 g0661(.A(new_n860), .B(new_n861), .C1(new_n820), .C2(G132), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT34), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n862), .B1(new_n857), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n853), .B1(new_n859), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n845), .B1(new_n865), .B2(new_n772), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n836), .B2(new_n770), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n842), .A2(new_n867), .ZN(G384));
  NOR2_X1   g0668(.A1(new_n763), .A2(new_n263), .ZN(new_n869));
  INV_X1    g0669(.A(G330), .ZN(new_n870));
  AND3_X1   g0670(.A1(new_n753), .A2(KEYINPUT31), .A3(new_n700), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n871), .A2(new_n754), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n837), .B1(new_n872), .B2(new_n743), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n275), .A2(new_n707), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n275), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n335), .A2(G179), .B1(new_n326), .B2(new_n276), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n332), .B1(new_n877), .B2(new_n331), .ZN(new_n878));
  NOR3_X1   g0678(.A1(new_n324), .A2(KEYINPUT74), .A3(new_n327), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n876), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n340), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n875), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NOR3_X1   g0682(.A1(new_n334), .A2(new_n340), .A3(new_n874), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n873), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n698), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n412), .A2(new_n413), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT37), .B1(new_n373), .B2(new_n395), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n420), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(KEYINPUT102), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT102), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n420), .A2(new_n886), .A3(new_n890), .A4(new_n887), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n406), .A2(new_n407), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n371), .A2(KEYINPUT101), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n404), .B1(new_n371), .B2(KEYINPUT101), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n372), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n398), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n893), .B1(new_n417), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n885), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(KEYINPUT37), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n892), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n409), .B1(new_n420), .B2(new_n422), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n419), .ZN(new_n904));
  INV_X1    g0704(.A(new_n899), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n902), .A2(new_n906), .A3(KEYINPUT38), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT38), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n889), .A2(new_n891), .B1(KEYINPUT37), .B2(new_n900), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n899), .B1(new_n903), .B2(new_n419), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n884), .B1(new_n907), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(KEYINPUT103), .B1(new_n912), .B2(KEYINPUT40), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n757), .A2(new_n836), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n880), .A2(new_n881), .A3(new_n875), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n874), .B1(new_n334), .B2(new_n340), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT38), .B1(new_n902), .B2(new_n906), .ZN(new_n918));
  NOR3_X1   g0718(.A1(new_n909), .A2(new_n910), .A3(new_n908), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT103), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT40), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n913), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n917), .A2(KEYINPUT40), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n886), .B(new_n670), .C1(new_n406), .C2(new_n407), .ZN(new_n927));
  AOI22_X1  g0727(.A1(new_n889), .A2(new_n891), .B1(KEYINPUT37), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n886), .B1(new_n671), .B2(new_n410), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n908), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n907), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n926), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n924), .A2(new_n932), .ZN(new_n933));
  XOR2_X1   g0733(.A(new_n933), .B(KEYINPUT104), .Z(new_n934));
  NAND2_X1  g0734(.A1(new_n674), .A2(new_n757), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n870), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n934), .B2(new_n936), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT39), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n927), .A2(KEYINPUT37), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n892), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n929), .ZN(new_n942));
  AOI21_X1  g0742(.A(KEYINPUT38), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n939), .B1(new_n943), .B2(new_n919), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n880), .A2(new_n700), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n907), .A2(new_n911), .A3(KEYINPUT39), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n671), .A2(new_n885), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n907), .A2(new_n911), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n478), .A2(new_n700), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n839), .A2(new_n951), .B1(new_n915), .B2(new_n916), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n948), .B1(new_n949), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n947), .A2(new_n953), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n669), .A2(new_n671), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n661), .A2(new_n662), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n450), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n683), .A2(KEYINPUT26), .ZN(new_n958));
  INV_X1    g0758(.A(new_n731), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n707), .B1(new_n960), .B2(new_n691), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(KEYINPUT29), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n490), .B1(new_n962), .B2(new_n739), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n957), .A2(new_n963), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n954), .B(new_n964), .Z(new_n965));
  AOI21_X1  g0765(.A(new_n869), .B1(new_n938), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n965), .B2(new_n938), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n500), .A2(KEYINPUT35), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n500), .A2(KEYINPUT35), .ZN(new_n969));
  NOR3_X1   g0769(.A1(new_n232), .A2(new_n231), .A3(new_n574), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT36), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n727), .A2(G77), .A3(new_n356), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(G50), .B2(new_n228), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n974), .A2(G1), .A3(new_n255), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n967), .A2(new_n972), .A3(new_n975), .ZN(G367));
  NOR2_X1   g0776(.A1(new_n555), .A2(new_n707), .ZN(new_n977));
  MUX2_X1   g0777(.A(new_n571), .B(new_n685), .S(new_n977), .Z(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n771), .ZN(new_n979));
  INV_X1    g0779(.A(new_n766), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n774), .A2(new_n242), .ZN(new_n981));
  INV_X1    g0781(.A(new_n773), .ZN(new_n982));
  INV_X1    g0782(.A(new_n453), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n982), .B1(new_n722), .B2(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n980), .B1(new_n981), .B2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(G311), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n350), .B1(new_n785), .B2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(G317), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n796), .A2(new_n574), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n806), .A2(new_n988), .B1(KEYINPUT46), .B2(new_n989), .ZN(new_n990));
  AOI211_X1 g0790(.A(new_n987), .B(new_n990), .C1(KEYINPUT46), .C2(new_n989), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n790), .A2(G294), .B1(new_n794), .B2(G97), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n471), .B2(new_n788), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(G283), .B2(new_n801), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n991), .B(new_n994), .C1(new_n603), .C2(new_n810), .ZN(new_n995));
  AOI22_X1  g0795(.A1(new_n809), .A2(G150), .B1(G68), .B2(new_n789), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT107), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n285), .B1(new_n793), .B2(new_n212), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n998), .A2(KEYINPUT108), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(KEYINPUT108), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n999), .B(new_n1000), .C1(new_n855), .C2(new_n202), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n796), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n790), .A2(G159), .B1(new_n1002), .B2(G58), .ZN(new_n1003));
  INV_X1    g0803(.A(G137), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1003), .B1(new_n856), .B2(new_n785), .C1(new_n806), .C2(new_n1004), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1001), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n995), .B1(new_n997), .B2(new_n1006), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1007), .B(KEYINPUT109), .Z(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT47), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n979), .B(new_n985), .C1(new_n1009), .C2(new_n843), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n734), .B1(new_n503), .B2(new_n707), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n733), .A2(new_n542), .A3(new_n700), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n720), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT45), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n720), .A2(KEYINPUT45), .A3(new_n1013), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT44), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n720), .B2(new_n1013), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n1013), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n706), .A2(new_n718), .ZN(new_n1022));
  OAI211_X1 g0822(.A(KEYINPUT44), .B(new_n1021), .C1(new_n1022), .C2(new_n714), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(KEYINPUT105), .B1(new_n1018), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1018), .A2(new_n1024), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(new_n712), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1018), .A2(new_n713), .A3(new_n1024), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1025), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT105), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1026), .A2(new_n1030), .A3(new_n713), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n706), .A2(new_n718), .ZN(new_n1032));
  AND3_X1   g0832(.A1(new_n1032), .A2(KEYINPUT106), .A3(new_n711), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n711), .B1(new_n1032), .B2(KEYINPUT106), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n717), .A2(new_n719), .ZN(new_n1035));
  OR3_X1    g0835(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1035), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n759), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1031), .A2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n760), .B1(new_n1029), .B2(new_n1039), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n723), .B(KEYINPUT41), .Z(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n765), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT43), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n978), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1022), .A2(new_n1013), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n1046), .A2(KEYINPUT42), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n540), .A2(new_n689), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n700), .B1(new_n1048), .B2(new_n544), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(new_n1046), .B2(KEYINPUT42), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1045), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n978), .A2(new_n1044), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1051), .B(new_n1052), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n713), .A2(new_n1021), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1053), .B(new_n1054), .Z(new_n1055));
  OAI21_X1  g0855(.A(new_n1010), .B1(new_n1043), .B2(new_n1055), .ZN(G387));
  NAND2_X1  g0856(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n706), .A2(new_n771), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n777), .A2(new_n724), .B1(G107), .B2(new_n223), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n239), .A2(new_n299), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT110), .ZN(new_n1061));
  AOI211_X1 g0861(.A(G45), .B(new_n725), .C1(G68), .C2(G77), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n425), .A2(G50), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT50), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n722), .B(new_n285), .C1(new_n1062), .C2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1059), .B1(new_n1061), .B2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n766), .B1(new_n1066), .B2(new_n982), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n788), .A2(new_n453), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n785), .A2(new_n359), .B1(new_n796), .B2(new_n212), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n1068), .B(new_n1069), .C1(new_n342), .C2(new_n790), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n820), .A2(G150), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n350), .B1(new_n794), .B2(G97), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(G50), .A2(new_n809), .B1(new_n801), .B2(G68), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1070), .A2(new_n1071), .A3(new_n1072), .A4(new_n1073), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n790), .A2(G311), .B1(new_n784), .B2(G322), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1075), .B1(new_n603), .B2(new_n855), .C1(new_n810), .C2(new_n988), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT48), .ZN(new_n1077));
  OR2_X1    g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n788), .A2(new_n847), .B1(new_n796), .B2(new_n823), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1078), .A2(KEYINPUT49), .A3(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n285), .B1(new_n794), .B2(G116), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1081), .B(new_n1082), .C1(new_n822), .C2(new_n806), .ZN(new_n1083));
  AOI21_X1  g0883(.A(KEYINPUT49), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1074), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1067), .B1(new_n1085), .B2(new_n772), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n1057), .A2(new_n765), .B1(new_n1058), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1038), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n723), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1057), .A2(new_n760), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1087), .B1(new_n1089), .B2(new_n1090), .ZN(G393));
  INV_X1    g0891(.A(new_n1028), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n713), .B1(new_n1018), .B2(new_n1024), .ZN(new_n1093));
  NOR3_X1   g0893(.A1(new_n1092), .A2(new_n764), .A3(new_n1093), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1013), .A2(new_n829), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT111), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n247), .A2(new_n774), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n982), .B1(new_n722), .B2(G97), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n980), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n809), .A2(G311), .B1(G317), .B2(new_n784), .ZN(new_n1100));
  XOR2_X1   g0900(.A(new_n1100), .B(KEYINPUT52), .Z(new_n1101));
  AOI22_X1  g0901(.A1(new_n789), .A2(G116), .B1(new_n1002), .B2(G283), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n603), .B2(new_n818), .ZN(new_n1103));
  INV_X1    g0903(.A(G322), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n350), .B(new_n795), .C1(new_n806), .C2(new_n1104), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n1103), .B(new_n1105), .C1(G294), .C2(new_n801), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n809), .A2(G159), .B1(G150), .B2(new_n784), .ZN(new_n1107));
  XOR2_X1   g0907(.A(new_n1107), .B(KEYINPUT51), .Z(new_n1108));
  AOI22_X1  g0908(.A1(new_n790), .A2(G50), .B1(new_n1002), .B2(G68), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n212), .B2(new_n788), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n285), .B1(new_n375), .B2(new_n793), .C1(new_n806), .C2(new_n856), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n1110), .B(new_n1111), .C1(new_n342), .C2(new_n801), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n1101), .A2(new_n1106), .B1(new_n1108), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1099), .B1(new_n1113), .B2(new_n843), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1096), .A2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1094), .A2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n723), .B1(new_n1117), .B2(new_n1038), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1029), .A2(new_n1039), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1116), .B1(new_n1118), .B2(new_n1119), .ZN(G390));
  NAND2_X1  g0920(.A1(new_n915), .A2(new_n916), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1121), .A2(G330), .A3(new_n873), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n952), .A2(new_n945), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(new_n944), .B2(new_n946), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n951), .B1(new_n961), .B2(new_n837), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n1121), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n945), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n931), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1123), .B1(new_n1125), .B2(new_n1130), .ZN(new_n1131));
  AND3_X1   g0931(.A1(new_n907), .A2(new_n911), .A3(KEYINPUT39), .ZN(new_n1132));
  AOI21_X1  g0932(.A(KEYINPUT39), .B1(new_n907), .B2(new_n930), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1122), .B(new_n1129), .C1(new_n1134), .C2(new_n1124), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1131), .A2(new_n1135), .A3(new_n765), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n766), .B1(new_n342), .B2(new_n844), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n809), .A2(G132), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n796), .A2(new_n426), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT53), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(KEYINPUT54), .B(G143), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1138), .B(new_n1140), .C1(new_n855), .C2(new_n1141), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(G159), .A2(new_n789), .B1(new_n790), .B2(G137), .ZN(new_n1143));
  INV_X1    g0943(.A(G128), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1143), .B1(new_n1144), .B2(new_n785), .ZN(new_n1145));
  INV_X1    g0945(.A(G125), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n285), .B1(new_n202), .B2(new_n793), .C1(new_n806), .C2(new_n1146), .ZN(new_n1147));
  NOR3_X1   g0947(.A1(new_n1142), .A2(new_n1145), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  OR2_X1    g0949(.A1(new_n1149), .A2(KEYINPUT113), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(G97), .A2(new_n801), .B1(new_n809), .B2(G116), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n818), .A2(new_n471), .B1(new_n785), .B2(new_n847), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n788), .A2(new_n212), .B1(new_n793), .B2(new_n228), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n820), .A2(G294), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n285), .B1(new_n1002), .B2(G87), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1151), .A2(new_n1154), .A3(new_n1155), .A4(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1149), .A2(KEYINPUT113), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1150), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1137), .B1(new_n1159), .B2(new_n772), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1160), .B1(new_n1134), .B2(new_n770), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n674), .B1(new_n738), .B2(new_n740), .ZN(new_n1162));
  OR2_X1    g0962(.A1(new_n490), .A2(new_n758), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1162), .A2(new_n673), .A3(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n757), .A2(G330), .A3(new_n836), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1165), .A2(new_n915), .A3(new_n916), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1122), .A2(new_n1166), .ZN(new_n1167));
  AND2_X1   g0967(.A1(new_n839), .A2(new_n951), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n691), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n700), .B1(new_n1171), .B2(new_n732), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n950), .B1(new_n1172), .B2(new_n836), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1122), .A2(new_n1173), .A3(new_n1166), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1164), .B1(new_n1170), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1131), .A2(new_n1135), .A3(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT112), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1176), .A2(new_n1177), .A3(new_n723), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1131), .A2(new_n1135), .ZN(new_n1179));
  AND3_X1   g0979(.A1(new_n1122), .A2(new_n1173), .A3(new_n1166), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1168), .B1(new_n1122), .B2(new_n1166), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n964), .B(new_n1163), .C1(new_n1180), .C2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1178), .A2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1177), .B1(new_n1176), .B2(new_n723), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1136), .B(new_n1161), .C1(new_n1184), .C2(new_n1185), .ZN(G378));
  NOR2_X1   g0986(.A1(new_n956), .A2(new_n660), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n433), .A2(new_n698), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT116), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(new_n1187), .B(new_n1189), .ZN(new_n1190));
  XOR2_X1   g0990(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1190), .B(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n870), .B1(new_n926), .B2(new_n931), .ZN(new_n1195));
  AND3_X1   g0995(.A1(new_n924), .A2(new_n954), .A3(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n954), .B1(new_n924), .B2(new_n1195), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1194), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1164), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1176), .A2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n921), .B1(new_n920), .B2(new_n922), .ZN(new_n1201));
  AOI211_X1 g1001(.A(KEYINPUT103), .B(KEYINPUT40), .C1(new_n949), .C2(new_n917), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1195), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n954), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n924), .A2(new_n954), .A3(new_n1195), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1205), .A2(new_n1206), .A3(new_n1193), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1198), .A2(new_n1200), .A3(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT57), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1198), .A2(new_n1207), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1200), .A2(KEYINPUT57), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n723), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  OR2_X1    g1013(.A1(new_n1210), .A2(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1198), .A2(new_n765), .A3(new_n1207), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n766), .B1(G50), .B2(new_n844), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n285), .A2(G41), .ZN(new_n1217));
  AOI211_X1 g1017(.A(G50), .B(new_n1217), .C1(new_n278), .C2(new_n298), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n785), .A2(new_n574), .B1(new_n228), .B2(new_n788), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n818), .A2(new_n494), .B1(new_n227), .B2(new_n793), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n1219), .B(new_n1220), .C1(G283), .C2(new_n820), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(G107), .A2(new_n809), .B1(new_n801), .B2(new_n983), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1217), .B1(new_n212), .B2(new_n796), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1223), .B(KEYINPUT114), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1221), .A2(new_n1222), .A3(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT58), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1218), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n790), .A2(G132), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n809), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n1228), .B1(new_n796), .B2(new_n1141), .C1(new_n1229), .C2(new_n1144), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(G150), .A2(new_n789), .B1(new_n784), .B2(G125), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(new_n1231), .B(KEYINPUT115), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n1230), .B(new_n1232), .C1(G137), .C2(new_n801), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1234), .A2(KEYINPUT59), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n820), .A2(G124), .ZN(new_n1236));
  AOI211_X1 g1036(.A(G33), .B(G41), .C1(new_n794), .C2(G159), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT59), .ZN(new_n1238));
  OAI211_X1 g1038(.A(new_n1236), .B(new_n1237), .C1(new_n1233), .C2(new_n1238), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n1227), .B1(new_n1226), .B2(new_n1225), .C1(new_n1235), .C2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1216), .B1(new_n1240), .B2(new_n772), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1241), .B1(new_n1193), .B2(new_n770), .ZN(new_n1242));
  AND2_X1   g1042(.A1(new_n1215), .A2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1214), .A2(new_n1243), .ZN(G375));
  NAND3_X1  g1044(.A1(new_n1170), .A2(new_n1164), .A3(new_n1174), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1182), .A2(new_n1042), .A3(new_n1245), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(new_n1246), .B(KEYINPUT117), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n764), .B1(new_n1170), .B2(new_n1174), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n915), .A2(new_n916), .A3(new_n769), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n766), .B1(G68), .B2(new_n844), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n801), .A2(G107), .B1(G116), .B2(new_n790), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1251), .B(KEYINPUT118), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1068), .B1(G294), .B2(new_n784), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1253), .B1(new_n1229), .B2(new_n847), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n285), .B1(new_n794), .B2(G77), .ZN(new_n1255));
  OR2_X1    g1055(.A1(new_n1255), .A2(KEYINPUT119), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(KEYINPUT119), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1254), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  OAI22_X1  g1058(.A1(new_n806), .A2(new_n589), .B1(new_n494), .B2(new_n796), .ZN(new_n1259));
  XOR2_X1   g1059(.A(new_n1259), .B(KEYINPUT120), .Z(new_n1260));
  NAND3_X1  g1060(.A1(new_n1252), .A2(new_n1258), .A3(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT121), .ZN(new_n1262));
  OR2_X1    g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  OAI22_X1  g1063(.A1(new_n818), .A2(new_n1141), .B1(new_n359), .B2(new_n796), .ZN(new_n1264));
  OAI221_X1 g1064(.A(new_n285), .B1(new_n227), .B2(new_n793), .C1(new_n806), .C2(new_n1144), .ZN(new_n1265));
  AOI211_X1 g1065(.A(new_n1264), .B(new_n1265), .C1(G132), .C2(new_n784), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n801), .A2(G150), .B1(G50), .B2(new_n789), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1267), .B(KEYINPUT122), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1266), .B(new_n1268), .C1(new_n1004), .C2(new_n810), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1263), .A2(new_n1269), .A3(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1250), .B1(new_n1271), .B2(new_n772), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1248), .B1(new_n1249), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1247), .A2(new_n1273), .ZN(new_n1274));
  XNOR2_X1  g1074(.A(new_n1274), .B(KEYINPUT123), .ZN(G381));
  OR2_X1    g1075(.A1(G393), .A2(G396), .ZN(new_n1276));
  OR4_X1    g1076(.A1(G384), .A2(G387), .A3(G390), .A4(new_n1276), .ZN(new_n1277));
  OR4_X1    g1077(.A1(G378), .A2(new_n1277), .A3(G375), .A4(G381), .ZN(G407));
  INV_X1    g1078(.A(G378), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n699), .A2(G213), .ZN(new_n1280));
  XOR2_X1   g1080(.A(new_n1280), .B(KEYINPUT124), .Z(new_n1281));
  NAND4_X1  g1081(.A1(new_n1214), .A2(new_n1279), .A3(new_n1243), .A4(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(G407), .A2(G213), .A3(new_n1282), .ZN(G409));
  OAI211_X1 g1083(.A(G378), .B(new_n1243), .C1(new_n1210), .C2(new_n1213), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1215), .B(new_n1242), .C1(new_n1208), .C2(new_n1041), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1279), .A2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1284), .A2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT60), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1245), .A2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n723), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1288), .B1(new_n1182), .B2(new_n1245), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1273), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(G384), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  OAI211_X1 g1094(.A(G384), .B(new_n1273), .C1(new_n1290), .C2(new_n1291), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1287), .A2(new_n1280), .A3(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT63), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT126), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n699), .A2(G213), .A3(G2897), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1294), .A2(new_n1295), .A3(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(KEYINPUT125), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT125), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1294), .A2(new_n1305), .A3(new_n1295), .A4(new_n1302), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1304), .A2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1281), .A2(G2897), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1308), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1301), .B1(new_n1307), .B2(new_n1310), .ZN(new_n1311));
  AOI211_X1 g1111(.A(KEYINPUT126), .B(new_n1309), .C1(new_n1304), .C2(new_n1306), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1287), .A2(new_n1280), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1281), .B1(new_n1284), .B2(new_n1286), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1316), .A2(KEYINPUT63), .A3(new_n1297), .ZN(new_n1317));
  INV_X1    g1117(.A(G390), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(G387), .A2(new_n1318), .ZN(new_n1319));
  XNOR2_X1  g1119(.A(G393), .B(new_n831), .ZN(new_n1320));
  OAI211_X1 g1120(.A(G390), .B(new_n1010), .C1(new_n1043), .C2(new_n1055), .ZN(new_n1321));
  AND3_X1   g1121(.A1(new_n1319), .A2(new_n1320), .A3(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1320), .B1(new_n1319), .B2(new_n1321), .ZN(new_n1323));
  NOR3_X1   g1123(.A1(new_n1322), .A2(new_n1323), .A3(KEYINPUT61), .ZN(new_n1324));
  NAND4_X1  g1124(.A1(new_n1300), .A2(new_n1315), .A3(new_n1317), .A4(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT61), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1307), .A2(new_n1310), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1326), .B1(new_n1316), .B2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT62), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1298), .A2(new_n1329), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1316), .A2(KEYINPUT62), .A3(new_n1297), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1328), .B1(new_n1330), .B2(new_n1331), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1325), .B1(new_n1332), .B2(new_n1333), .ZN(G405));
  INV_X1    g1134(.A(KEYINPUT127), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1297), .A2(new_n1335), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1336), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1320), .ZN(new_n1338));
  XNOR2_X1  g1138(.A(new_n1053), .B(new_n1054), .ZN(new_n1339));
  AND2_X1   g1139(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1339), .B1(new_n1340), .B2(new_n765), .ZN(new_n1341));
  AOI21_X1  g1141(.A(G390), .B1(new_n1341), .B2(new_n1010), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1321), .ZN(new_n1343));
  OAI21_X1  g1143(.A(new_n1338), .B1(new_n1342), .B2(new_n1343), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1319), .A2(new_n1320), .A3(new_n1321), .ZN(new_n1345));
  INV_X1    g1145(.A(new_n1336), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1344), .A2(new_n1345), .A3(new_n1346), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1337), .A2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(G375), .A2(new_n1279), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1297), .A2(new_n1335), .ZN(new_n1350));
  AND2_X1   g1150(.A1(new_n1284), .A2(new_n1350), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1349), .A2(new_n1351), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1348), .A2(new_n1352), .ZN(new_n1353));
  NAND4_X1  g1153(.A1(new_n1337), .A2(new_n1347), .A3(new_n1349), .A4(new_n1351), .ZN(new_n1354));
  AND2_X1   g1154(.A1(new_n1353), .A2(new_n1354), .ZN(G402));
endmodule


