//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 0 0 1 0 0 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 1 1 0 0 0 1 0 0 1 1 1 0 0 1 1 0 1 1 1 0 0 0 1 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:45 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1268, new_n1269, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1336, new_n1337, new_n1338;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  INV_X1    g0014(.A(new_n201), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G50), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(new_n211), .A2(new_n212), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT64), .Z(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n209), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n218), .B1(new_n212), .B2(new_n211), .C1(new_n225), .C2(KEYINPUT1), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XOR2_X1   g0027(.A(G238), .B(G244), .Z(new_n228));
  XNOR2_X1  g0028(.A(G226), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT66), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(G41), .ZN(new_n245));
  INV_X1    g0045(.A(G45), .ZN(new_n246));
  AOI21_X1  g0046(.A(G1), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(G274), .ZN(new_n248));
  INV_X1    g0048(.A(new_n247), .ZN(new_n249));
  INV_X1    g0049(.A(new_n213), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G33), .A2(G41), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G238), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n248), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  OR2_X1    g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  AOI21_X1  g0057(.A(G1698), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(KEYINPUT73), .A3(G226), .ZN(new_n259));
  INV_X1    g0059(.A(G1698), .ZN(new_n260));
  AND2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  OAI211_X1 g0062(.A(G226), .B(new_n260), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT73), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(G33), .A2(G97), .ZN(new_n266));
  OAI211_X1 g0066(.A(G232), .B(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n267));
  NAND4_X1  g0067(.A1(new_n259), .A2(new_n265), .A3(new_n266), .A4(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n255), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT13), .ZN(new_n271));
  OAI21_X1  g0071(.A(KEYINPUT74), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  OAI211_X1 g0072(.A(new_n266), .B(new_n267), .C1(new_n263), .C2(new_n264), .ZN(new_n273));
  AOI21_X1  g0073(.A(KEYINPUT73), .B1(new_n258), .B2(G226), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n269), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n255), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT74), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n277), .A2(new_n278), .A3(KEYINPUT13), .ZN(new_n279));
  AOI22_X1  g0079(.A1(new_n272), .A2(new_n279), .B1(new_n271), .B2(new_n270), .ZN(new_n280));
  INV_X1    g0080(.A(G169), .ZN(new_n281));
  OAI21_X1  g0081(.A(KEYINPUT14), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n270), .A2(new_n271), .ZN(new_n283));
  NOR3_X1   g0083(.A1(new_n270), .A2(KEYINPUT74), .A3(new_n271), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n278), .B1(new_n277), .B2(KEYINPUT13), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT14), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n286), .A2(new_n287), .A3(G169), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n277), .A2(KEYINPUT13), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n289), .A2(new_n283), .A3(G179), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n282), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n213), .ZN(new_n293));
  INV_X1    g0093(.A(G33), .ZN(new_n294));
  OAI21_X1  g0094(.A(KEYINPUT67), .B1(new_n294), .B2(G20), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT67), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n296), .A2(new_n207), .A3(G33), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n295), .A2(new_n297), .A3(G77), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n298), .B1(new_n207), .B2(G68), .ZN(new_n299));
  NOR2_X1   g0099(.A1(G20), .A2(G33), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  OAI22_X1  g0101(.A1(new_n299), .A2(KEYINPUT75), .B1(new_n202), .B2(new_n301), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n299), .A2(KEYINPUT75), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n293), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT11), .ZN(new_n305));
  OR2_X1    g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(new_n305), .ZN(new_n307));
  AND2_X1   g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G13), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n309), .A2(G1), .ZN(new_n310));
  INV_X1    g0110(.A(G68), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n310), .A2(G20), .A3(new_n311), .ZN(new_n312));
  XNOR2_X1  g0112(.A(new_n312), .B(KEYINPUT12), .ZN(new_n313));
  INV_X1    g0113(.A(new_n293), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n314), .A2(KEYINPUT70), .A3(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT70), .ZN(new_n317));
  INV_X1    g0117(.A(new_n315), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n317), .B1(new_n318), .B2(new_n293), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n206), .A2(G20), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n316), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n313), .B1(new_n321), .B2(new_n311), .ZN(new_n322));
  XNOR2_X1  g0122(.A(new_n322), .B(KEYINPUT76), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n308), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n291), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n314), .A2(new_n315), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n320), .A2(G50), .ZN(new_n327));
  OAI22_X1  g0127(.A1(new_n326), .A2(new_n327), .B1(G50), .B2(new_n315), .ZN(new_n328));
  INV_X1    g0128(.A(G58), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT8), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT8), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G58), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n333), .A2(new_n295), .A3(new_n297), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n300), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n314), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n328), .A2(new_n336), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n261), .A2(new_n262), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n258), .A2(G222), .B1(new_n338), .B2(G77), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n260), .B1(new_n256), .B2(new_n257), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G223), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n252), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(G226), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n248), .B1(new_n253), .B2(new_n343), .ZN(new_n344));
  OR2_X1    g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(G169), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n342), .A2(new_n344), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(G179), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n337), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(G77), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n318), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n351), .B1(new_n321), .B2(new_n350), .ZN(new_n352));
  XNOR2_X1  g0152(.A(KEYINPUT15), .B(G87), .ZN(new_n353));
  NOR3_X1   g0153(.A1(new_n353), .A2(G20), .A3(new_n294), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n207), .A2(new_n350), .ZN(new_n355));
  OR2_X1    g0155(.A1(new_n300), .A2(KEYINPUT68), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n300), .A2(KEYINPUT68), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n355), .B1(new_n358), .B2(new_n333), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n354), .B1(new_n359), .B2(KEYINPUT69), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT69), .ZN(new_n361));
  INV_X1    g0161(.A(new_n333), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n362), .B1(new_n356), .B2(new_n357), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n361), .B1(new_n363), .B2(new_n355), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n352), .B1(new_n365), .B2(new_n293), .ZN(new_n366));
  INV_X1    g0166(.A(G244), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n248), .B1(new_n253), .B2(new_n367), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n258), .A2(G232), .B1(new_n338), .B2(G107), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n340), .A2(G238), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI211_X1 g0171(.A(G190), .B(new_n368), .C1(new_n371), .C2(new_n269), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n269), .ZN(new_n373));
  INV_X1    g0173(.A(new_n368), .ZN(new_n374));
  AOI21_X1  g0174(.A(G200), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n366), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(G179), .ZN(new_n377));
  AOI211_X1 g0177(.A(new_n377), .B(new_n368), .C1(new_n371), .C2(new_n269), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n281), .B1(new_n373), .B2(new_n374), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n314), .B1(new_n360), .B2(new_n364), .ZN(new_n380));
  OAI22_X1  g0180(.A1(new_n378), .A2(new_n379), .B1(new_n380), .B2(new_n352), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n376), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT72), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n345), .A2(new_n383), .A3(G200), .ZN(new_n384));
  INV_X1    g0184(.A(G200), .ZN(new_n385));
  OAI21_X1  g0185(.A(KEYINPUT72), .B1(new_n347), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT71), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n389), .B1(new_n337), .B2(KEYINPUT9), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT9), .ZN(new_n391));
  NOR4_X1   g0191(.A1(new_n328), .A2(new_n336), .A3(KEYINPUT71), .A4(new_n391), .ZN(new_n392));
  OR2_X1    g0192(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT10), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n347), .A2(G190), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n391), .B1(new_n336), .B2(new_n328), .ZN(new_n396));
  AND2_X1   g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n388), .A2(new_n393), .A3(new_n394), .A4(new_n397), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n395), .B(new_n396), .C1(new_n390), .C2(new_n392), .ZN(new_n399));
  OAI21_X1  g0199(.A(KEYINPUT10), .B1(new_n387), .B2(new_n399), .ZN(new_n400));
  AOI211_X1 g0200(.A(new_n349), .B(new_n382), .C1(new_n398), .C2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n286), .A2(G200), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n289), .A2(new_n283), .A3(G190), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n402), .A2(new_n323), .A3(new_n308), .A4(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n333), .A2(new_n320), .ZN(new_n405));
  OAI22_X1  g0205(.A1(new_n326), .A2(new_n405), .B1(new_n315), .B2(new_n333), .ZN(new_n406));
  AOI21_X1  g0206(.A(KEYINPUT7), .B1(new_n338), .B2(new_n207), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT7), .ZN(new_n408));
  NOR4_X1   g0208(.A1(new_n261), .A2(new_n262), .A3(new_n408), .A4(G20), .ZN(new_n409));
  OAI21_X1  g0209(.A(G68), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n329), .A2(new_n311), .ZN(new_n411));
  OAI21_X1  g0211(.A(G20), .B1(new_n411), .B2(new_n201), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n300), .A2(G159), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n410), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT16), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n314), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n256), .A2(KEYINPUT77), .A3(new_n257), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT77), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(new_n261), .B2(new_n262), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n419), .A2(new_n421), .A3(new_n207), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n409), .B1(new_n422), .B2(new_n408), .ZN(new_n423));
  OAI211_X1 g0223(.A(KEYINPUT16), .B(new_n415), .C1(new_n423), .C2(new_n311), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n406), .B1(new_n418), .B2(new_n424), .ZN(new_n425));
  OAI211_X1 g0225(.A(G226), .B(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT79), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(G33), .A2(G87), .ZN(new_n430));
  OAI211_X1 g0230(.A(G223), .B(new_n260), .C1(new_n261), .C2(new_n262), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n430), .B(new_n431), .C1(new_n426), .C2(new_n427), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n269), .B1(new_n429), .B2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(G190), .ZN(new_n434));
  INV_X1    g0234(.A(G232), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n248), .B1(new_n253), .B2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n433), .A2(new_n434), .A3(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n340), .A2(KEYINPUT79), .A3(G226), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n439), .A2(new_n428), .A3(new_n430), .A4(new_n431), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n436), .B1(new_n440), .B2(new_n269), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n438), .B1(new_n441), .B2(G200), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n425), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT17), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n425), .A2(KEYINPUT17), .A3(new_n442), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n256), .A2(new_n257), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n408), .B1(new_n448), .B2(G20), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n338), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n311), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n417), .B1(new_n451), .B2(new_n414), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n424), .A2(new_n293), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n406), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(KEYINPUT78), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT78), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n425), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n433), .A2(new_n377), .A3(new_n437), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n459), .B1(new_n441), .B2(G169), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n456), .A2(new_n458), .A3(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT18), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n456), .A2(new_n458), .A3(KEYINPUT18), .A4(new_n461), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n447), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AND4_X1   g0266(.A1(new_n325), .A2(new_n401), .A3(new_n404), .A4(new_n466), .ZN(new_n467));
  OAI211_X1 g0267(.A(G250), .B(new_n260), .C1(new_n261), .C2(new_n262), .ZN(new_n468));
  OAI211_X1 g0268(.A(G257), .B(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n469));
  INV_X1    g0269(.A(G294), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n468), .B(new_n469), .C1(new_n294), .C2(new_n470), .ZN(new_n471));
  XNOR2_X1  g0271(.A(KEYINPUT5), .B(G41), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n246), .A2(G1), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n472), .A2(new_n473), .B1(new_n250), .B2(new_n251), .ZN(new_n474));
  AOI22_X1  g0274(.A1(new_n471), .A2(new_n269), .B1(G264), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n206), .A2(G45), .ZN(new_n476));
  OR2_X1    g0276(.A1(KEYINPUT5), .A2(G41), .ZN(new_n477));
  NAND2_X1  g0277(.A1(KEYINPUT5), .A2(G41), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(G274), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n475), .A2(new_n434), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(G200), .B1(new_n475), .B2(new_n480), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n206), .A2(G33), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n315), .A2(new_n484), .A3(new_n213), .A4(new_n292), .ZN(new_n485));
  AND2_X1   g0285(.A1(new_n485), .A2(KEYINPUT81), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n485), .A2(KEYINPUT81), .ZN(new_n487));
  OAI21_X1  g0287(.A(G107), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(G107), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n310), .A2(G20), .A3(new_n489), .ZN(new_n490));
  XOR2_X1   g0290(.A(new_n490), .B(KEYINPUT25), .Z(new_n491));
  OAI211_X1 g0291(.A(new_n207), .B(G87), .C1(new_n261), .C2(new_n262), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT22), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT22), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n448), .A2(new_n494), .A3(new_n207), .A4(G87), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT23), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n497), .B1(new_n207), .B2(G107), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n489), .A2(KEYINPUT23), .A3(G20), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(G33), .A2(G116), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n500), .B1(G20), .B2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n496), .A2(new_n503), .A3(KEYINPUT24), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n293), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n502), .B1(new_n493), .B2(new_n495), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n506), .A2(KEYINPUT24), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n488), .B(new_n491), .C1(new_n505), .C2(new_n507), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n483), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT89), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n475), .A2(new_n377), .A3(new_n480), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(G169), .B1(new_n475), .B2(new_n480), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n510), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n471), .A2(new_n269), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n474), .A2(G264), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n515), .A2(new_n516), .A3(new_n480), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n281), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n518), .A2(KEYINPUT89), .A3(new_n511), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n514), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n509), .B1(new_n520), .B2(new_n508), .ZN(new_n521));
  OAI211_X1 g0321(.A(G238), .B(new_n260), .C1(new_n261), .C2(new_n262), .ZN(new_n522));
  OAI211_X1 g0322(.A(G244), .B(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n522), .A2(new_n523), .A3(new_n501), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n269), .ZN(new_n525));
  NAND2_X1  g0325(.A1(KEYINPUT83), .A2(G250), .ZN(new_n526));
  INV_X1    g0326(.A(G274), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n473), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT83), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n476), .A2(new_n530), .A3(G250), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n269), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n525), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(G200), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n532), .B1(new_n524), .B2(new_n269), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G190), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n448), .A2(new_n207), .A3(G68), .ZN(new_n538));
  INV_X1    g0338(.A(G87), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(KEYINPUT85), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT85), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(G87), .ZN(new_n542));
  NOR2_X1   g0342(.A1(G97), .A2(G107), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n540), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT19), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n207), .B1(new_n266), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n545), .B1(new_n266), .B2(G20), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n538), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n549), .A2(new_n293), .B1(new_n318), .B2(new_n353), .ZN(new_n550));
  XNOR2_X1  g0350(.A(new_n485), .B(KEYINPUT81), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(G87), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n535), .A2(new_n537), .A3(new_n550), .A4(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n534), .A2(new_n281), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT86), .ZN(new_n555));
  XNOR2_X1  g0355(.A(new_n353), .B(new_n555), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n556), .B(KEYINPUT87), .C1(new_n486), .C2(new_n487), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n550), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(KEYINPUT87), .B1(new_n551), .B2(new_n556), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n554), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT84), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n536), .A2(new_n561), .A3(new_n377), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n561), .B1(new_n536), .B2(new_n377), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n553), .B1(new_n560), .B2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n474), .A2(G270), .B1(G274), .B2(new_n479), .ZN(new_n567));
  OAI211_X1 g0367(.A(G264), .B(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n568));
  OAI211_X1 g0368(.A(G257), .B(new_n260), .C1(new_n261), .C2(new_n262), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n256), .A2(G303), .A3(new_n257), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n269), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n567), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(G200), .ZN(new_n574));
  NAND2_X1  g0374(.A1(G33), .A2(G283), .ZN(new_n575));
  INV_X1    g0375(.A(G97), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n575), .B1(new_n576), .B2(G33), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n207), .ZN(new_n578));
  INV_X1    g0378(.A(G116), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n207), .A2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(KEYINPUT20), .B1(new_n582), .B2(new_n293), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n580), .B1(new_n577), .B2(new_n207), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT20), .ZN(new_n585));
  NOR3_X1   g0385(.A1(new_n584), .A2(new_n585), .A3(new_n314), .ZN(new_n586));
  OR2_X1    g0386(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n316), .A2(new_n319), .A3(G116), .A4(new_n484), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n318), .A2(new_n579), .ZN(new_n589));
  AND2_X1   g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n574), .A2(new_n587), .A3(KEYINPUT88), .A4(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT88), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n588), .B(new_n589), .C1(new_n583), .C2(new_n586), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n385), .B1(new_n567), .B2(new_n572), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n567), .A2(new_n572), .A3(G190), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n591), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n571), .A2(new_n269), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n472), .A2(new_n473), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n599), .A2(G270), .A3(new_n252), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n480), .ZN(new_n601));
  OAI211_X1 g0401(.A(KEYINPUT21), .B(G169), .C1(new_n598), .C2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n567), .A2(new_n572), .A3(G179), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n281), .B1(new_n567), .B2(new_n572), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n593), .A2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT21), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n604), .A2(new_n593), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(G97), .B1(new_n486), .B2(new_n487), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(G97), .B2(new_n315), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT6), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n576), .A2(new_n489), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n611), .B1(new_n612), .B2(new_n543), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT80), .ZN(new_n614));
  NAND2_X1  g0414(.A1(KEYINPUT6), .A2(G97), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n614), .B1(new_n615), .B2(G107), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n489), .A2(KEYINPUT80), .A3(KEYINPUT6), .A4(G97), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n207), .B1(new_n613), .B2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(G107), .B1(new_n407), .B2(new_n409), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n620), .B(new_n621), .C1(new_n350), .C2(new_n301), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n610), .B1(new_n293), .B2(new_n622), .ZN(new_n623));
  OAI211_X1 g0423(.A(G250), .B(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n624));
  OAI211_X1 g0424(.A(G244), .B(new_n260), .C1(new_n261), .C2(new_n262), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT4), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(KEYINPUT82), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n575), .B(new_n624), .C1(new_n625), .C2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n627), .B1(new_n258), .B2(G244), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n269), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n599), .A2(G257), .A3(new_n252), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n632), .A2(new_n480), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n631), .A2(new_n633), .A3(new_n434), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n632), .A2(new_n480), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n258), .A2(G244), .A3(new_n627), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n625), .A2(new_n628), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n636), .A2(new_n637), .A3(new_n575), .A4(new_n624), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n635), .B1(new_n638), .B2(new_n269), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n634), .B1(new_n639), .B2(G200), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n623), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n315), .A2(G97), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n642), .B1(new_n551), .B2(G97), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n489), .B1(new_n449), .B2(new_n450), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n301), .A2(new_n350), .ZN(new_n645));
  NOR3_X1   g0445(.A1(new_n644), .A2(new_n619), .A3(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n643), .B1(new_n646), .B2(new_n314), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n631), .A2(new_n633), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n648), .A2(new_n377), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n281), .B1(new_n631), .B2(new_n633), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n647), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  AND4_X1   g0451(.A1(new_n597), .A2(new_n608), .A3(new_n641), .A4(new_n651), .ZN(new_n652));
  AND4_X1   g0452(.A1(new_n467), .A2(new_n521), .A3(new_n566), .A4(new_n652), .ZN(G372));
  NAND2_X1  g0453(.A1(new_n550), .A2(new_n552), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n536), .A2(new_n385), .ZN(new_n655));
  OAI21_X1  g0455(.A(KEYINPUT90), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT90), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n535), .A2(new_n657), .A3(new_n550), .A4(new_n552), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n656), .A2(new_n537), .A3(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT26), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(new_n660), .A3(new_n641), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n488), .A2(new_n491), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n506), .A2(KEYINPUT24), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n314), .B1(new_n506), .B2(KEYINPUT24), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n665), .B1(new_n481), .B2(new_n482), .ZN(new_n666));
  AOI211_X1 g0466(.A(new_n607), .B(new_n281), .C1(new_n567), .C2(new_n572), .ZN(new_n667));
  INV_X1    g0467(.A(new_n603), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n593), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n606), .A2(new_n607), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n518), .A2(new_n511), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n665), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n666), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n661), .B1(new_n674), .B2(new_n651), .ZN(new_n675));
  OAI21_X1  g0475(.A(KEYINPUT26), .B1(new_n565), .B2(new_n651), .ZN(new_n676));
  OAI221_X1 g0476(.A(new_n554), .B1(G179), .B2(new_n534), .C1(new_n558), .C2(new_n559), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n467), .B1(new_n675), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(KEYINPUT18), .B1(new_n425), .B2(new_n460), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n461), .A2(new_n455), .A3(new_n463), .ZN(new_n681));
  INV_X1    g0481(.A(new_n381), .ZN(new_n682));
  AOI22_X1  g0482(.A1(new_n324), .A2(new_n291), .B1(new_n404), .B2(new_n682), .ZN(new_n683));
  OAI211_X1 g0483(.A(new_n680), .B(new_n681), .C1(new_n683), .C2(new_n447), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n398), .A2(new_n400), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n349), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n679), .A2(new_n686), .ZN(G369));
  INV_X1    g0487(.A(KEYINPUT27), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n310), .A2(new_n688), .A3(new_n207), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(G213), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n688), .B1(new_n310), .B2(new_n207), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  OR2_X1    g0492(.A1(new_n692), .A2(KEYINPUT91), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(KEYINPUT91), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n693), .A2(G343), .A3(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n508), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n521), .A2(new_n671), .A3(new_n695), .A4(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n673), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n698), .B1(new_n699), .B2(new_n696), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n700), .A2(KEYINPUT92), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(KEYINPUT92), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n695), .B1(new_n587), .B2(new_n590), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n704), .B1(new_n608), .B2(new_n597), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n705), .B1(new_n608), .B2(new_n704), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(G330), .ZN(new_n707));
  INV_X1    g0507(.A(new_n519), .ZN(new_n708));
  AOI21_X1  g0508(.A(KEYINPUT89), .B1(new_n518), .B2(new_n511), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n508), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  AOI22_X1  g0511(.A1(new_n521), .A2(new_n697), .B1(new_n711), .B2(new_n696), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n707), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n703), .A2(new_n714), .ZN(G399));
  INV_X1    g0515(.A(new_n210), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(G41), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(KEYINPUT93), .B1(new_n718), .B2(new_n216), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n544), .A2(G116), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n717), .A2(new_n721), .A3(new_n206), .ZN(new_n722));
  MUX2_X1   g0522(.A(new_n719), .B(KEYINPUT93), .S(new_n722), .Z(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT28), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n475), .A2(new_n536), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n725), .A2(new_n668), .A3(KEYINPUT30), .A4(new_n639), .ZN(new_n726));
  AOI21_X1  g0526(.A(G179), .B1(new_n567), .B2(new_n572), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n648), .A2(new_n727), .A3(new_n517), .A4(new_n534), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n475), .A2(new_n536), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n730), .A2(new_n648), .A3(new_n603), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(KEYINPUT30), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT94), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n729), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(KEYINPUT94), .B1(new_n731), .B2(KEYINPUT30), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n695), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n652), .A2(new_n521), .A3(new_n566), .A4(new_n695), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n736), .B1(new_n737), .B2(KEYINPUT31), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n732), .A2(new_n729), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT31), .ZN(new_n740));
  NOR3_X1   g0540(.A1(new_n739), .A2(new_n740), .A3(new_n695), .ZN(new_n741));
  OR2_X1    g0541(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G330), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT95), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n659), .A2(new_n677), .ZN(new_n745));
  OAI211_X1 g0545(.A(new_n647), .B(KEYINPUT26), .C1(new_n649), .C2(new_n650), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n744), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n746), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n748), .A2(KEYINPUT95), .A3(new_n659), .A4(new_n677), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n660), .B1(new_n565), .B2(new_n651), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n747), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n745), .A2(new_n509), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n710), .A2(new_n608), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n641), .A2(new_n651), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT96), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n641), .A2(new_n651), .A3(KEYINPUT96), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n752), .A2(new_n753), .A3(new_n756), .A4(new_n757), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n751), .A2(new_n758), .A3(new_n677), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n759), .A2(KEYINPUT29), .A3(new_n695), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n695), .B1(new_n675), .B2(new_n678), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT29), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n743), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n724), .B1(new_n766), .B2(G1), .ZN(G364));
  INV_X1    g0567(.A(new_n707), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n309), .A2(G20), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n206), .B1(new_n769), .B2(G45), .ZN(new_n770));
  AND2_X1   g0570(.A1(new_n718), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n768), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(G330), .B2(new_n706), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n771), .B(KEYINPUT97), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n213), .B1(G20), .B2(new_n281), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n207), .A2(new_n434), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n779), .A2(new_n377), .A3(G200), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G322), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n377), .A2(new_n385), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n778), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(G326), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n781), .A2(new_n782), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n207), .A2(G190), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR3_X1   g0588(.A1(new_n788), .A2(new_n377), .A3(G200), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n448), .B(new_n786), .C1(G311), .C2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G179), .A2(G200), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT99), .ZN(new_n792));
  OAI21_X1  g0592(.A(G20), .B1(new_n792), .B2(new_n434), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G294), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n792), .A2(new_n788), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G329), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n385), .A2(G179), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n787), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(G283), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  XOR2_X1   g0600(.A(KEYINPUT33), .B(G317), .Z(new_n801));
  NAND2_X1  g0601(.A1(new_n783), .A2(new_n787), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n778), .A2(new_n797), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n800), .B(new_n803), .C1(G303), .C2(new_n805), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n790), .A2(new_n794), .A3(new_n796), .A4(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n795), .A2(G159), .ZN(new_n808));
  XOR2_X1   g0608(.A(new_n808), .B(KEYINPUT32), .Z(new_n809));
  INV_X1    g0609(.A(new_n784), .ZN(new_n810));
  INV_X1    g0610(.A(new_n798), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n810), .A2(G50), .B1(new_n811), .B2(G107), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n812), .B1(new_n329), .B2(new_n781), .ZN(new_n813));
  INV_X1    g0613(.A(new_n789), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n448), .B1(new_n814), .B2(new_n350), .ZN(new_n815));
  AND2_X1   g0615(.A1(new_n540), .A2(new_n542), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n816), .A2(new_n804), .B1(new_n802), .B2(new_n311), .ZN(new_n817));
  NOR3_X1   g0617(.A1(new_n813), .A2(new_n815), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n793), .A2(G97), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n809), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n777), .B1(new_n807), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(G13), .A2(G33), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n823), .A2(G20), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n824), .A2(new_n776), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n419), .A2(new_n421), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n716), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n828), .B1(new_n246), .B2(new_n217), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT98), .ZN(new_n830));
  OR2_X1    g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n829), .A2(new_n830), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n831), .B(new_n832), .C1(new_n246), .C2(new_n243), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n716), .A2(new_n338), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n834), .A2(G355), .B1(new_n579), .B2(new_n716), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n775), .B(new_n821), .C1(new_n825), .C2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n824), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n837), .B1(new_n706), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n773), .A2(new_n839), .ZN(G396));
  INV_X1    g0640(.A(new_n743), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n381), .A2(new_n696), .ZN(new_n842));
  OAI21_X1  g0642(.A(KEYINPUT103), .B1(new_n366), .B2(new_n695), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT103), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n696), .B(new_n844), .C1(new_n380), .C2(new_n352), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n843), .A2(new_n376), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n842), .B1(new_n846), .B2(new_n381), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n761), .B(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n771), .B1(new_n841), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n841), .A2(new_n848), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n847), .A2(new_n823), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n777), .A2(new_n823), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n798), .A2(new_n539), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n810), .A2(G303), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(new_n814), .B2(new_n579), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n854), .B(new_n856), .C1(G294), .C2(new_n780), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n448), .B1(new_n805), .B2(G107), .ZN(new_n858));
  XOR2_X1   g0658(.A(new_n802), .B(KEYINPUT100), .Z(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n860), .A2(G283), .B1(G311), .B2(new_n795), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n857), .A2(new_n819), .A3(new_n858), .A4(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n802), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n780), .A2(G143), .B1(G150), .B2(new_n863), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n789), .A2(G159), .B1(new_n810), .B2(G137), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT34), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI22_X1  g0668(.A1(new_n804), .A2(new_n202), .B1(new_n798), .B2(new_n311), .ZN(new_n869));
  INV_X1    g0669(.A(new_n826), .ZN(new_n870));
  AOI211_X1 g0670(.A(new_n869), .B(new_n870), .C1(G132), .C2(new_n795), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n793), .ZN(new_n873));
  OAI22_X1  g0673(.A1(new_n866), .A2(new_n867), .B1(new_n329), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n862), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n875), .A2(KEYINPUT101), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n776), .B1(new_n875), .B2(KEYINPUT101), .ZN(new_n877));
  OAI221_X1 g0677(.A(new_n774), .B1(G77), .B2(new_n853), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n878), .B(KEYINPUT102), .ZN(new_n879));
  OAI22_X1  g0679(.A1(new_n850), .A2(new_n851), .B1(new_n852), .B2(new_n879), .ZN(G384));
  NAND2_X1  g0680(.A1(new_n613), .A2(new_n618), .ZN(new_n881));
  OAI211_X1 g0681(.A(G116), .B(new_n214), .C1(new_n881), .C2(KEYINPUT35), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(KEYINPUT35), .B2(new_n881), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n883), .B(KEYINPUT36), .ZN(new_n884));
  OR3_X1    g0684(.A1(new_n216), .A2(new_n350), .A3(new_n411), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n202), .A2(G68), .ZN(new_n886));
  AOI211_X1 g0686(.A(new_n206), .B(G13), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n325), .A2(new_n696), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT39), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n424), .A2(new_n293), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n415), .B1(new_n423), .B2(new_n311), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n417), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n406), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n693), .A2(new_n694), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n443), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n894), .A2(new_n460), .ZN(new_n897));
  OAI21_X1  g0697(.A(KEYINPUT37), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n895), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n456), .A2(new_n458), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT37), .B1(new_n425), .B2(new_n442), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n462), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n898), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n894), .A2(new_n895), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n903), .B1(new_n466), .B2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT38), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n903), .B(KEYINPUT38), .C1(new_n466), .C2(new_n905), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n890), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n900), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n681), .A2(new_n680), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n911), .B1(new_n447), .B2(new_n912), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n462), .A2(new_n900), .A3(new_n901), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT37), .ZN(new_n915));
  AND3_X1   g0715(.A1(new_n442), .A2(new_n454), .A3(new_n453), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n425), .A2(new_n460), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n915), .B1(new_n918), .B2(new_n900), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n913), .B1(new_n914), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n907), .ZN(new_n921));
  AND3_X1   g0721(.A1(new_n921), .A2(new_n890), .A3(new_n909), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n889), .B1(new_n910), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n324), .A2(new_n696), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n325), .A2(new_n404), .A3(new_n924), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n403), .A2(new_n306), .A3(new_n323), .A4(new_n307), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n926), .B1(G200), .B2(new_n286), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n324), .B(new_n696), .C1(new_n291), .C2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n695), .B(new_n847), .C1(new_n675), .C2(new_n678), .ZN(new_n930));
  INV_X1    g0730(.A(new_n842), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n908), .A2(new_n909), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n933), .A2(new_n934), .B1(new_n912), .B2(new_n895), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n923), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n760), .A2(new_n467), .A3(new_n763), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n686), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n936), .B(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT40), .ZN(new_n940));
  INV_X1    g0740(.A(new_n447), .ZN(new_n941));
  AOI211_X1 g0741(.A(KEYINPUT78), .B(new_n406), .C1(new_n418), .C2(new_n424), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n457), .B1(new_n453), .B2(new_n454), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(KEYINPUT18), .B1(new_n944), .B2(new_n461), .ZN(new_n945));
  INV_X1    g0745(.A(new_n465), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n941), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n904), .ZN(new_n948));
  AOI21_X1  g0748(.A(KEYINPUT38), .B1(new_n948), .B2(new_n903), .ZN(new_n949));
  INV_X1    g0749(.A(new_n909), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n736), .A2(KEYINPUT31), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n929), .B(new_n847), .C1(new_n738), .C2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n940), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n940), .B1(new_n921), .B2(new_n909), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n738), .A2(new_n952), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n955), .A2(new_n847), .A3(new_n929), .A4(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n956), .A2(new_n467), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n958), .B(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(G330), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n939), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n206), .B2(new_n769), .ZN(new_n963));
  NOR3_X1   g0763(.A1(new_n939), .A2(new_n960), .A3(new_n961), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n888), .B1(new_n963), .B2(new_n964), .ZN(G367));
  OAI211_X1 g0765(.A(new_n756), .B(new_n757), .C1(new_n623), .C2(new_n695), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n651), .A2(new_n695), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT104), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n651), .B1(new_n970), .B2(new_n710), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n695), .ZN(new_n972));
  OAI21_X1  g0772(.A(KEYINPUT42), .B1(new_n970), .B2(new_n698), .ZN(new_n973));
  OR3_X1    g0773(.A1(new_n970), .A2(KEYINPUT42), .A3(new_n698), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n695), .B1(new_n550), .B2(new_n552), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n976), .B1(new_n659), .B2(new_n677), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(new_n677), .B2(new_n976), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n978), .A2(KEYINPUT43), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n978), .A2(KEYINPUT43), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT105), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n975), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n714), .A2(new_n970), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n980), .B1(new_n975), .B2(new_n982), .ZN(new_n987));
  OR3_X1    g0787(.A1(new_n984), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n986), .B1(new_n984), .B2(new_n987), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n717), .B(KEYINPUT41), .Z(new_n990));
  NAND3_X1  g0790(.A1(new_n701), .A2(new_n970), .A3(new_n702), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT44), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n991), .B(new_n992), .ZN(new_n993));
  AND2_X1   g0793(.A1(new_n700), .A2(KEYINPUT92), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n700), .A2(KEYINPUT92), .ZN(new_n995));
  OAI211_X1 g0795(.A(KEYINPUT45), .B(new_n969), .C1(new_n994), .C2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(KEYINPUT45), .B1(new_n703), .B2(new_n969), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n993), .B(new_n714), .C1(new_n997), .C2(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n991), .B(KEYINPUT44), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n998), .A2(new_n997), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n713), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n671), .A2(new_n695), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n712), .A2(KEYINPUT106), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(new_n698), .ZN(new_n1005));
  AOI21_X1  g0805(.A(KEYINPUT106), .B1(new_n712), .B2(new_n1003), .ZN(new_n1006));
  OR2_X1    g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(new_n707), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1008), .A2(new_n765), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n999), .A2(new_n1002), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n990), .B1(new_n1010), .B2(new_n766), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n770), .B(KEYINPUT107), .Z(new_n1012));
  OAI211_X1 g0812(.A(new_n988), .B(new_n989), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n860), .A2(G159), .B1(G137), .B2(new_n795), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n338), .B1(new_n811), .B2(G77), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n789), .A2(G50), .B1(new_n810), .B2(G143), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n780), .A2(G150), .B1(G58), .B2(new_n805), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n873), .A2(new_n311), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n860), .A2(G294), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n795), .A2(G317), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n798), .A2(new_n576), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(G311), .B2(new_n810), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(G303), .A2(new_n780), .B1(new_n789), .B2(G283), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1020), .A2(new_n1021), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n793), .A2(G107), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n805), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT46), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n804), .B2(new_n579), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1026), .A2(new_n870), .A3(new_n1027), .A4(new_n1029), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n1018), .A2(new_n1019), .B1(new_n1025), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT47), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1033), .A2(new_n776), .A3(new_n1034), .ZN(new_n1035));
  AND2_X1   g0835(.A1(new_n827), .A2(new_n235), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n825), .B1(new_n210), .B2(new_n353), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1035), .B(new_n774), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT108), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n838), .B2(new_n978), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1013), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(KEYINPUT109), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT109), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1013), .A2(new_n1043), .A3(new_n1040), .ZN(new_n1044));
  AND2_X1   g0844(.A1(new_n1042), .A2(new_n1044), .ZN(G387));
  INV_X1    g0845(.A(new_n1009), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1008), .A2(new_n765), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1046), .A2(new_n1047), .A3(new_n717), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1008), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n712), .A2(new_n824), .ZN(new_n1050));
  AOI211_X1 g0850(.A(G45), .B(new_n721), .C1(G68), .C2(G77), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n333), .A2(new_n202), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT50), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n828), .B1(new_n1051), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT110), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n1055), .A2(new_n1056), .B1(G45), .B2(new_n232), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n1056), .B2(new_n1055), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n834), .A2(new_n721), .B1(new_n489), .B2(new_n716), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  AND2_X1   g0860(.A1(new_n1060), .A2(new_n825), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n814), .A2(new_n311), .B1(new_n362), .B2(new_n802), .ZN(new_n1062));
  INV_X1    g0862(.A(G159), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n784), .A2(new_n1063), .B1(new_n804), .B2(new_n350), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n1022), .B(new_n870), .C1(G50), .C2(new_n780), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n793), .A2(new_n556), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(KEYINPUT111), .B(G150), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n795), .A2(new_n1068), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .A4(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(G311), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n859), .A2(new_n1071), .B1(new_n782), .B2(new_n784), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT112), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(G317), .A2(new_n780), .B1(new_n789), .B2(G303), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  OR2_X1    g0876(.A1(new_n1076), .A2(KEYINPUT48), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n793), .A2(G283), .B1(G294), .B2(new_n805), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(new_n1076), .B2(KEYINPUT48), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1077), .A2(KEYINPUT49), .A3(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n826), .B1(G116), .B2(new_n811), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n795), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1081), .B(new_n1082), .C1(new_n785), .C2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(KEYINPUT49), .B1(new_n1077), .B2(new_n1080), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1070), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n775), .B(new_n1061), .C1(new_n1086), .C2(new_n776), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n1049), .A2(new_n1012), .B1(new_n1050), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1048), .A2(new_n1088), .ZN(G393));
  NAND2_X1  g0889(.A1(new_n999), .A2(new_n1002), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n1046), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1091), .A2(new_n717), .A3(new_n1010), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n999), .A2(new_n1002), .A3(new_n1012), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n240), .A2(new_n828), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n825), .B1(new_n576), .B2(new_n210), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n774), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n814), .A2(new_n362), .B1(new_n539), .B2(new_n798), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n870), .B(new_n1097), .C1(G68), .C2(new_n805), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n780), .A2(G159), .B1(new_n810), .B2(G150), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1099), .A2(KEYINPUT51), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(G50), .B2(new_n860), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n1099), .A2(KEYINPUT51), .B1(G143), .B2(new_n795), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n793), .A2(G77), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1098), .A2(new_n1101), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n338), .B1(new_n489), .B2(new_n798), .C1(new_n814), .C2(new_n470), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(G303), .B2(new_n860), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n780), .A2(G311), .B1(new_n810), .B2(G317), .ZN(new_n1107));
  XOR2_X1   g0907(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n1108));
  XNOR2_X1  g0908(.A(new_n1107), .B(new_n1108), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1106), .B(new_n1109), .C1(new_n579), .C2(new_n873), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n795), .A2(G322), .B1(G283), .B2(new_n805), .ZN(new_n1111));
  XOR2_X1   g0911(.A(new_n1111), .B(KEYINPUT114), .Z(new_n1112));
  OAI21_X1  g0912(.A(new_n1104), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1096), .B1(new_n1113), .B2(new_n776), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n969), .B2(new_n838), .ZN(new_n1115));
  AND2_X1   g0915(.A1(new_n1093), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1092), .A2(new_n1116), .ZN(G390));
  OAI21_X1  g0917(.A(KEYINPUT39), .B1(new_n949), .B2(new_n950), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n921), .A2(new_n909), .A3(new_n890), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1118), .A2(new_n822), .A3(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n774), .B1(new_n333), .B2(new_n853), .ZN(new_n1121));
  XOR2_X1   g0921(.A(new_n1121), .B(KEYINPUT115), .Z(new_n1122));
  AND2_X1   g0922(.A1(new_n795), .A2(G125), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n780), .A2(G132), .B1(new_n810), .B2(G128), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(KEYINPUT54), .B(G143), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1124), .B1(new_n814), .B2(new_n1125), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n1123), .B(new_n1126), .C1(G137), .C2(new_n860), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n805), .A2(new_n1068), .ZN(new_n1128));
  XOR2_X1   g0928(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n1129));
  OR2_X1    g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n338), .B1(new_n811), .B2(G50), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1130), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(new_n793), .B2(G159), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n859), .A2(new_n489), .B1(new_n1083), .B2(new_n470), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n338), .B1(new_n798), .B2(new_n311), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n781), .A2(new_n579), .B1(new_n814), .B2(new_n576), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n784), .A2(new_n799), .B1(new_n804), .B2(new_n539), .ZN(new_n1138));
  NOR4_X1   g0938(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n1127), .A2(new_n1134), .B1(new_n1139), .B2(new_n1103), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1120), .B(new_n1122), .C1(new_n777), .C2(new_n1140), .ZN(new_n1141));
  OAI211_X1 g0941(.A(G330), .B(new_n847), .C1(new_n738), .C2(new_n952), .ZN(new_n1142));
  AND2_X1   g0942(.A1(new_n925), .A2(new_n928), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n889), .B1(new_n929), .B2(new_n932), .ZN(new_n1145));
  NOR3_X1   g0945(.A1(new_n910), .A2(new_n922), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n846), .A2(new_n381), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n759), .A2(new_n695), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1143), .B1(new_n931), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n921), .A2(new_n909), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n889), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1144), .B1(new_n1146), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n929), .A2(new_n932), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(new_n1151), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1118), .A2(new_n1156), .A3(new_n1119), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n742), .A2(G330), .A3(new_n847), .A4(new_n929), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1157), .B(new_n1158), .C1(new_n1149), .C2(new_n1152), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1154), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1012), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1141), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n686), .B(new_n937), .C1(new_n959), .C2(new_n961), .ZN(new_n1163));
  OAI211_X1 g0963(.A(G330), .B(new_n847), .C1(new_n738), .C2(new_n741), .ZN(new_n1164));
  AND2_X1   g0964(.A1(new_n1164), .A2(new_n1143), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n932), .B1(new_n1165), .B2(new_n1144), .ZN(new_n1166));
  AND2_X1   g0966(.A1(new_n1148), .A2(new_n931), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1158), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1163), .B1(new_n1166), .B2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1170), .A2(new_n1154), .A3(new_n1159), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1170), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n718), .B1(new_n1160), .B2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1162), .B1(new_n1171), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(G378));
  NAND3_X1  g0975(.A1(new_n954), .A2(G330), .A3(new_n957), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n895), .A2(new_n337), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n349), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1179), .B1(new_n685), .B2(new_n1180), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n349), .B(new_n1178), .C1(new_n398), .C2(new_n400), .ZN(new_n1182));
  XOR2_X1   g0982(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1183));
  OR3_X1    g0983(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1183), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  AND3_X1   g0987(.A1(new_n923), .A2(new_n935), .A3(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1187), .B1(new_n923), .B2(new_n935), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1177), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1151), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n912), .A2(new_n895), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n951), .B2(new_n1155), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1186), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n923), .A2(new_n935), .A3(new_n1187), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1194), .A2(new_n1176), .A3(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1190), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(new_n1012), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n771), .B1(G50), .B2(new_n853), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n245), .B1(new_n798), .B2(new_n329), .C1(new_n350), .C2(new_n804), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n826), .B(new_n1200), .C1(G283), .C2(new_n795), .ZN(new_n1201));
  XOR2_X1   g1001(.A(new_n1201), .B(KEYINPUT118), .Z(new_n1202));
  AOI22_X1  g1002(.A1(new_n780), .A2(G107), .B1(new_n810), .B2(G116), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n576), .B2(new_n802), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n1019), .B(new_n1204), .C1(new_n556), .C2(new_n789), .ZN(new_n1205));
  AND2_X1   g1005(.A1(new_n1202), .A2(new_n1205), .ZN(new_n1206));
  OR2_X1    g1006(.A1(new_n1206), .A2(KEYINPUT58), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(KEYINPUT58), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n826), .A2(G33), .ZN(new_n1209));
  AOI21_X1  g1009(.A(G50), .B1(new_n1209), .B2(new_n245), .ZN(new_n1210));
  XOR2_X1   g1010(.A(new_n1210), .B(KEYINPUT117), .Z(new_n1211));
  INV_X1    g1011(.A(new_n1125), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n805), .A2(new_n1212), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT119), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n793), .A2(G150), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n780), .A2(G128), .B1(new_n810), .B2(G125), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n789), .A2(G137), .B1(new_n863), .B2(G132), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .A4(new_n1217), .ZN(new_n1218));
  OR2_X1    g1018(.A1(new_n1218), .A2(KEYINPUT59), .ZN(new_n1219));
  AOI211_X1 g1019(.A(G33), .B(G41), .C1(new_n811), .C2(G159), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(KEYINPUT120), .B(G124), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1220), .B1(new_n1083), .B2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(new_n1218), .B2(KEYINPUT59), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1211), .B1(new_n1219), .B2(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1207), .A2(new_n1208), .A3(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1199), .B1(new_n1225), .B2(new_n776), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1226), .B1(new_n1186), .B2(new_n823), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1198), .A2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1163), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1171), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1197), .A2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(KEYINPUT57), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT57), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1197), .A2(new_n1230), .A3(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1232), .A2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1228), .B1(new_n1235), .B2(new_n717), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(G375));
  OAI21_X1  g1037(.A(new_n774), .B1(G68), .B2(new_n853), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n860), .A2(G116), .B1(G303), .B2(new_n795), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n448), .B1(new_n811), .B2(G77), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n781), .A2(new_n799), .B1(new_n814), .B2(new_n489), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n784), .A2(new_n470), .B1(new_n804), .B2(new_n576), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1239), .A2(new_n1067), .A3(new_n1240), .A4(new_n1243), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n860), .A2(new_n1212), .B1(G128), .B2(new_n795), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n810), .A2(G132), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(G137), .A2(new_n780), .B1(new_n789), .B2(G150), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n804), .A2(new_n1063), .B1(new_n798), .B2(new_n329), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n870), .A2(new_n1248), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1245), .A2(new_n1246), .A3(new_n1247), .A4(new_n1249), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n873), .A2(new_n202), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1244), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1238), .B1(new_n1252), .B2(new_n776), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1253), .B1(new_n929), .B2(new_n823), .ZN(new_n1254));
  AND2_X1   g1054(.A1(new_n1166), .A2(new_n1169), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1254), .B1(new_n1255), .B2(new_n1161), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n990), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1166), .A2(new_n1163), .A3(new_n1169), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1172), .A2(new_n1258), .A3(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1257), .A2(new_n1260), .ZN(G381));
  NAND4_X1  g1061(.A1(new_n1088), .A2(new_n839), .A3(new_n773), .A4(new_n1048), .ZN(new_n1262));
  OR3_X1    g1062(.A1(G390), .A2(G384), .A3(new_n1262), .ZN(new_n1263));
  NOR3_X1   g1063(.A1(G387), .A2(G381), .A3(new_n1263), .ZN(new_n1264));
  XOR2_X1   g1064(.A(new_n1264), .B(KEYINPUT121), .Z(new_n1265));
  NAND2_X1  g1065(.A1(new_n1236), .A2(new_n1174), .ZN(new_n1266));
  OR2_X1    g1066(.A1(new_n1265), .A2(new_n1266), .ZN(G407));
  INV_X1    g1067(.A(G343), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1236), .A2(new_n1268), .A3(new_n1174), .ZN(new_n1269));
  OAI211_X1 g1069(.A(G213), .B(new_n1269), .C1(new_n1265), .C2(new_n1266), .ZN(G409));
  NAND3_X1  g1070(.A1(new_n1013), .A2(new_n1040), .A3(G390), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT125), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1013), .A2(G390), .A3(KEYINPUT125), .A4(new_n1040), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(G390), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1042), .A2(new_n1044), .A3(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(G393), .A2(G396), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(new_n1262), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1275), .A2(new_n1277), .A3(new_n1279), .ZN(new_n1280));
  XOR2_X1   g1080(.A(new_n1279), .B(KEYINPUT124), .Z(new_n1281));
  AOI21_X1  g1081(.A(G390), .B1(new_n1013), .B2(new_n1040), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1271), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1281), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1280), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT61), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(new_n1259), .B(KEYINPUT60), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1288), .A2(new_n717), .A3(new_n1172), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1257), .ZN(new_n1290));
  INV_X1    g1090(.A(G384), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1289), .A2(G384), .A3(new_n1257), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1268), .A2(G213), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(G2897), .ZN(new_n1297));
  XNOR2_X1  g1097(.A(new_n1294), .B(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1228), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1197), .A2(new_n1230), .A3(new_n1258), .ZN(new_n1300));
  AOI21_X1  g1100(.A(G378), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  AND3_X1   g1101(.A1(new_n1197), .A2(new_n1230), .A3(new_n1233), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1233), .B1(new_n1197), .B2(new_n1230), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n717), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1304), .A2(G378), .A3(new_n1299), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT122), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1304), .A2(G378), .A3(KEYINPUT122), .A4(new_n1299), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1301), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1298), .B1(new_n1309), .B2(new_n1296), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1301), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1296), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1294), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  OAI211_X1 g1115(.A(new_n1287), .B(new_n1310), .C1(new_n1315), .C2(KEYINPUT62), .ZN(new_n1316));
  AND2_X1   g1116(.A1(new_n1315), .A2(KEYINPUT62), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1286), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1318));
  XOR2_X1   g1118(.A(KEYINPUT123), .B(KEYINPUT63), .Z(new_n1319));
  AOI21_X1  g1119(.A(new_n1319), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT63), .ZN(new_n1321));
  NOR4_X1   g1121(.A1(new_n1309), .A2(new_n1321), .A3(new_n1296), .A4(new_n1294), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1320), .A2(new_n1322), .ZN(new_n1323));
  AND3_X1   g1123(.A1(new_n1310), .A2(new_n1285), .A3(new_n1287), .ZN(new_n1324));
  AOI21_X1  g1124(.A(KEYINPUT126), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1325));
  AOI21_X1  g1125(.A(KEYINPUT122), .B1(new_n1236), .B2(G378), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1308), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1312), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1328));
  NAND4_X1  g1128(.A1(new_n1328), .A2(KEYINPUT63), .A3(new_n1295), .A4(new_n1314), .ZN(new_n1329));
  NOR3_X1   g1129(.A1(new_n1309), .A2(new_n1296), .A3(new_n1294), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1329), .B1(new_n1330), .B2(new_n1319), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1310), .A2(new_n1285), .A3(new_n1287), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT126), .ZN(new_n1333));
  NOR3_X1   g1133(.A1(new_n1331), .A2(new_n1332), .A3(new_n1333), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1318), .B1(new_n1325), .B2(new_n1334), .ZN(G405));
  XNOR2_X1  g1135(.A(new_n1285), .B(new_n1294), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1311), .B1(G378), .B2(new_n1236), .ZN(new_n1337));
  XNOR2_X1  g1137(.A(new_n1337), .B(KEYINPUT127), .ZN(new_n1338));
  XNOR2_X1  g1138(.A(new_n1336), .B(new_n1338), .ZN(G402));
endmodule


