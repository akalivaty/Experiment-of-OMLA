//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 1 0 1 0 1 0 0 0 1 1 1 0 0 1 1 1 1 1 0 1 1 0 1 0 1 1 0 0 0 0 0 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:02 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(G119), .B(G128), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n190), .B(KEYINPUT72), .ZN(new_n191));
  XOR2_X1   g005(.A(KEYINPUT24), .B(G110), .Z(new_n192));
  INV_X1    g006(.A(KEYINPUT23), .ZN(new_n193));
  INV_X1    g007(.A(G119), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n193), .B1(new_n194), .B2(G128), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(KEYINPUT23), .A3(G119), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n195), .B(new_n197), .C1(G119), .C2(new_n196), .ZN(new_n198));
  OAI22_X1  g012(.A1(new_n191), .A2(new_n192), .B1(G110), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G140), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G125), .ZN(new_n201));
  INV_X1    g015(.A(G125), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G140), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n201), .A2(new_n203), .A3(KEYINPUT16), .ZN(new_n204));
  OR3_X1    g018(.A1(new_n202), .A2(KEYINPUT16), .A3(G140), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(new_n205), .A3(G146), .ZN(new_n206));
  XNOR2_X1  g020(.A(G125), .B(G140), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n199), .A2(new_n206), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n191), .A2(new_n192), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n204), .A2(new_n205), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(new_n208), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(new_n206), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n198), .A2(G110), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n211), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n210), .A2(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n217), .A2(KEYINPUT74), .ZN(new_n218));
  INV_X1    g032(.A(G953), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(G221), .A3(G234), .ZN(new_n220));
  XNOR2_X1  g034(.A(new_n220), .B(KEYINPUT73), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT22), .B(G137), .ZN(new_n222));
  XNOR2_X1  g036(.A(new_n221), .B(new_n222), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n218), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n218), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n217), .A2(KEYINPUT74), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n224), .B1(new_n227), .B2(new_n223), .ZN(new_n228));
  AOI21_X1  g042(.A(KEYINPUT25), .B1(new_n228), .B2(new_n188), .ZN(new_n229));
  INV_X1    g043(.A(new_n223), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n230), .B1(new_n225), .B2(new_n226), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT25), .ZN(new_n232));
  NOR4_X1   g046(.A1(new_n231), .A2(new_n232), .A3(G902), .A4(new_n224), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n189), .B1(new_n229), .B2(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n189), .A2(G902), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n228), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n238));
  OR3_X1    g052(.A1(new_n238), .A2(KEYINPUT2), .A3(G113), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n238), .B1(KEYINPUT2), .B2(G113), .ZN(new_n240));
  AOI22_X1  g054(.A1(new_n239), .A2(new_n240), .B1(KEYINPUT2), .B2(G113), .ZN(new_n241));
  XNOR2_X1  g055(.A(G116), .B(G119), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n194), .A2(G116), .ZN(new_n244));
  INV_X1    g058(.A(G116), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G119), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n247), .B(KEYINPUT68), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n243), .B1(new_n248), .B2(new_n241), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  AND2_X1   g064(.A1(KEYINPUT11), .A2(G134), .ZN(new_n251));
  OR2_X1    g065(.A1(KEYINPUT11), .A2(G134), .ZN(new_n252));
  INV_X1    g066(.A(G137), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  AND2_X1   g069(.A1(KEYINPUT64), .A2(G137), .ZN(new_n256));
  NOR2_X1   g070(.A1(KEYINPUT64), .A2(G137), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(KEYINPUT65), .B1(new_n258), .B2(new_n251), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT64), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(new_n253), .ZN(new_n261));
  NAND2_X1  g075(.A1(KEYINPUT64), .A2(G137), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n261), .A2(new_n251), .A3(KEYINPUT65), .A4(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n255), .B1(new_n259), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G131), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n261), .A2(new_n251), .A3(new_n262), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT65), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n254), .B1(new_n269), .B2(new_n263), .ZN(new_n270));
  INV_X1    g084(.A(G131), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n266), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g087(.A(G143), .B(G146), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n274), .A2(KEYINPUT0), .A3(G128), .ZN(new_n275));
  XNOR2_X1  g089(.A(KEYINPUT0), .B(G128), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n275), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n208), .A2(G143), .ZN(new_n279));
  INV_X1    g093(.A(G143), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G146), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n279), .A2(KEYINPUT1), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n282), .A2(new_n283), .A3(G128), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n279), .B(new_n281), .C1(KEYINPUT1), .C2(new_n196), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n271), .B1(G134), .B2(G137), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n261), .A2(new_n262), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n287), .B1(new_n288), .B2(G134), .ZN(new_n289));
  AND2_X1   g103(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  AOI22_X1  g104(.A1(new_n273), .A2(new_n278), .B1(new_n290), .B2(new_n272), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n250), .B1(new_n291), .B2(KEYINPUT30), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n270), .A2(new_n271), .ZN(new_n293));
  AOI211_X1 g107(.A(G131), .B(new_n254), .C1(new_n269), .C2(new_n263), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n278), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n272), .A2(new_n286), .A3(new_n289), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT30), .ZN(new_n298));
  AOI21_X1  g112(.A(KEYINPUT66), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT66), .ZN(new_n300));
  AOI211_X1 g114(.A(new_n300), .B(KEYINPUT30), .C1(new_n295), .C2(new_n296), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n292), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT31), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n295), .A2(new_n250), .A3(new_n296), .ZN(new_n304));
  NOR2_X1   g118(.A1(G237), .A2(G953), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G210), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n306), .B(KEYINPUT27), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT26), .B(G101), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n307), .B(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n304), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n302), .A2(new_n303), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n309), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT28), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n297), .A2(new_n249), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n314), .B1(new_n315), .B2(new_n304), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n304), .A2(new_n314), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n313), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n312), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT69), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n300), .B1(new_n291), .B2(KEYINPUT30), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n297), .A2(KEYINPUT66), .A3(new_n298), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n310), .B1(new_n324), .B2(new_n292), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n321), .B1(new_n325), .B2(new_n303), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n302), .A2(new_n311), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n327), .A2(KEYINPUT69), .A3(KEYINPUT31), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n320), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  NOR2_X1   g143(.A1(G472), .A2(G902), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  AND3_X1   g146(.A1(new_n295), .A2(new_n250), .A3(new_n296), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n250), .B1(new_n295), .B2(new_n296), .ZN(new_n334));
  OAI21_X1  g148(.A(KEYINPUT28), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n335), .A2(KEYINPUT29), .A3(new_n317), .A4(new_n309), .ZN(new_n336));
  XOR2_X1   g150(.A(new_n336), .B(KEYINPUT71), .Z(new_n337));
  NOR2_X1   g151(.A1(new_n316), .A2(new_n318), .ZN(new_n338));
  AOI21_X1  g152(.A(KEYINPUT29), .B1(new_n338), .B2(new_n309), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n302), .A2(new_n304), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(new_n313), .ZN(new_n341));
  AOI21_X1  g155(.A(G902), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n337), .A2(new_n342), .ZN(new_n343));
  AOI22_X1  g157(.A1(new_n332), .A2(KEYINPUT32), .B1(new_n343), .B2(G472), .ZN(new_n344));
  OAI21_X1  g158(.A(KEYINPUT70), .B1(new_n329), .B2(new_n331), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n312), .A2(new_n319), .ZN(new_n346));
  AOI21_X1  g160(.A(KEYINPUT69), .B1(new_n327), .B2(KEYINPUT31), .ZN(new_n347));
  AOI211_X1 g161(.A(new_n321), .B(new_n303), .C1(new_n302), .C2(new_n311), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n346), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT70), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n349), .A2(new_n350), .A3(new_n330), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT32), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n345), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n237), .B1(new_n344), .B2(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n196), .A2(G143), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n280), .A2(G128), .ZN(new_n356));
  NOR3_X1   g170(.A1(new_n355), .A2(new_n356), .A3(G134), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n356), .B1(KEYINPUT13), .B2(new_n355), .ZN(new_n358));
  NOR3_X1   g172(.A1(new_n355), .A2(KEYINPUT93), .A3(KEYINPUT13), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT93), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n280), .A2(G128), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT13), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n358), .B1(new_n359), .B2(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n357), .B1(new_n364), .B2(G134), .ZN(new_n365));
  INV_X1    g179(.A(G122), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT91), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT91), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G122), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n245), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n245), .A2(G122), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(KEYINPUT92), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT92), .ZN(new_n374));
  XNOR2_X1  g188(.A(KEYINPUT91), .B(G122), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n374), .B(new_n371), .C1(new_n375), .C2(new_n245), .ZN(new_n376));
  AND3_X1   g190(.A1(new_n373), .A2(G107), .A3(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(G107), .B1(new_n373), .B2(new_n376), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n365), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n373), .A2(new_n376), .ZN(new_n380));
  INV_X1    g194(.A(G107), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OR3_X1    g196(.A1(new_n371), .A2(KEYINPUT94), .A3(KEYINPUT14), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n367), .A2(new_n369), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G116), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n371), .A2(KEYINPUT14), .ZN(new_n386));
  OAI21_X1  g200(.A(KEYINPUT94), .B1(new_n371), .B2(KEYINPUT14), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n383), .A2(new_n385), .A3(new_n386), .A4(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(G107), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n355), .A2(new_n356), .ZN(new_n390));
  XOR2_X1   g204(.A(new_n390), .B(G134), .Z(new_n391));
  NAND3_X1  g205(.A1(new_n382), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n379), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(KEYINPUT9), .B(G234), .ZN(new_n394));
  NOR3_X1   g208(.A1(new_n394), .A2(new_n187), .A3(G953), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n379), .A2(new_n392), .A3(new_n395), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n188), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n400), .A2(KEYINPUT95), .ZN(new_n401));
  INV_X1    g215(.A(G478), .ZN(new_n402));
  OR2_X1    g216(.A1(new_n402), .A2(KEYINPUT15), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n401), .B(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(G237), .ZN(new_n405));
  AND4_X1   g219(.A1(G143), .A2(new_n405), .A3(new_n219), .A4(G214), .ZN(new_n406));
  AOI21_X1  g220(.A(G143), .B1(new_n305), .B2(G214), .ZN(new_n407));
  OAI211_X1 g221(.A(KEYINPUT17), .B(G131), .C1(new_n406), .C2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n213), .A2(new_n206), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT88), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT88), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n213), .A2(new_n408), .A3(new_n411), .A4(new_n206), .ZN(new_n412));
  NOR3_X1   g226(.A1(new_n406), .A2(new_n407), .A3(G131), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n405), .A2(new_n219), .A3(G214), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n280), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n305), .A2(G143), .A3(G214), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n271), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n413), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT17), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n410), .A2(new_n412), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT90), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n201), .A2(new_n203), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(G146), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n209), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT86), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT86), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n424), .A2(new_n209), .A3(new_n427), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n415), .A2(KEYINPUT18), .A3(G131), .A4(new_n416), .ZN(new_n429));
  NAND2_X1  g243(.A1(KEYINPUT18), .A2(G131), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n430), .B1(new_n406), .B2(new_n407), .ZN(new_n431));
  AOI22_X1  g245(.A1(new_n426), .A2(new_n428), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  AND3_X1   g247(.A1(new_n421), .A2(new_n422), .A3(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n422), .B1(new_n421), .B2(new_n433), .ZN(new_n436));
  XNOR2_X1  g250(.A(G113), .B(G122), .ZN(new_n437));
  INV_X1    g251(.A(G104), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n437), .B(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n421), .A2(new_n433), .ZN(new_n441));
  INV_X1    g255(.A(new_n439), .ZN(new_n442));
  OAI21_X1  g256(.A(KEYINPUT89), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AOI22_X1  g257(.A1(KEYINPUT88), .A2(new_n409), .B1(new_n418), .B2(new_n419), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n432), .B1(new_n444), .B2(new_n412), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT89), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n445), .A2(new_n446), .A3(new_n439), .ZN(new_n447));
  AOI22_X1  g261(.A1(new_n435), .A2(new_n440), .B1(new_n443), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(G475), .B1(new_n448), .B2(G902), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT87), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n207), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n451), .B(KEYINPUT19), .ZN(new_n452));
  OAI221_X1 g266(.A(new_n206), .B1(new_n417), .B2(new_n413), .C1(new_n452), .C2(G146), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n439), .B1(new_n453), .B2(new_n433), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n454), .B1(new_n443), .B2(new_n447), .ZN(new_n455));
  NOR2_X1   g269(.A1(G475), .A2(G902), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  NOR3_X1   g271(.A1(new_n455), .A2(KEYINPUT20), .A3(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT20), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n446), .B1(new_n445), .B2(new_n439), .ZN(new_n460));
  AND4_X1   g274(.A1(new_n446), .A2(new_n421), .A3(new_n439), .A4(new_n433), .ZN(new_n461));
  AND2_X1   g275(.A1(new_n453), .A2(new_n433), .ZN(new_n462));
  OAI22_X1  g276(.A1(new_n460), .A2(new_n461), .B1(new_n439), .B2(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n459), .B1(new_n463), .B2(new_n456), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n449), .B1(new_n458), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(G234), .A2(G237), .ZN(new_n466));
  AND3_X1   g280(.A1(new_n466), .A2(G952), .A3(new_n219), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n466), .A2(G902), .A3(G953), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n468), .B(KEYINPUT96), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT21), .B(G898), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n467), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR3_X1   g285(.A1(new_n404), .A2(new_n465), .A3(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(G221), .B1(new_n394), .B2(G902), .ZN(new_n473));
  INV_X1    g287(.A(G469), .ZN(new_n474));
  XNOR2_X1  g288(.A(G110), .B(G140), .ZN(new_n475));
  INV_X1    g289(.A(G227), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n476), .A2(G953), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n475), .B(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(KEYINPUT3), .B1(new_n438), .B2(G107), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT3), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n480), .A2(new_n381), .A3(G104), .ZN(new_n481));
  INV_X1    g295(.A(G101), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n438), .A2(G107), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n479), .A2(new_n481), .A3(new_n482), .A4(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n438), .A2(G107), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n381), .A2(G104), .ZN(new_n486));
  OAI21_X1  g300(.A(G101), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n286), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n284), .A2(new_n285), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n488), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n273), .B(new_n493), .C1(KEYINPUT77), .C2(KEYINPUT12), .ZN(new_n494));
  AND2_X1   g308(.A1(new_n273), .A2(new_n493), .ZN(new_n495));
  XOR2_X1   g309(.A(KEYINPUT77), .B(KEYINPUT12), .Z(new_n496));
  OAI21_X1  g310(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  OR3_X1    g312(.A1(new_n293), .A2(new_n294), .A3(KEYINPUT76), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n273), .A2(KEYINPUT76), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT10), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n490), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(G101), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n505), .A2(KEYINPUT4), .A3(new_n484), .ZN(new_n506));
  XNOR2_X1  g320(.A(KEYINPUT75), .B(KEYINPUT4), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n504), .A2(G101), .A3(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n278), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n286), .A2(new_n489), .A3(KEYINPUT10), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n503), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n501), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n478), .B1(new_n498), .B2(new_n512), .ZN(new_n513));
  AND2_X1   g327(.A1(new_n503), .A2(new_n510), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n514), .A2(new_n499), .A3(new_n509), .A4(new_n500), .ZN(new_n515));
  INV_X1    g329(.A(new_n478), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n511), .A2(KEYINPUT78), .A3(new_n273), .ZN(new_n517));
  AOI21_X1  g331(.A(KEYINPUT78), .B1(new_n511), .B2(new_n273), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n515), .B(new_n516), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n513), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(KEYINPUT79), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT79), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n513), .A2(new_n519), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n474), .B1(new_n524), .B2(new_n188), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n515), .B1(new_n517), .B2(new_n518), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n478), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n497), .A2(new_n515), .A3(new_n516), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  XOR2_X1   g343(.A(KEYINPUT80), .B(G469), .Z(new_n530));
  NAND3_X1  g344(.A1(new_n529), .A2(new_n188), .A3(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n473), .B1(new_n525), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(G210), .B1(G237), .B2(G902), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT5), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n536), .A2(new_n194), .A3(G116), .ZN(new_n537));
  AND2_X1   g351(.A1(new_n537), .A2(G113), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n242), .B(KEYINPUT68), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n538), .B1(new_n539), .B2(new_n536), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(KEYINPUT81), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT81), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n542), .B(new_n538), .C1(new_n539), .C2(new_n536), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n541), .A2(new_n543), .A3(new_n243), .A4(new_n488), .ZN(new_n544));
  XNOR2_X1  g358(.A(G110), .B(G122), .ZN(new_n545));
  XOR2_X1   g359(.A(new_n545), .B(KEYINPUT8), .Z(new_n546));
  OAI21_X1  g360(.A(new_n538), .B1(new_n536), .B2(new_n247), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n243), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n546), .B1(new_n548), .B2(new_n489), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n544), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT83), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n544), .A2(KEYINPUT83), .A3(new_n549), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n286), .A2(new_n202), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n555), .B1(new_n202), .B2(new_n277), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n219), .A2(G224), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT7), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n556), .B(new_n558), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n541), .A2(new_n543), .A3(new_n243), .A4(new_n489), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n249), .A2(new_n506), .A3(new_n508), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n560), .A2(new_n545), .A3(new_n561), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(G902), .B1(new_n554), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n560), .A2(new_n561), .ZN(new_n565));
  INV_X1    g379(.A(new_n545), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n567), .A2(KEYINPUT6), .A3(new_n562), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n557), .B(KEYINPUT82), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n556), .B(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT6), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n565), .A2(new_n571), .A3(new_n566), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n568), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n564), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT85), .ZN(new_n575));
  OAI211_X1 g389(.A(KEYINPUT84), .B(new_n535), .C1(new_n574), .C2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n535), .A2(KEYINPUT84), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n564), .A2(new_n573), .A3(KEYINPUT85), .A4(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n564), .A2(new_n573), .A3(new_n534), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n575), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n576), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(G214), .B1(G237), .B2(G902), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n533), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n354), .A2(new_n472), .A3(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(KEYINPUT97), .B(G101), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n585), .B(new_n586), .ZN(G3));
  OAI21_X1  g401(.A(G472), .B1(new_n329), .B2(G902), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n345), .A2(new_n588), .A3(new_n351), .ZN(new_n589));
  NOR3_X1   g403(.A1(new_n589), .A2(new_n533), .A3(new_n237), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n574), .A2(KEYINPUT98), .A3(new_n535), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n579), .ZN(new_n592));
  AOI21_X1  g406(.A(KEYINPUT98), .B1(new_n574), .B2(new_n535), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n582), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(KEYINPUT20), .B1(new_n455), .B2(new_n457), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n463), .A2(new_n459), .A3(new_n456), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n460), .A2(new_n461), .ZN(new_n597));
  NOR3_X1   g411(.A1(new_n434), .A2(new_n436), .A3(new_n439), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n188), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g413(.A1(new_n595), .A2(new_n596), .B1(new_n599), .B2(G475), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n402), .A2(G902), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT33), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(KEYINPUT99), .ZN(new_n604));
  OR2_X1    g418(.A1(new_n603), .A2(KEYINPUT99), .ZN(new_n605));
  AND3_X1   g419(.A1(new_n379), .A2(new_n392), .A3(new_n395), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n395), .B1(new_n379), .B2(new_n392), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n604), .B(new_n605), .C1(new_n606), .C2(new_n607), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n397), .A2(KEYINPUT99), .A3(new_n603), .A4(new_n398), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n602), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(KEYINPUT100), .B(G478), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n612), .B1(new_n399), .B2(new_n188), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  NOR4_X1   g428(.A1(new_n594), .A2(new_n471), .A3(new_n600), .A4(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n590), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(KEYINPUT101), .ZN(new_n617));
  XNOR2_X1  g431(.A(KEYINPUT34), .B(G104), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G6));
  INV_X1    g433(.A(KEYINPUT102), .ZN(new_n620));
  OAI21_X1  g434(.A(KEYINPUT103), .B1(new_n458), .B2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT103), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n596), .A2(KEYINPUT102), .A3(new_n622), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n621), .A2(new_n464), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n464), .B1(new_n621), .B2(new_n623), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n449), .B(new_n404), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n626), .A2(new_n594), .A3(new_n471), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n590), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT35), .B(G107), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G9));
  INV_X1    g444(.A(new_n589), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n230), .A2(KEYINPUT36), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n217), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n235), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n234), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n584), .A2(new_n472), .A3(new_n631), .A4(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT37), .B(G110), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G12));
  OAI211_X1 g452(.A(new_n473), .B(new_n635), .C1(new_n525), .C2(new_n532), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n639), .B1(new_n344), .B2(new_n353), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT104), .B(G900), .Z(new_n641));
  NAND2_X1  g455(.A1(new_n469), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n467), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n626), .A2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n594), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n640), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G128), .ZN(G30));
  INV_X1    g463(.A(new_n533), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT40), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n644), .B(KEYINPUT39), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n404), .A2(new_n465), .ZN(new_n654));
  INV_X1    g468(.A(new_n582), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AND2_X1   g470(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n652), .ZN(new_n658));
  OAI21_X1  g472(.A(KEYINPUT40), .B1(new_n533), .B2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n581), .B(KEYINPUT38), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n332), .A2(KEYINPUT32), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n340), .A2(new_n309), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n315), .A2(new_n304), .ZN(new_n664));
  OAI211_X1 g478(.A(new_n663), .B(new_n188), .C1(new_n664), .C2(new_n309), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(G472), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n353), .A2(new_n662), .A3(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n635), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n657), .A2(new_n661), .A3(KEYINPUT105), .A4(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT105), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n653), .A2(new_n659), .A3(new_n660), .A4(new_n656), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n672), .B1(new_n673), .B2(new_n669), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(new_n280), .ZN(G45));
  NOR2_X1   g490(.A1(new_n600), .A2(new_n614), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n644), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n640), .A2(new_n647), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G146), .ZN(G48));
  NAND2_X1  g495(.A1(new_n344), .A2(new_n353), .ZN(new_n682));
  INV_X1    g496(.A(new_n237), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n529), .A2(new_n188), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(G469), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n686), .A2(new_n473), .A3(new_n531), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(new_n615), .ZN(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT41), .B(G113), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G15));
  NAND2_X1  g505(.A1(new_n688), .A2(new_n627), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G116), .ZN(G18));
  NAND2_X1  g507(.A1(new_n472), .A2(new_n635), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n694), .A2(new_n594), .A3(new_n687), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n682), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT106), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G119), .ZN(G21));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n594), .A2(new_n687), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n654), .A2(new_n471), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n327), .A2(KEYINPUT31), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n331), .B1(new_n346), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n349), .A2(new_n188), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n704), .B1(new_n705), .B2(G472), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n683), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n699), .B1(new_n702), .B2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n707), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n709), .A2(KEYINPUT107), .A3(new_n700), .A4(new_n701), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(KEYINPUT108), .B(G122), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G24));
  AND2_X1   g527(.A1(new_n706), .A2(new_n635), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n714), .A2(new_n679), .A3(new_n700), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G125), .ZN(G27));
  NAND4_X1  g530(.A1(new_n576), .A2(new_n582), .A3(new_n578), .A4(new_n580), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n473), .ZN(new_n719));
  INV_X1    g533(.A(new_n520), .ZN(new_n720));
  OAI21_X1  g534(.A(G469), .B1(new_n720), .B2(G902), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n719), .B1(new_n721), .B2(new_n531), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  NOR4_X1   g537(.A1(new_n684), .A2(KEYINPUT42), .A3(new_n678), .A4(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n723), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n343), .A2(G472), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n352), .B1(new_n329), .B2(new_n331), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n662), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n728), .A2(KEYINPUT109), .A3(new_n683), .ZN(new_n729));
  AOI21_X1  g543(.A(KEYINPUT109), .B1(new_n728), .B2(new_n683), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n679), .B(new_n725), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n724), .B1(new_n731), .B2(KEYINPUT42), .ZN(new_n732));
  XOR2_X1   g546(.A(KEYINPUT110), .B(G131), .Z(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(G33));
  NAND3_X1  g548(.A1(new_n354), .A2(new_n725), .A3(new_n646), .ZN(new_n735));
  XNOR2_X1  g549(.A(KEYINPUT111), .B(G134), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G36));
  INV_X1    g551(.A(KEYINPUT43), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n608), .A2(new_n609), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n601), .ZN(new_n740));
  INV_X1    g554(.A(new_n613), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT112), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  OAI21_X1  g557(.A(KEYINPUT112), .B1(new_n610), .B2(new_n613), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n738), .B1(new_n745), .B2(new_n465), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT113), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n738), .B1(new_n740), .B2(new_n741), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n595), .A2(new_n596), .ZN(new_n749));
  AND4_X1   g563(.A1(new_n747), .A2(new_n748), .A3(new_n749), .A4(new_n449), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n747), .B1(new_n600), .B2(new_n748), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n746), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n589), .A2(new_n752), .A3(KEYINPUT44), .A4(new_n635), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n718), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(KEYINPUT114), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT114), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n753), .A2(new_n756), .A3(new_n718), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n589), .A2(new_n752), .A3(new_n635), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT44), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n755), .A2(new_n757), .A3(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT115), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n474), .A2(new_n188), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT45), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n524), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n474), .B1(new_n720), .B2(KEYINPUT45), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n764), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n768), .A2(KEYINPUT46), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n531), .B1(new_n768), .B2(KEYINPUT46), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(new_n473), .A3(new_n652), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n755), .A2(KEYINPUT115), .A3(new_n757), .A4(new_n760), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n763), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  XOR2_X1   g589(.A(KEYINPUT116), .B(G137), .Z(new_n776));
  XNOR2_X1  g590(.A(new_n775), .B(new_n776), .ZN(G39));
  OAI21_X1  g591(.A(new_n473), .B1(new_n769), .B2(new_n770), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT47), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OAI211_X1 g594(.A(KEYINPUT47), .B(new_n473), .C1(new_n769), .C2(new_n770), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR4_X1   g596(.A1(new_n682), .A2(new_n683), .A3(new_n678), .A4(new_n717), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G140), .ZN(G42));
  INV_X1    g599(.A(new_n614), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n683), .A2(new_n582), .A3(new_n473), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n686), .A2(new_n531), .ZN(new_n788));
  AOI211_X1 g602(.A(new_n465), .B(new_n787), .C1(KEYINPUT49), .C2(new_n788), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n789), .B1(KEYINPUT49), .B2(new_n788), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n790), .A2(new_n667), .A3(new_n660), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT117), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n706), .A2(new_n679), .A3(new_n635), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n793), .A2(new_n594), .A3(new_n687), .ZN(new_n794));
  AOI211_X1 g608(.A(new_n594), .B(new_n639), .C1(new_n353), .C2(new_n344), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n794), .B1(new_n795), .B2(new_n646), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT119), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n594), .A2(new_n654), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n722), .A2(new_n644), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n667), .A2(new_n798), .A3(new_n668), .A4(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n796), .A2(new_n797), .A3(new_n680), .A4(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n648), .A2(new_n680), .A3(new_n715), .A4(new_n800), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(KEYINPUT119), .ZN(new_n803));
  AOI21_X1  g617(.A(KEYINPUT52), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n804), .B1(KEYINPUT52), .B2(new_n802), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT120), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n696), .A2(KEYINPUT106), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT106), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n808), .B1(new_n695), .B2(new_n682), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n711), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n688), .B1(new_n615), .B2(new_n627), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n806), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n697), .A2(new_n811), .A3(KEYINPUT120), .A4(new_n711), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n731), .A2(KEYINPUT42), .ZN(new_n816));
  INV_X1    g630(.A(new_n724), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n793), .A2(new_n723), .ZN(new_n818));
  OR2_X1    g632(.A1(new_n624), .A2(new_n625), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(new_n449), .ZN(new_n820));
  NOR4_X1   g634(.A1(new_n820), .A2(new_n404), .A3(new_n645), .A4(new_n717), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n818), .B1(new_n821), .B2(new_n640), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n816), .A2(new_n817), .A3(new_n735), .A4(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n465), .A2(new_n614), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n824), .B1(new_n465), .B2(new_n404), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n583), .A2(new_n471), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n590), .A2(new_n826), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n585), .A2(new_n827), .A3(new_n636), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(KEYINPUT53), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n823), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n805), .A2(new_n815), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n801), .A2(new_n803), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT52), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n697), .A2(new_n828), .A3(new_n711), .A4(new_n811), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n823), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n801), .A2(new_n803), .A3(KEYINPUT52), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n834), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT54), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n831), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n838), .A2(new_n839), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT118), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n844), .B1(new_n823), .B2(new_n835), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n836), .A2(KEYINPUT118), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n805), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n843), .B1(new_n847), .B2(new_n839), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n842), .B1(new_n848), .B2(new_n841), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n752), .A2(new_n467), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n709), .A2(new_n850), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n660), .A2(new_n582), .A3(new_n687), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XOR2_X1   g667(.A(new_n853), .B(KEYINPUT50), .Z(new_n854));
  NOR2_X1   g668(.A1(new_n717), .A2(new_n687), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n850), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n855), .A2(new_n683), .A3(new_n467), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n857), .A2(new_n667), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n465), .A2(new_n786), .ZN(new_n859));
  AOI22_X1  g673(.A1(new_n856), .A2(new_n714), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n788), .A2(new_n473), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n718), .B(new_n851), .C1(new_n782), .C2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n854), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT51), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n863), .A2(new_n864), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n851), .A2(new_n700), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n858), .A2(new_n677), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n867), .A2(new_n868), .A3(G952), .A4(new_n219), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n856), .B1(new_n729), .B2(new_n730), .ZN(new_n870));
  OR2_X1    g684(.A1(new_n870), .A2(KEYINPUT48), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(KEYINPUT48), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n869), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n865), .A2(new_n866), .A3(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n849), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(G952), .A2(G953), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n792), .B1(new_n875), .B2(new_n876), .ZN(G75));
  NOR2_X1   g691(.A1(new_n219), .A2(G952), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n804), .A2(new_n835), .A3(new_n823), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT53), .B1(new_n879), .B2(new_n837), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n802), .A2(KEYINPUT52), .ZN(new_n881));
  AND4_X1   g695(.A1(new_n834), .A2(new_n815), .A3(new_n830), .A4(new_n881), .ZN(new_n882));
  OAI211_X1 g696(.A(G210), .B(G902), .C1(new_n880), .C2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT56), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n568), .A2(new_n572), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n886), .B(new_n570), .Z(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT55), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n878), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(new_n888), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n883), .A2(KEYINPUT121), .A3(new_n884), .A4(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n883), .A2(new_n884), .A3(new_n890), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT121), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n889), .A2(new_n891), .A3(new_n894), .ZN(G51));
  XNOR2_X1  g709(.A(new_n764), .B(KEYINPUT57), .ZN(new_n896));
  INV_X1    g710(.A(new_n842), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n841), .B1(new_n831), .B2(new_n840), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(new_n529), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n188), .B1(new_n831), .B2(new_n840), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n901), .A2(new_n766), .A3(new_n767), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n878), .B1(new_n900), .B2(new_n902), .ZN(G54));
  NAND2_X1  g717(.A1(KEYINPUT58), .A2(G475), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT122), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n901), .A2(new_n463), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n463), .B1(new_n901), .B2(new_n905), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n906), .A2(new_n907), .A3(new_n878), .ZN(G60));
  NAND2_X1  g722(.A1(G478), .A2(G902), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n909), .B(KEYINPUT59), .Z(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n739), .B1(new_n849), .B2(new_n911), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n739), .B(new_n911), .C1(new_n897), .C2(new_n898), .ZN(new_n913));
  INV_X1    g727(.A(new_n878), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n912), .A2(new_n915), .ZN(G63));
  INV_X1    g730(.A(KEYINPUT61), .ZN(new_n917));
  NAND2_X1  g731(.A1(G217), .A2(G902), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT60), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n919), .B1(new_n831), .B2(new_n840), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n633), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n914), .B1(new_n920), .B2(new_n228), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n917), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OR2_X1    g738(.A1(new_n920), .A2(new_n228), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n925), .A2(KEYINPUT61), .A3(new_n914), .A4(new_n921), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n924), .A2(new_n926), .ZN(G66));
  INV_X1    g741(.A(G224), .ZN(new_n928));
  OAI21_X1  g742(.A(G953), .B1(new_n470), .B2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n835), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n929), .B1(new_n930), .B2(G953), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n886), .B1(G898), .B2(new_n219), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n931), .B(new_n932), .ZN(G69));
  OAI21_X1  g747(.A(new_n324), .B1(new_n298), .B2(new_n297), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(new_n452), .Z(new_n935));
  INV_X1    g749(.A(KEYINPUT123), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n648), .A2(new_n680), .A3(new_n715), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n937), .A2(new_n671), .A3(new_n674), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(KEYINPUT62), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT62), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n937), .A2(new_n671), .A3(new_n674), .A4(new_n940), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n533), .A2(new_n658), .A3(new_n825), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n354), .A2(new_n942), .A3(new_n718), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n939), .A2(new_n784), .A3(new_n941), .A4(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(new_n775), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n936), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n784), .A2(new_n943), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n947), .B1(KEYINPUT62), .B2(new_n938), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n948), .A2(KEYINPUT123), .A3(new_n775), .A4(new_n941), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n946), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n935), .B1(new_n950), .B2(G953), .ZN(new_n951));
  INV_X1    g765(.A(new_n935), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n219), .A2(G900), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n732), .A2(new_n735), .ZN(new_n954));
  INV_X1    g768(.A(new_n784), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n729), .A2(new_n730), .ZN(new_n956));
  INV_X1    g770(.A(new_n798), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n772), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n954), .A2(new_n955), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(KEYINPUT125), .B1(new_n775), .B2(new_n937), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n774), .A2(new_n773), .ZN(new_n961));
  AOI22_X1  g775(.A1(new_n754), .A2(KEYINPUT114), .B1(new_n759), .B2(new_n758), .ZN(new_n962));
  AOI21_X1  g776(.A(KEYINPUT115), .B1(new_n962), .B2(new_n757), .ZN(new_n963));
  OAI211_X1 g777(.A(KEYINPUT125), .B(new_n937), .C1(new_n961), .C2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n959), .B1(new_n960), .B2(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n953), .B1(new_n966), .B2(new_n219), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT126), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n952), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n953), .ZN(new_n970));
  INV_X1    g784(.A(new_n954), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n955), .A2(new_n958), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n937), .B1(new_n961), .B2(new_n963), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT125), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n973), .B1(new_n976), .B2(new_n964), .ZN(new_n977));
  OAI211_X1 g791(.A(new_n968), .B(new_n970), .C1(new_n977), .C2(G953), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n951), .B1(new_n969), .B2(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n953), .B1(new_n476), .B2(G953), .ZN(new_n981));
  XNOR2_X1  g795(.A(KEYINPUT124), .B(KEYINPUT127), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n981), .B(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n980), .A2(new_n984), .ZN(new_n985));
  OAI211_X1 g799(.A(new_n951), .B(new_n983), .C1(new_n969), .C2(new_n979), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(G72));
  NAND2_X1  g801(.A1(new_n950), .A2(new_n930), .ZN(new_n988));
  NAND2_X1  g802(.A1(G472), .A2(G902), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT63), .Z(new_n990));
  AOI21_X1  g804(.A(new_n663), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n977), .A2(new_n930), .ZN(new_n992));
  AOI211_X1 g806(.A(new_n309), .B(new_n340), .C1(new_n992), .C2(new_n990), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n341), .A2(new_n327), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(new_n990), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n914), .B1(new_n848), .B2(new_n995), .ZN(new_n996));
  NOR3_X1   g810(.A1(new_n991), .A2(new_n993), .A3(new_n996), .ZN(G57));
endmodule


