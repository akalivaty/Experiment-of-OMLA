

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U546 ( .A(KEYINPUT65), .B(G2104), .Z(n517) );
  XNOR2_X1 U547 ( .A(n688), .B(KEYINPUT104), .ZN(n690) );
  NOR2_X2 U548 ( .A1(n517), .A2(n518), .ZN(n702) );
  XNOR2_X1 U549 ( .A(n617), .B(KEYINPUT26), .ZN(n618) );
  INV_X1 U550 ( .A(KEYINPUT30), .ZN(n653) );
  XNOR2_X1 U551 ( .A(n653), .B(KEYINPUT103), .ZN(n654) );
  XNOR2_X1 U552 ( .A(n655), .B(n654), .ZN(n656) );
  INV_X1 U553 ( .A(KEYINPUT29), .ZN(n644) );
  XNOR2_X1 U554 ( .A(n645), .B(n644), .ZN(n650) );
  NAND2_X1 U555 ( .A1(n669), .A2(G8), .ZN(n670) );
  INV_X1 U556 ( .A(n855), .ZN(n689) );
  AND2_X1 U557 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U558 ( .A1(G651), .A2(n583), .ZN(n800) );
  AND2_X1 U559 ( .A1(G2105), .A2(G2104), .ZN(n991) );
  NAND2_X1 U560 ( .A1(n991), .A2(G114), .ZN(n513) );
  XNOR2_X1 U561 ( .A(n513), .B(KEYINPUT92), .ZN(n516) );
  NOR2_X1 U562 ( .A1(G2105), .A2(G2104), .ZN(n514) );
  XOR2_X1 U563 ( .A(KEYINPUT17), .B(n514), .Z(n530) );
  NAND2_X1 U564 ( .A1(G138), .A2(n995), .ZN(n515) );
  NAND2_X1 U565 ( .A1(n516), .A2(n515), .ZN(n523) );
  INV_X1 U566 ( .A(G2105), .ZN(n518) );
  NAND2_X1 U567 ( .A1(G126), .A2(n702), .ZN(n521) );
  NAND2_X1 U568 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U569 ( .A(KEYINPUT67), .B(n519), .ZN(n699) );
  NAND2_X1 U570 ( .A1(G102), .A2(n699), .ZN(n520) );
  NAND2_X1 U571 ( .A1(n521), .A2(n520), .ZN(n522) );
  NOR2_X1 U572 ( .A1(n523), .A2(n522), .ZN(G164) );
  NAND2_X1 U573 ( .A1(G125), .A2(n702), .ZN(n524) );
  XNOR2_X1 U574 ( .A(n524), .B(KEYINPUT66), .ZN(n528) );
  NAND2_X1 U575 ( .A1(G101), .A2(n699), .ZN(n526) );
  INV_X1 U576 ( .A(KEYINPUT23), .ZN(n525) );
  XNOR2_X1 U577 ( .A(n526), .B(n525), .ZN(n527) );
  NAND2_X1 U578 ( .A1(n528), .A2(n527), .ZN(n534) );
  NAND2_X1 U579 ( .A1(n991), .A2(G113), .ZN(n529) );
  XNOR2_X1 U580 ( .A(n529), .B(KEYINPUT68), .ZN(n532) );
  BUF_X1 U581 ( .A(n530), .Z(n995) );
  NAND2_X1 U582 ( .A1(G137), .A2(n995), .ZN(n531) );
  NAND2_X1 U583 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X2 U584 ( .A1(n534), .A2(n533), .ZN(G160) );
  NOR2_X1 U585 ( .A1(G651), .A2(G543), .ZN(n792) );
  NAND2_X1 U586 ( .A1(G86), .A2(n792), .ZN(n537) );
  INV_X1 U587 ( .A(G651), .ZN(n539) );
  NOR2_X1 U588 ( .A1(G543), .A2(n539), .ZN(n535) );
  XOR2_X1 U589 ( .A(KEYINPUT1), .B(n535), .Z(n793) );
  NAND2_X1 U590 ( .A1(G61), .A2(n793), .ZN(n536) );
  NAND2_X1 U591 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U592 ( .A(KEYINPUT82), .B(n538), .ZN(n542) );
  XOR2_X1 U593 ( .A(G543), .B(KEYINPUT0), .Z(n583) );
  NOR2_X1 U594 ( .A1(n583), .A2(n539), .ZN(n796) );
  NAND2_X1 U595 ( .A1(n796), .A2(G73), .ZN(n540) );
  XOR2_X1 U596 ( .A(KEYINPUT2), .B(n540), .Z(n541) );
  NOR2_X1 U597 ( .A1(n542), .A2(n541), .ZN(n544) );
  NAND2_X1 U598 ( .A1(n800), .A2(G48), .ZN(n543) );
  NAND2_X1 U599 ( .A1(n544), .A2(n543), .ZN(G305) );
  NAND2_X1 U600 ( .A1(G65), .A2(n793), .ZN(n545) );
  XOR2_X1 U601 ( .A(KEYINPUT72), .B(n545), .Z(n550) );
  NAND2_X1 U602 ( .A1(G91), .A2(n792), .ZN(n547) );
  NAND2_X1 U603 ( .A1(G78), .A2(n796), .ZN(n546) );
  NAND2_X1 U604 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U605 ( .A(KEYINPUT71), .B(n548), .Z(n549) );
  NOR2_X1 U606 ( .A1(n550), .A2(n549), .ZN(n552) );
  NAND2_X1 U607 ( .A1(n800), .A2(G53), .ZN(n551) );
  NAND2_X1 U608 ( .A1(n552), .A2(n551), .ZN(G299) );
  NAND2_X1 U609 ( .A1(G90), .A2(n792), .ZN(n554) );
  NAND2_X1 U610 ( .A1(G77), .A2(n796), .ZN(n553) );
  NAND2_X1 U611 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U612 ( .A(n555), .B(KEYINPUT9), .ZN(n557) );
  NAND2_X1 U613 ( .A1(G64), .A2(n793), .ZN(n556) );
  NAND2_X1 U614 ( .A1(n557), .A2(n556), .ZN(n560) );
  NAND2_X1 U615 ( .A1(G52), .A2(n800), .ZN(n558) );
  XNOR2_X1 U616 ( .A(KEYINPUT69), .B(n558), .ZN(n559) );
  NOR2_X1 U617 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U618 ( .A(KEYINPUT70), .B(n561), .ZN(G171) );
  NAND2_X1 U619 ( .A1(n800), .A2(G51), .ZN(n562) );
  XNOR2_X1 U620 ( .A(KEYINPUT77), .B(n562), .ZN(n565) );
  NAND2_X1 U621 ( .A1(n793), .A2(G63), .ZN(n563) );
  XOR2_X1 U622 ( .A(KEYINPUT76), .B(n563), .Z(n564) );
  NOR2_X1 U623 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U624 ( .A(n566), .B(KEYINPUT6), .ZN(n572) );
  NAND2_X1 U625 ( .A1(n792), .A2(G89), .ZN(n567) );
  XNOR2_X1 U626 ( .A(n567), .B(KEYINPUT4), .ZN(n569) );
  NAND2_X1 U627 ( .A1(G76), .A2(n796), .ZN(n568) );
  NAND2_X1 U628 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U629 ( .A(KEYINPUT5), .B(n570), .ZN(n571) );
  NAND2_X1 U630 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U631 ( .A(n573), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U632 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U633 ( .A1(G88), .A2(n792), .ZN(n574) );
  XNOR2_X1 U634 ( .A(n574), .B(KEYINPUT84), .ZN(n581) );
  NAND2_X1 U635 ( .A1(G75), .A2(n796), .ZN(n576) );
  NAND2_X1 U636 ( .A1(G50), .A2(n800), .ZN(n575) );
  NAND2_X1 U637 ( .A1(n576), .A2(n575), .ZN(n579) );
  NAND2_X1 U638 ( .A1(G62), .A2(n793), .ZN(n577) );
  XNOR2_X1 U639 ( .A(KEYINPUT83), .B(n577), .ZN(n578) );
  NOR2_X1 U640 ( .A1(n579), .A2(n578), .ZN(n580) );
  NAND2_X1 U641 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U642 ( .A(KEYINPUT85), .B(n582), .ZN(G166) );
  XNOR2_X1 U643 ( .A(G166), .B(KEYINPUT93), .ZN(G303) );
  NAND2_X1 U644 ( .A1(G49), .A2(n800), .ZN(n585) );
  NAND2_X1 U645 ( .A1(G87), .A2(n583), .ZN(n584) );
  NAND2_X1 U646 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U647 ( .A1(n793), .A2(n586), .ZN(n588) );
  NAND2_X1 U648 ( .A1(G651), .A2(G74), .ZN(n587) );
  NAND2_X1 U649 ( .A1(n588), .A2(n587), .ZN(G288) );
  NAND2_X1 U650 ( .A1(G85), .A2(n792), .ZN(n590) );
  NAND2_X1 U651 ( .A1(G72), .A2(n796), .ZN(n589) );
  NAND2_X1 U652 ( .A1(n590), .A2(n589), .ZN(n594) );
  NAND2_X1 U653 ( .A1(G47), .A2(n800), .ZN(n592) );
  NAND2_X1 U654 ( .A1(G60), .A2(n793), .ZN(n591) );
  NAND2_X1 U655 ( .A1(n592), .A2(n591), .ZN(n593) );
  OR2_X1 U656 ( .A1(n594), .A2(n593), .ZN(G290) );
  NOR2_X1 U657 ( .A1(G164), .A2(G1384), .ZN(n725) );
  NAND2_X1 U658 ( .A1(G160), .A2(G40), .ZN(n726) );
  INV_X1 U659 ( .A(n726), .ZN(n616) );
  NAND2_X1 U660 ( .A1(n725), .A2(n616), .ZN(n663) );
  NAND2_X1 U661 ( .A1(G8), .A2(n663), .ZN(n651) );
  NOR2_X1 U662 ( .A1(G1981), .A2(G305), .ZN(n595) );
  XOR2_X1 U663 ( .A(n595), .B(KEYINPUT24), .Z(n596) );
  NOR2_X1 U664 ( .A1(n651), .A2(n596), .ZN(n692) );
  NAND2_X1 U665 ( .A1(G66), .A2(n793), .ZN(n603) );
  NAND2_X1 U666 ( .A1(G92), .A2(n792), .ZN(n598) );
  NAND2_X1 U667 ( .A1(G79), .A2(n796), .ZN(n597) );
  NAND2_X1 U668 ( .A1(n598), .A2(n597), .ZN(n601) );
  NAND2_X1 U669 ( .A1(G54), .A2(n800), .ZN(n599) );
  XNOR2_X1 U670 ( .A(KEYINPUT75), .B(n599), .ZN(n600) );
  NOR2_X1 U671 ( .A1(n601), .A2(n600), .ZN(n602) );
  NAND2_X1 U672 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U673 ( .A(n604), .B(KEYINPUT15), .ZN(n1009) );
  XNOR2_X1 U674 ( .A(KEYINPUT73), .B(KEYINPUT13), .ZN(n609) );
  NAND2_X1 U675 ( .A1(n792), .A2(G81), .ZN(n605) );
  XNOR2_X1 U676 ( .A(n605), .B(KEYINPUT12), .ZN(n607) );
  NAND2_X1 U677 ( .A1(G68), .A2(n796), .ZN(n606) );
  NAND2_X1 U678 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U679 ( .A(n609), .B(n608), .ZN(n612) );
  NAND2_X1 U680 ( .A1(n793), .A2(G56), .ZN(n610) );
  XOR2_X1 U681 ( .A(KEYINPUT14), .B(n610), .Z(n611) );
  NOR2_X1 U682 ( .A1(n612), .A2(n611), .ZN(n614) );
  NAND2_X1 U683 ( .A1(n800), .A2(G43), .ZN(n613) );
  NAND2_X1 U684 ( .A1(n614), .A2(n613), .ZN(n1008) );
  INV_X1 U685 ( .A(KEYINPUT64), .ZN(n619) );
  AND2_X1 U686 ( .A1(n725), .A2(G1996), .ZN(n615) );
  NAND2_X1 U687 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U688 ( .A(n619), .B(n618), .ZN(n623) );
  INV_X1 U689 ( .A(KEYINPUT100), .ZN(n621) );
  NAND2_X1 U690 ( .A1(G1341), .A2(n663), .ZN(n620) );
  XNOR2_X1 U691 ( .A(n621), .B(n620), .ZN(n622) );
  NOR2_X1 U692 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U693 ( .A(n624), .B(KEYINPUT101), .ZN(n625) );
  NOR2_X1 U694 ( .A1(n1008), .A2(n625), .ZN(n631) );
  NAND2_X1 U695 ( .A1(n1009), .A2(n631), .ZN(n630) );
  INV_X1 U696 ( .A(n663), .ZN(n646) );
  AND2_X1 U697 ( .A1(n646), .A2(G2067), .ZN(n626) );
  XOR2_X1 U698 ( .A(n626), .B(KEYINPUT102), .Z(n628) );
  NAND2_X1 U699 ( .A1(n663), .A2(G1348), .ZN(n627) );
  NAND2_X1 U700 ( .A1(n628), .A2(n627), .ZN(n629) );
  NAND2_X1 U701 ( .A1(n630), .A2(n629), .ZN(n633) );
  OR2_X1 U702 ( .A1(n1009), .A2(n631), .ZN(n632) );
  NAND2_X1 U703 ( .A1(n633), .A2(n632), .ZN(n638) );
  INV_X1 U704 ( .A(G299), .ZN(n807) );
  NAND2_X1 U705 ( .A1(n646), .A2(G2072), .ZN(n634) );
  XNOR2_X1 U706 ( .A(n634), .B(KEYINPUT27), .ZN(n636) );
  INV_X1 U707 ( .A(G1956), .ZN(n875) );
  NOR2_X1 U708 ( .A1(n875), .A2(n646), .ZN(n635) );
  NOR2_X1 U709 ( .A1(n636), .A2(n635), .ZN(n639) );
  NAND2_X1 U710 ( .A1(n807), .A2(n639), .ZN(n637) );
  NAND2_X1 U711 ( .A1(n638), .A2(n637), .ZN(n643) );
  NOR2_X1 U712 ( .A1(n807), .A2(n639), .ZN(n641) );
  XNOR2_X1 U713 ( .A(KEYINPUT99), .B(KEYINPUT28), .ZN(n640) );
  XNOR2_X1 U714 ( .A(n641), .B(n640), .ZN(n642) );
  NAND2_X1 U715 ( .A1(n643), .A2(n642), .ZN(n645) );
  INV_X1 U716 ( .A(G1961), .ZN(n884) );
  NAND2_X1 U717 ( .A1(n663), .A2(n884), .ZN(n648) );
  XNOR2_X1 U718 ( .A(G2078), .B(KEYINPUT25), .ZN(n900) );
  NAND2_X1 U719 ( .A1(n646), .A2(n900), .ZN(n647) );
  NAND2_X1 U720 ( .A1(n648), .A2(n647), .ZN(n657) );
  NAND2_X1 U721 ( .A1(n657), .A2(G171), .ZN(n649) );
  NAND2_X1 U722 ( .A1(n650), .A2(n649), .ZN(n662) );
  NOR2_X1 U723 ( .A1(G1966), .A2(n651), .ZN(n674) );
  NOR2_X1 U724 ( .A1(G2084), .A2(n663), .ZN(n671) );
  NOR2_X1 U725 ( .A1(n674), .A2(n671), .ZN(n652) );
  NAND2_X1 U726 ( .A1(G8), .A2(n652), .ZN(n655) );
  NOR2_X1 U727 ( .A1(G168), .A2(n656), .ZN(n659) );
  NOR2_X1 U728 ( .A1(n657), .A2(G171), .ZN(n658) );
  NOR2_X1 U729 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U730 ( .A(KEYINPUT31), .B(n660), .Z(n661) );
  NAND2_X1 U731 ( .A1(n662), .A2(n661), .ZN(n672) );
  NAND2_X1 U732 ( .A1(n672), .A2(G286), .ZN(n668) );
  NOR2_X1 U733 ( .A1(G1971), .A2(n651), .ZN(n665) );
  NOR2_X1 U734 ( .A1(G2090), .A2(n663), .ZN(n664) );
  NOR2_X1 U735 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U736 ( .A1(n666), .A2(G303), .ZN(n667) );
  NAND2_X1 U737 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U738 ( .A(n670), .B(KEYINPUT32), .ZN(n678) );
  NAND2_X1 U739 ( .A1(G8), .A2(n671), .ZN(n676) );
  INV_X1 U740 ( .A(n672), .ZN(n673) );
  NOR2_X1 U741 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U742 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U743 ( .A1(n678), .A2(n677), .ZN(n695) );
  NOR2_X1 U744 ( .A1(G1976), .A2(G288), .ZN(n684) );
  NOR2_X1 U745 ( .A1(G1971), .A2(G303), .ZN(n679) );
  NOR2_X1 U746 ( .A1(n684), .A2(n679), .ZN(n865) );
  NAND2_X1 U747 ( .A1(n695), .A2(n865), .ZN(n680) );
  NAND2_X1 U748 ( .A1(G1976), .A2(G288), .ZN(n852) );
  NAND2_X1 U749 ( .A1(n680), .A2(n852), .ZN(n681) );
  NOR2_X1 U750 ( .A1(KEYINPUT33), .A2(n681), .ZN(n682) );
  INV_X1 U751 ( .A(n651), .ZN(n683) );
  NAND2_X1 U752 ( .A1(n682), .A2(n683), .ZN(n687) );
  NAND2_X1 U753 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U754 ( .A1(n685), .A2(KEYINPUT33), .ZN(n686) );
  NAND2_X1 U755 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U756 ( .A(G1981), .B(G305), .ZN(n855) );
  NOR2_X1 U757 ( .A1(n692), .A2(n691), .ZN(n731) );
  NOR2_X1 U758 ( .A1(G2090), .A2(G303), .ZN(n693) );
  NAND2_X1 U759 ( .A1(G8), .A2(n693), .ZN(n694) );
  NAND2_X1 U760 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U761 ( .A1(n651), .A2(n696), .ZN(n729) );
  INV_X1 U762 ( .A(G1996), .ZN(n716) );
  NAND2_X1 U763 ( .A1(G117), .A2(n991), .ZN(n698) );
  NAND2_X1 U764 ( .A1(G141), .A2(n995), .ZN(n697) );
  NAND2_X1 U765 ( .A1(n698), .A2(n697), .ZN(n707) );
  BUF_X1 U766 ( .A(n699), .Z(n994) );
  NAND2_X1 U767 ( .A1(G105), .A2(n994), .ZN(n700) );
  XNOR2_X1 U768 ( .A(n700), .B(KEYINPUT38), .ZN(n701) );
  XNOR2_X1 U769 ( .A(KEYINPUT98), .B(n701), .ZN(n705) );
  NAND2_X1 U770 ( .A1(G129), .A2(n702), .ZN(n703) );
  XOR2_X1 U771 ( .A(KEYINPUT97), .B(n703), .Z(n704) );
  NAND2_X1 U772 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U773 ( .A1(n707), .A2(n706), .ZN(n979) );
  AND2_X1 U774 ( .A1(n716), .A2(n979), .ZN(n940) );
  INV_X1 U775 ( .A(G1991), .ZN(n898) );
  NAND2_X1 U776 ( .A1(n702), .A2(G119), .ZN(n714) );
  NAND2_X1 U777 ( .A1(G107), .A2(n991), .ZN(n709) );
  NAND2_X1 U778 ( .A1(G131), .A2(n995), .ZN(n708) );
  NAND2_X1 U779 ( .A1(n709), .A2(n708), .ZN(n712) );
  NAND2_X1 U780 ( .A1(G95), .A2(n994), .ZN(n710) );
  XNOR2_X1 U781 ( .A(KEYINPUT95), .B(n710), .ZN(n711) );
  NOR2_X1 U782 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U783 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U784 ( .A(KEYINPUT96), .B(n715), .Z(n719) );
  NOR2_X1 U785 ( .A1(n898), .A2(n719), .ZN(n718) );
  NOR2_X1 U786 ( .A1(n716), .A2(n979), .ZN(n717) );
  NOR2_X1 U787 ( .A1(n718), .A2(n717), .ZN(n742) );
  INV_X1 U788 ( .A(n742), .ZN(n933) );
  NOR2_X1 U789 ( .A1(G1986), .A2(G290), .ZN(n720) );
  INV_X1 U790 ( .A(n719), .ZN(n980) );
  NOR2_X1 U791 ( .A1(G1991), .A2(n980), .ZN(n931) );
  NOR2_X1 U792 ( .A1(n720), .A2(n931), .ZN(n721) );
  XOR2_X1 U793 ( .A(KEYINPUT105), .B(n721), .Z(n722) );
  NOR2_X1 U794 ( .A1(n933), .A2(n722), .ZN(n723) );
  NOR2_X1 U795 ( .A1(n940), .A2(n723), .ZN(n724) );
  XNOR2_X1 U796 ( .A(KEYINPUT39), .B(n724), .ZN(n728) );
  NOR2_X1 U797 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U798 ( .A(n727), .B(KEYINPUT94), .ZN(n752) );
  NAND2_X1 U799 ( .A1(n728), .A2(n752), .ZN(n741) );
  AND2_X1 U800 ( .A1(n729), .A2(n741), .ZN(n730) );
  NAND2_X1 U801 ( .A1(n731), .A2(n730), .ZN(n749) );
  NAND2_X1 U802 ( .A1(n995), .A2(G140), .ZN(n733) );
  NAND2_X1 U803 ( .A1(n994), .A2(G104), .ZN(n732) );
  NAND2_X1 U804 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U805 ( .A(KEYINPUT34), .B(n734), .ZN(n739) );
  NAND2_X1 U806 ( .A1(G128), .A2(n702), .ZN(n736) );
  NAND2_X1 U807 ( .A1(G116), .A2(n991), .ZN(n735) );
  NAND2_X1 U808 ( .A1(n736), .A2(n735), .ZN(n737) );
  XOR2_X1 U809 ( .A(KEYINPUT35), .B(n737), .Z(n738) );
  NOR2_X1 U810 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U811 ( .A(KEYINPUT36), .B(n740), .ZN(n981) );
  XNOR2_X1 U812 ( .A(G2067), .B(KEYINPUT37), .ZN(n750) );
  NOR2_X1 U813 ( .A1(n981), .A2(n750), .ZN(n932) );
  NAND2_X1 U814 ( .A1(n932), .A2(n752), .ZN(n747) );
  INV_X1 U815 ( .A(n741), .ZN(n745) );
  XOR2_X1 U816 ( .A(G1986), .B(G290), .Z(n848) );
  NAND2_X1 U817 ( .A1(n742), .A2(n848), .ZN(n743) );
  NAND2_X1 U818 ( .A1(n743), .A2(n752), .ZN(n744) );
  OR2_X1 U819 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U820 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U821 ( .A1(n749), .A2(n748), .ZN(n754) );
  AND2_X1 U822 ( .A1(n750), .A2(n981), .ZN(n751) );
  XNOR2_X1 U823 ( .A(n751), .B(KEYINPUT106), .ZN(n943) );
  NAND2_X1 U824 ( .A1(n943), .A2(n752), .ZN(n753) );
  NAND2_X1 U825 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U826 ( .A(n755), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U827 ( .A(G1348), .B(G2427), .ZN(n765) );
  XOR2_X1 U828 ( .A(G2451), .B(G2430), .Z(n757) );
  XNOR2_X1 U829 ( .A(G1341), .B(G2443), .ZN(n756) );
  XNOR2_X1 U830 ( .A(n757), .B(n756), .ZN(n761) );
  XOR2_X1 U831 ( .A(G2438), .B(G2435), .Z(n759) );
  XNOR2_X1 U832 ( .A(KEYINPUT107), .B(G2454), .ZN(n758) );
  XNOR2_X1 U833 ( .A(n759), .B(n758), .ZN(n760) );
  XOR2_X1 U834 ( .A(n761), .B(n760), .Z(n763) );
  XNOR2_X1 U835 ( .A(G2446), .B(KEYINPUT108), .ZN(n762) );
  XNOR2_X1 U836 ( .A(n763), .B(n762), .ZN(n764) );
  XNOR2_X1 U837 ( .A(n765), .B(n764), .ZN(n766) );
  AND2_X1 U838 ( .A1(n766), .A2(G14), .ZN(G401) );
  AND2_X1 U839 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U840 ( .A1(G123), .A2(n702), .ZN(n767) );
  XNOR2_X1 U841 ( .A(n767), .B(KEYINPUT18), .ZN(n774) );
  NAND2_X1 U842 ( .A1(G111), .A2(n991), .ZN(n769) );
  NAND2_X1 U843 ( .A1(G99), .A2(n994), .ZN(n768) );
  NAND2_X1 U844 ( .A1(n769), .A2(n768), .ZN(n772) );
  NAND2_X1 U845 ( .A1(G135), .A2(n995), .ZN(n770) );
  XNOR2_X1 U846 ( .A(KEYINPUT79), .B(n770), .ZN(n771) );
  NOR2_X1 U847 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U848 ( .A1(n774), .A2(n773), .ZN(n985) );
  XNOR2_X1 U849 ( .A(G2096), .B(n985), .ZN(n775) );
  OR2_X1 U850 ( .A1(G2100), .A2(n775), .ZN(G156) );
  INV_X1 U851 ( .A(G132), .ZN(G219) );
  INV_X1 U852 ( .A(G82), .ZN(G220) );
  INV_X1 U853 ( .A(G120), .ZN(G236) );
  INV_X1 U854 ( .A(G69), .ZN(G235) );
  INV_X1 U855 ( .A(G108), .ZN(G238) );
  NAND2_X1 U856 ( .A1(G7), .A2(G661), .ZN(n776) );
  XNOR2_X1 U857 ( .A(n776), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U858 ( .A(G223), .ZN(n834) );
  NAND2_X1 U859 ( .A1(n834), .A2(G567), .ZN(n777) );
  XOR2_X1 U860 ( .A(KEYINPUT11), .B(n777), .Z(G234) );
  INV_X1 U861 ( .A(G860), .ZN(n783) );
  NOR2_X1 U862 ( .A1(n1008), .A2(n783), .ZN(n778) );
  XOR2_X1 U863 ( .A(KEYINPUT74), .B(n778), .Z(G153) );
  INV_X1 U864 ( .A(G171), .ZN(G301) );
  NAND2_X1 U865 ( .A1(G301), .A2(G868), .ZN(n780) );
  OR2_X1 U866 ( .A1(n1009), .A2(G868), .ZN(n779) );
  NAND2_X1 U867 ( .A1(n780), .A2(n779), .ZN(G284) );
  INV_X1 U868 ( .A(G868), .ZN(n815) );
  NOR2_X1 U869 ( .A1(G286), .A2(n815), .ZN(n782) );
  NOR2_X1 U870 ( .A1(G868), .A2(G299), .ZN(n781) );
  NOR2_X1 U871 ( .A1(n782), .A2(n781), .ZN(G297) );
  NAND2_X1 U872 ( .A1(G559), .A2(n783), .ZN(n784) );
  XNOR2_X1 U873 ( .A(KEYINPUT78), .B(n784), .ZN(n785) );
  NAND2_X1 U874 ( .A1(n785), .A2(n1009), .ZN(n786) );
  XNOR2_X1 U875 ( .A(KEYINPUT16), .B(n786), .ZN(G148) );
  NOR2_X1 U876 ( .A1(G868), .A2(n1008), .ZN(n789) );
  NAND2_X1 U877 ( .A1(G868), .A2(n1009), .ZN(n787) );
  NOR2_X1 U878 ( .A1(G559), .A2(n787), .ZN(n788) );
  NOR2_X1 U879 ( .A1(n789), .A2(n788), .ZN(G282) );
  NAND2_X1 U880 ( .A1(G559), .A2(n1009), .ZN(n790) );
  XNOR2_X1 U881 ( .A(n790), .B(n1008), .ZN(n812) );
  XNOR2_X1 U882 ( .A(KEYINPUT80), .B(n812), .ZN(n791) );
  NOR2_X1 U883 ( .A1(G860), .A2(n791), .ZN(n803) );
  NAND2_X1 U884 ( .A1(G93), .A2(n792), .ZN(n795) );
  NAND2_X1 U885 ( .A1(G67), .A2(n793), .ZN(n794) );
  NAND2_X1 U886 ( .A1(n795), .A2(n794), .ZN(n799) );
  NAND2_X1 U887 ( .A1(G80), .A2(n796), .ZN(n797) );
  XNOR2_X1 U888 ( .A(KEYINPUT81), .B(n797), .ZN(n798) );
  NOR2_X1 U889 ( .A1(n799), .A2(n798), .ZN(n802) );
  NAND2_X1 U890 ( .A1(n800), .A2(G55), .ZN(n801) );
  NAND2_X1 U891 ( .A1(n802), .A2(n801), .ZN(n814) );
  XOR2_X1 U892 ( .A(n803), .B(n814), .Z(G145) );
  XNOR2_X1 U893 ( .A(G166), .B(G305), .ZN(n811) );
  XNOR2_X1 U894 ( .A(KEYINPUT19), .B(KEYINPUT86), .ZN(n805) );
  XNOR2_X1 U895 ( .A(G288), .B(KEYINPUT87), .ZN(n804) );
  XNOR2_X1 U896 ( .A(n805), .B(n804), .ZN(n806) );
  XNOR2_X1 U897 ( .A(n807), .B(n806), .ZN(n809) );
  XNOR2_X1 U898 ( .A(G290), .B(n814), .ZN(n808) );
  XNOR2_X1 U899 ( .A(n809), .B(n808), .ZN(n810) );
  XNOR2_X1 U900 ( .A(n811), .B(n810), .ZN(n1007) );
  XNOR2_X1 U901 ( .A(n812), .B(n1007), .ZN(n813) );
  NAND2_X1 U902 ( .A1(n813), .A2(G868), .ZN(n817) );
  NAND2_X1 U903 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U904 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U905 ( .A(KEYINPUT88), .B(n818), .ZN(G295) );
  NAND2_X1 U906 ( .A1(G2078), .A2(G2084), .ZN(n819) );
  XOR2_X1 U907 ( .A(KEYINPUT20), .B(n819), .Z(n820) );
  NAND2_X1 U908 ( .A1(G2090), .A2(n820), .ZN(n821) );
  XNOR2_X1 U909 ( .A(n821), .B(KEYINPUT90), .ZN(n823) );
  XOR2_X1 U910 ( .A(KEYINPUT21), .B(KEYINPUT89), .Z(n822) );
  XNOR2_X1 U911 ( .A(n823), .B(n822), .ZN(n824) );
  NAND2_X1 U912 ( .A1(n824), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U913 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U914 ( .A1(G235), .A2(G236), .ZN(n825) );
  XNOR2_X1 U915 ( .A(n825), .B(KEYINPUT91), .ZN(n826) );
  NOR2_X1 U916 ( .A1(G238), .A2(n826), .ZN(n827) );
  NAND2_X1 U917 ( .A1(G57), .A2(n827), .ZN(n955) );
  NAND2_X1 U918 ( .A1(G567), .A2(n955), .ZN(n832) );
  NOR2_X1 U919 ( .A1(G220), .A2(G219), .ZN(n828) );
  XOR2_X1 U920 ( .A(KEYINPUT22), .B(n828), .Z(n829) );
  NOR2_X1 U921 ( .A1(G218), .A2(n829), .ZN(n830) );
  NAND2_X1 U922 ( .A1(G96), .A2(n830), .ZN(n956) );
  NAND2_X1 U923 ( .A1(G2106), .A2(n956), .ZN(n831) );
  NAND2_X1 U924 ( .A1(n832), .A2(n831), .ZN(n978) );
  NAND2_X1 U925 ( .A1(G483), .A2(G661), .ZN(n833) );
  NOR2_X1 U926 ( .A1(n978), .A2(n833), .ZN(n838) );
  NAND2_X1 U927 ( .A1(n838), .A2(G36), .ZN(G176) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n834), .ZN(G217) );
  NAND2_X1 U929 ( .A1(G15), .A2(G2), .ZN(n835) );
  XNOR2_X1 U930 ( .A(KEYINPUT109), .B(n835), .ZN(n836) );
  NAND2_X1 U931 ( .A1(n836), .A2(G661), .ZN(G259) );
  NAND2_X1 U932 ( .A1(G3), .A2(G1), .ZN(n837) );
  NAND2_X1 U933 ( .A1(n838), .A2(n837), .ZN(G188) );
  NAND2_X1 U935 ( .A1(G112), .A2(n991), .ZN(n840) );
  NAND2_X1 U936 ( .A1(G100), .A2(n994), .ZN(n839) );
  NAND2_X1 U937 ( .A1(n840), .A2(n839), .ZN(n841) );
  XNOR2_X1 U938 ( .A(KEYINPUT116), .B(n841), .ZN(n847) );
  NAND2_X1 U939 ( .A1(n702), .A2(G124), .ZN(n842) );
  XNOR2_X1 U940 ( .A(n842), .B(KEYINPUT44), .ZN(n844) );
  NAND2_X1 U941 ( .A1(G136), .A2(n995), .ZN(n843) );
  NAND2_X1 U942 ( .A1(n844), .A2(n843), .ZN(n845) );
  XOR2_X1 U943 ( .A(KEYINPUT115), .B(n845), .Z(n846) );
  NOR2_X1 U944 ( .A1(n847), .A2(n846), .ZN(G162) );
  XNOR2_X1 U945 ( .A(G16), .B(KEYINPUT56), .ZN(n868) );
  XNOR2_X1 U946 ( .A(G301), .B(n884), .ZN(n849) );
  NAND2_X1 U947 ( .A1(n849), .A2(n848), .ZN(n851) );
  XNOR2_X1 U948 ( .A(G1341), .B(n1008), .ZN(n850) );
  NOR2_X1 U949 ( .A1(n851), .A2(n850), .ZN(n853) );
  NAND2_X1 U950 ( .A1(n853), .A2(n852), .ZN(n864) );
  XOR2_X1 U951 ( .A(G168), .B(G1966), .Z(n854) );
  NOR2_X1 U952 ( .A1(n855), .A2(n854), .ZN(n856) );
  XOR2_X1 U953 ( .A(KEYINPUT57), .B(n856), .Z(n862) );
  XNOR2_X1 U954 ( .A(G1348), .B(n1009), .ZN(n858) );
  NAND2_X1 U955 ( .A1(G1971), .A2(G303), .ZN(n857) );
  NAND2_X1 U956 ( .A1(n858), .A2(n857), .ZN(n860) );
  XNOR2_X1 U957 ( .A(G1956), .B(G299), .ZN(n859) );
  NOR2_X1 U958 ( .A1(n860), .A2(n859), .ZN(n861) );
  NAND2_X1 U959 ( .A1(n862), .A2(n861), .ZN(n863) );
  NOR2_X1 U960 ( .A1(n864), .A2(n863), .ZN(n866) );
  NAND2_X1 U961 ( .A1(n866), .A2(n865), .ZN(n867) );
  NAND2_X1 U962 ( .A1(n868), .A2(n867), .ZN(n869) );
  XNOR2_X1 U963 ( .A(KEYINPUT124), .B(n869), .ZN(n953) );
  XOR2_X1 U964 ( .A(G1986), .B(G24), .Z(n871) );
  XOR2_X1 U965 ( .A(G1971), .B(G22), .Z(n870) );
  NAND2_X1 U966 ( .A1(n871), .A2(n870), .ZN(n873) );
  XNOR2_X1 U967 ( .A(G23), .B(G1976), .ZN(n872) );
  NOR2_X1 U968 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U969 ( .A(KEYINPUT58), .B(n874), .Z(n891) );
  XNOR2_X1 U970 ( .A(G20), .B(n875), .ZN(n879) );
  XNOR2_X1 U971 ( .A(G1341), .B(G19), .ZN(n877) );
  XNOR2_X1 U972 ( .A(G6), .B(G1981), .ZN(n876) );
  NOR2_X1 U973 ( .A1(n877), .A2(n876), .ZN(n878) );
  NAND2_X1 U974 ( .A1(n879), .A2(n878), .ZN(n882) );
  XOR2_X1 U975 ( .A(KEYINPUT59), .B(G1348), .Z(n880) );
  XNOR2_X1 U976 ( .A(G4), .B(n880), .ZN(n881) );
  NOR2_X1 U977 ( .A1(n882), .A2(n881), .ZN(n883) );
  XNOR2_X1 U978 ( .A(KEYINPUT60), .B(n883), .ZN(n886) );
  XNOR2_X1 U979 ( .A(n884), .B(G5), .ZN(n885) );
  NAND2_X1 U980 ( .A1(n886), .A2(n885), .ZN(n888) );
  XNOR2_X1 U981 ( .A(G21), .B(G1966), .ZN(n887) );
  NOR2_X1 U982 ( .A1(n888), .A2(n887), .ZN(n889) );
  XNOR2_X1 U983 ( .A(KEYINPUT125), .B(n889), .ZN(n890) );
  NOR2_X1 U984 ( .A1(n891), .A2(n890), .ZN(n892) );
  XNOR2_X1 U985 ( .A(KEYINPUT126), .B(n892), .ZN(n893) );
  XNOR2_X1 U986 ( .A(n893), .B(KEYINPUT61), .ZN(n895) );
  INV_X1 U987 ( .A(G16), .ZN(n894) );
  NAND2_X1 U988 ( .A1(n895), .A2(n894), .ZN(n896) );
  NAND2_X1 U989 ( .A1(G11), .A2(n896), .ZN(n951) );
  XNOR2_X1 U990 ( .A(G2084), .B(G34), .ZN(n897) );
  XNOR2_X1 U991 ( .A(n897), .B(KEYINPUT54), .ZN(n915) );
  XNOR2_X1 U992 ( .A(G2090), .B(G35), .ZN(n912) );
  XNOR2_X1 U993 ( .A(G25), .B(n898), .ZN(n899) );
  NAND2_X1 U994 ( .A1(n899), .A2(G28), .ZN(n909) );
  XOR2_X1 U995 ( .A(n900), .B(G27), .Z(n902) );
  XNOR2_X1 U996 ( .A(G32), .B(G1996), .ZN(n901) );
  NOR2_X1 U997 ( .A1(n902), .A2(n901), .ZN(n903) );
  XNOR2_X1 U998 ( .A(KEYINPUT122), .B(n903), .ZN(n907) );
  XNOR2_X1 U999 ( .A(G2067), .B(G26), .ZN(n905) );
  XNOR2_X1 U1000 ( .A(G33), .B(G2072), .ZN(n904) );
  NOR2_X1 U1001 ( .A1(n905), .A2(n904), .ZN(n906) );
  NAND2_X1 U1002 ( .A1(n907), .A2(n906), .ZN(n908) );
  NOR2_X1 U1003 ( .A1(n909), .A2(n908), .ZN(n910) );
  XNOR2_X1 U1004 ( .A(KEYINPUT53), .B(n910), .ZN(n911) );
  NOR2_X1 U1005 ( .A1(n912), .A2(n911), .ZN(n913) );
  XNOR2_X1 U1006 ( .A(n913), .B(KEYINPUT123), .ZN(n914) );
  NOR2_X1 U1007 ( .A1(n915), .A2(n914), .ZN(n916) );
  NOR2_X1 U1008 ( .A1(G29), .A2(n916), .ZN(n917) );
  XNOR2_X1 U1009 ( .A(n917), .B(KEYINPUT55), .ZN(n949) );
  NAND2_X1 U1010 ( .A1(G103), .A2(n994), .ZN(n919) );
  NAND2_X1 U1011 ( .A1(G139), .A2(n995), .ZN(n918) );
  NAND2_X1 U1012 ( .A1(n919), .A2(n918), .ZN(n924) );
  NAND2_X1 U1013 ( .A1(G127), .A2(n702), .ZN(n921) );
  NAND2_X1 U1014 ( .A1(G115), .A2(n991), .ZN(n920) );
  NAND2_X1 U1015 ( .A1(n921), .A2(n920), .ZN(n922) );
  XOR2_X1 U1016 ( .A(KEYINPUT47), .B(n922), .Z(n923) );
  NOR2_X1 U1017 ( .A1(n924), .A2(n923), .ZN(n986) );
  XNOR2_X1 U1018 ( .A(G2072), .B(n986), .ZN(n927) );
  XOR2_X1 U1019 ( .A(G164), .B(G2078), .Z(n925) );
  XNOR2_X1 U1020 ( .A(KEYINPUT121), .B(n925), .ZN(n926) );
  NAND2_X1 U1021 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1022 ( .A(n928), .B(KEYINPUT50), .ZN(n938) );
  XNOR2_X1 U1023 ( .A(G160), .B(G2084), .ZN(n929) );
  NAND2_X1 U1024 ( .A1(n929), .A2(n985), .ZN(n930) );
  NOR2_X1 U1025 ( .A1(n931), .A2(n930), .ZN(n935) );
  NOR2_X1 U1026 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1027 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1028 ( .A(KEYINPUT120), .B(n936), .ZN(n937) );
  NOR2_X1 U1029 ( .A1(n938), .A2(n937), .ZN(n945) );
  XOR2_X1 U1030 ( .A(G2090), .B(G162), .Z(n939) );
  NOR2_X1 U1031 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1032 ( .A(n941), .B(KEYINPUT51), .ZN(n942) );
  NOR2_X1 U1033 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1034 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1035 ( .A(KEYINPUT52), .B(n946), .ZN(n947) );
  NAND2_X1 U1036 ( .A1(G29), .A2(n947), .ZN(n948) );
  NAND2_X1 U1037 ( .A1(n949), .A2(n948), .ZN(n950) );
  NOR2_X1 U1038 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1039 ( .A1(n953), .A2(n952), .ZN(n954) );
  XOR2_X1 U1040 ( .A(KEYINPUT62), .B(n954), .Z(G311) );
  XNOR2_X1 U1041 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1042 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1043 ( .A1(n956), .A2(n955), .ZN(G325) );
  INV_X1 U1044 ( .A(G325), .ZN(G261) );
  XOR2_X1 U1045 ( .A(KEYINPUT113), .B(KEYINPUT42), .Z(n958) );
  XNOR2_X1 U1046 ( .A(G2072), .B(G2096), .ZN(n957) );
  XNOR2_X1 U1047 ( .A(n958), .B(n957), .ZN(n968) );
  XOR2_X1 U1048 ( .A(KEYINPUT114), .B(G2678), .Z(n960) );
  XNOR2_X1 U1049 ( .A(G2090), .B(KEYINPUT111), .ZN(n959) );
  XNOR2_X1 U1050 ( .A(n960), .B(n959), .ZN(n964) );
  XOR2_X1 U1051 ( .A(KEYINPUT112), .B(G2100), .Z(n962) );
  XNOR2_X1 U1052 ( .A(G2067), .B(KEYINPUT43), .ZN(n961) );
  XNOR2_X1 U1053 ( .A(n962), .B(n961), .ZN(n963) );
  XOR2_X1 U1054 ( .A(n964), .B(n963), .Z(n966) );
  XNOR2_X1 U1055 ( .A(G2078), .B(G2084), .ZN(n965) );
  XNOR2_X1 U1056 ( .A(n966), .B(n965), .ZN(n967) );
  XOR2_X1 U1057 ( .A(n968), .B(n967), .Z(G227) );
  XOR2_X1 U1058 ( .A(G1986), .B(G1971), .Z(n970) );
  XNOR2_X1 U1059 ( .A(G1961), .B(G1996), .ZN(n969) );
  XNOR2_X1 U1060 ( .A(n970), .B(n969), .ZN(n971) );
  XOR2_X1 U1061 ( .A(n971), .B(KEYINPUT41), .Z(n973) );
  XNOR2_X1 U1062 ( .A(G1966), .B(G1976), .ZN(n972) );
  XNOR2_X1 U1063 ( .A(n973), .B(n972), .ZN(n977) );
  XOR2_X1 U1064 ( .A(G2474), .B(G1991), .Z(n975) );
  XNOR2_X1 U1065 ( .A(G1956), .B(G1981), .ZN(n974) );
  XNOR2_X1 U1066 ( .A(n975), .B(n974), .ZN(n976) );
  XNOR2_X1 U1067 ( .A(n977), .B(n976), .ZN(G229) );
  XOR2_X1 U1068 ( .A(KEYINPUT110), .B(n978), .Z(G319) );
  XOR2_X1 U1069 ( .A(n980), .B(n979), .Z(n983) );
  XOR2_X1 U1070 ( .A(n981), .B(G160), .Z(n982) );
  XNOR2_X1 U1071 ( .A(n983), .B(n982), .ZN(n984) );
  XNOR2_X1 U1072 ( .A(n985), .B(n984), .ZN(n988) );
  XNOR2_X1 U1073 ( .A(G162), .B(n986), .ZN(n987) );
  XNOR2_X1 U1074 ( .A(n988), .B(n987), .ZN(n1005) );
  XOR2_X1 U1075 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n990) );
  XNOR2_X1 U1076 ( .A(KEYINPUT118), .B(KEYINPUT117), .ZN(n989) );
  XNOR2_X1 U1077 ( .A(n990), .B(n989), .ZN(n1002) );
  NAND2_X1 U1078 ( .A1(G130), .A2(n702), .ZN(n993) );
  NAND2_X1 U1079 ( .A1(G118), .A2(n991), .ZN(n992) );
  NAND2_X1 U1080 ( .A1(n993), .A2(n992), .ZN(n1000) );
  NAND2_X1 U1081 ( .A1(G106), .A2(n994), .ZN(n997) );
  NAND2_X1 U1082 ( .A1(G142), .A2(n995), .ZN(n996) );
  NAND2_X1 U1083 ( .A1(n997), .A2(n996), .ZN(n998) );
  XOR2_X1 U1084 ( .A(n998), .B(KEYINPUT45), .Z(n999) );
  NOR2_X1 U1085 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1086 ( .A(n1002), .B(n1001), .Z(n1003) );
  XOR2_X1 U1087 ( .A(G164), .B(n1003), .Z(n1004) );
  XNOR2_X1 U1088 ( .A(n1005), .B(n1004), .ZN(n1006) );
  NOR2_X1 U1089 ( .A1(G37), .A2(n1006), .ZN(G395) );
  XNOR2_X1 U1090 ( .A(n1008), .B(n1007), .ZN(n1011) );
  XNOR2_X1 U1091 ( .A(G301), .B(n1009), .ZN(n1010) );
  XNOR2_X1 U1092 ( .A(n1011), .B(n1010), .ZN(n1012) );
  XNOR2_X1 U1093 ( .A(G286), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1094 ( .A1(G37), .A2(n1013), .ZN(G397) );
  NOR2_X1 U1095 ( .A1(G227), .A2(G229), .ZN(n1014) );
  XNOR2_X1 U1096 ( .A(n1014), .B(KEYINPUT49), .ZN(n1015) );
  NOR2_X1 U1097 ( .A1(G401), .A2(n1015), .ZN(n1016) );
  NAND2_X1 U1098 ( .A1(n1016), .A2(G319), .ZN(n1017) );
  XNOR2_X1 U1099 ( .A(KEYINPUT119), .B(n1017), .ZN(n1019) );
  NOR2_X1 U1100 ( .A1(G395), .A2(G397), .ZN(n1018) );
  NAND2_X1 U1101 ( .A1(n1019), .A2(n1018), .ZN(G225) );
  INV_X1 U1102 ( .A(G225), .ZN(G308) );
  INV_X1 U1103 ( .A(G57), .ZN(G237) );
endmodule

