//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 0 0 0 0 0 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 0 1 1 1 1 0 0 1 0 0 1 0 1 1 1 0 1 0 0 0 1 1 0 0 0 1 1 1 0 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n816, new_n817, new_n818, new_n820, new_n821,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202));
  XOR2_X1   g001(.A(new_n202), .B(KEYINPUT13), .Z(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT83), .ZN(new_n205));
  XNOR2_X1  g004(.A(G15gat), .B(G22gat), .ZN(new_n206));
  OR2_X1    g005(.A1(new_n206), .A2(G1gat), .ZN(new_n207));
  INV_X1    g006(.A(G8gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT16), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n206), .B1(new_n209), .B2(G1gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n207), .A2(new_n208), .A3(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n208), .B1(new_n207), .B2(new_n210), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n205), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n213), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n215), .A2(KEYINPUT83), .A3(new_n211), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  NOR2_X1   g016(.A1(G29gat), .A2(G36gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT14), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n218), .B(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(G29gat), .A2(G36gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G43gat), .B(G50gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT15), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  OR2_X1    g025(.A1(new_n223), .A2(KEYINPUT15), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n221), .B(KEYINPUT82), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n227), .A2(new_n220), .A3(new_n224), .A4(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n217), .A2(new_n226), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n226), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n214), .A2(new_n216), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n204), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT84), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(G113gat), .B(G141gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n236), .B(G197gat), .ZN(new_n237));
  XOR2_X1   g036(.A(KEYINPUT11), .B(G169gat), .Z(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n239), .B(KEYINPUT12), .Z(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT17), .ZN(new_n242));
  AND3_X1   g041(.A1(new_n229), .A2(new_n226), .A3(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n242), .B1(new_n229), .B2(new_n226), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n215), .B(new_n211), .C1(new_n243), .C2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n245), .A2(new_n232), .A3(new_n202), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT18), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  OR2_X1    g047(.A1(new_n246), .A2(new_n247), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n235), .A2(new_n241), .A3(new_n248), .A4(new_n249), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n233), .A2(new_n234), .ZN(new_n251));
  AOI211_X1 g050(.A(KEYINPUT84), .B(new_n204), .C1(new_n230), .C2(new_n232), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n249), .A2(new_n248), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n240), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n250), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G57gat), .B(G64gat), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT9), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(G71gat), .ZN(new_n260));
  INV_X1    g059(.A(G78gat), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NOR2_X1   g061(.A1(G71gat), .A2(G78gat), .ZN(new_n263));
  NOR3_X1   g062(.A1(new_n259), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n257), .A2(KEYINPUT85), .ZN(new_n266));
  OR2_X1    g065(.A1(G57gat), .A2(G64gat), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT85), .ZN(new_n268));
  NAND2_X1  g067(.A1(G57gat), .A2(G64gat), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n266), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n262), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n263), .A2(KEYINPUT9), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n271), .A2(KEYINPUT86), .A3(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(KEYINPUT86), .B1(new_n271), .B2(new_n274), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n265), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT21), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(G231gat), .A2(G233gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n280), .B(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(G127gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n217), .B1(new_n279), .B2(new_n278), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n284), .B(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n287), .B(G155gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(G183gat), .B(G211gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  OR2_X1    g089(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n286), .A2(new_n290), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(G99gat), .A2(G106gat), .ZN(new_n294));
  INV_X1    g093(.A(G85gat), .ZN(new_n295));
  INV_X1    g094(.A(G92gat), .ZN(new_n296));
  AOI22_X1  g095(.A1(KEYINPUT8), .A2(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND4_X1  g096(.A1(KEYINPUT87), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n298));
  NAND3_X1  g097(.A1(KEYINPUT87), .A2(G85gat), .A3(G92gat), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT7), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n297), .A2(new_n298), .A3(new_n301), .ZN(new_n302));
  OR2_X1    g101(.A1(G99gat), .A2(G106gat), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n302), .A2(new_n294), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT88), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n294), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n297), .A2(new_n306), .A3(new_n298), .A4(new_n301), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n304), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  OR2_X1    g107(.A1(new_n307), .A2(new_n305), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(new_n231), .ZN(new_n311));
  AND2_X1   g110(.A1(G232gat), .A2(G233gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT41), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n243), .A2(new_n244), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n311), .B(new_n313), .C1(new_n314), .C2(new_n310), .ZN(new_n315));
  XNOR2_X1  g114(.A(G190gat), .B(G218gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n315), .A2(new_n316), .ZN(new_n319));
  AOI21_X1  g118(.A(KEYINPUT89), .B1(new_n315), .B2(new_n316), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n312), .A2(KEYINPUT41), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n321), .B(G134gat), .ZN(new_n322));
  INV_X1    g121(.A(G162gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n322), .B(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  OAI22_X1  g124(.A1(new_n318), .A2(new_n319), .B1(new_n320), .B2(new_n325), .ZN(new_n326));
  OR2_X1    g125(.A1(new_n315), .A2(new_n316), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n327), .A2(new_n317), .A3(KEYINPUT89), .A4(new_n324), .ZN(new_n328));
  AND2_X1   g127(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n293), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(G230gat), .A2(G233gat), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT90), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n278), .A2(new_n334), .A3(new_n309), .A4(new_n308), .ZN(new_n335));
  INV_X1    g134(.A(new_n270), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n268), .B1(new_n267), .B2(new_n269), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n274), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT86), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n264), .B1(new_n340), .B2(new_n275), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT90), .B1(new_n341), .B2(new_n310), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT10), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n341), .A2(new_n307), .A3(new_n304), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n335), .A2(new_n342), .A3(new_n343), .A4(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n341), .A2(new_n310), .A3(KEYINPUT10), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n333), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n335), .A2(new_n344), .A3(new_n342), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n347), .B1(new_n333), .B2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G120gat), .B(G148gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(G176gat), .B(G204gat), .ZN(new_n351));
  XOR2_X1   g150(.A(new_n350), .B(new_n351), .Z(new_n352));
  OR2_X1    g151(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n349), .A2(new_n352), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n331), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(G78gat), .B(G106gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n357), .B(G22gat), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(G228gat), .A2(G233gat), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(KEYINPUT77), .B(G162gat), .ZN(new_n362));
  INV_X1    g161(.A(G155gat), .ZN(new_n363));
  OAI21_X1  g162(.A(KEYINPUT2), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n323), .A2(G155gat), .ZN(new_n365));
  INV_X1    g164(.A(G141gat), .ZN(new_n366));
  INV_X1    g165(.A(G148gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n363), .A2(G162gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(G141gat), .A2(G148gat), .ZN(new_n370));
  AND4_X1   g169(.A1(new_n365), .A2(new_n368), .A3(new_n369), .A4(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G155gat), .B(G162gat), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT2), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(KEYINPUT76), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT76), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT2), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n368), .A2(new_n375), .A3(new_n377), .A4(new_n370), .ZN(new_n378));
  AOI22_X1  g177(.A1(new_n364), .A2(new_n371), .B1(new_n373), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT22), .ZN(new_n380));
  XNOR2_X1  g179(.A(KEYINPUT73), .B(G218gat), .ZN(new_n381));
  INV_X1    g180(.A(G211gat), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n380), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G211gat), .B(G218gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(G197gat), .B(G204gat), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT74), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n384), .B1(new_n383), .B2(new_n385), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n383), .A2(new_n385), .ZN(new_n391));
  INV_X1    g190(.A(new_n384), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n393), .A2(new_n387), .A3(new_n386), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT29), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n390), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT3), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n379), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n390), .A2(new_n394), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n373), .A2(new_n378), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n323), .A2(KEYINPUT77), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT77), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(G162gat), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n374), .B1(new_n404), .B2(G155gat), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n368), .A2(new_n365), .A3(new_n369), .A4(new_n370), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n400), .B(new_n397), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n395), .ZN(new_n408));
  AND2_X1   g207(.A1(new_n399), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n361), .B1(new_n398), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n399), .A2(new_n408), .ZN(new_n411));
  INV_X1    g210(.A(new_n386), .ZN(new_n412));
  AOI21_X1  g211(.A(KEYINPUT29), .B1(new_n412), .B2(KEYINPUT80), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT80), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n393), .A2(new_n414), .A3(new_n386), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT3), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n411), .B(new_n360), .C1(new_n379), .C2(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(KEYINPUT31), .B(G50gat), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  AND3_X1   g218(.A1(new_n410), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n419), .B1(new_n410), .B2(new_n417), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n359), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n410), .A2(new_n417), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n418), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n410), .A2(new_n417), .A3(new_n419), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n424), .A2(new_n358), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n422), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT36), .ZN(new_n428));
  XNOR2_X1  g227(.A(G15gat), .B(G43gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n429), .B(KEYINPUT71), .ZN(new_n430));
  XNOR2_X1  g229(.A(G71gat), .B(G99gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n430), .B(new_n431), .ZN(new_n432));
  OR2_X1    g231(.A1(new_n432), .A2(KEYINPUT72), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(KEYINPUT72), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n433), .A2(KEYINPUT33), .A3(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT70), .ZN(new_n436));
  NAND2_X1  g235(.A1(G169gat), .A2(G176gat), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT64), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(KEYINPUT64), .A2(G169gat), .A3(G176gat), .ZN(new_n440));
  INV_X1    g239(.A(G169gat), .ZN(new_n441));
  INV_X1    g240(.A(G176gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT23), .ZN(new_n444));
  AOI22_X1  g243(.A1(new_n439), .A2(new_n440), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT24), .ZN(new_n446));
  INV_X1    g245(.A(G183gat), .ZN(new_n447));
  INV_X1    g246(.A(G190gat), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(KEYINPUT24), .B1(new_n448), .B2(G183gat), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n447), .A2(G190gat), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NOR2_X1   g251(.A1(G169gat), .A2(G176gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT23), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n445), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT25), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n453), .A2(KEYINPUT65), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT65), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n459), .B1(G169gat), .B2(G176gat), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n458), .A2(KEYINPUT23), .A3(new_n460), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n445), .A2(new_n452), .A3(new_n461), .A4(KEYINPUT25), .ZN(new_n462));
  XOR2_X1   g261(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n463));
  INV_X1    g262(.A(KEYINPUT27), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(G183gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n447), .A2(KEYINPUT27), .ZN(new_n466));
  AOI21_X1  g265(.A(KEYINPUT66), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(KEYINPUT66), .B1(new_n447), .B2(KEYINPUT27), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(new_n448), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n463), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n465), .A2(new_n466), .A3(KEYINPUT28), .A4(new_n448), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI22_X1  g271(.A1(new_n439), .A2(new_n440), .B1(new_n443), .B2(KEYINPUT26), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT26), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n458), .A2(new_n474), .A3(new_n460), .ZN(new_n475));
  AOI22_X1  g274(.A1(new_n473), .A2(new_n475), .B1(G183gat), .B2(G190gat), .ZN(new_n476));
  AOI22_X1  g275(.A1(new_n457), .A2(new_n462), .B1(new_n472), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT1), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n478), .B1(G113gat), .B2(G120gat), .ZN(new_n479));
  AND2_X1   g278(.A1(G113gat), .A2(G120gat), .ZN(new_n480));
  OAI21_X1  g279(.A(KEYINPUT68), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  XNOR2_X1  g280(.A(G127gat), .B(G134gat), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n482), .B(KEYINPUT68), .C1(new_n480), .C2(new_n479), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n436), .B1(new_n477), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n457), .A2(new_n462), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n476), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n484), .A2(new_n485), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n490), .A2(KEYINPUT70), .A3(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n488), .A2(new_n486), .A3(new_n489), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT69), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT69), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n477), .A2(new_n495), .A3(new_n486), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n487), .A2(new_n492), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(G227gat), .A2(G233gat), .ZN(new_n498));
  OAI211_X1 g297(.A(KEYINPUT32), .B(new_n435), .C1(new_n497), .C2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n487), .A2(new_n492), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n494), .A2(new_n496), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n498), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT32), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n432), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n502), .A2(KEYINPUT33), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n499), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT34), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n507), .B1(new_n497), .B2(new_n498), .ZN(new_n508));
  AND4_X1   g307(.A1(new_n507), .A2(new_n500), .A3(new_n501), .A4(new_n498), .ZN(new_n509));
  OR2_X1    g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n508), .A2(new_n509), .ZN(new_n512));
  OAI21_X1  g311(.A(KEYINPUT32), .B1(new_n497), .B2(new_n498), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT33), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n514), .B1(new_n497), .B2(new_n498), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n513), .A2(new_n515), .A3(new_n432), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n512), .B1(new_n516), .B2(new_n499), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n428), .B1(new_n511), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n506), .A2(new_n510), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n516), .A2(new_n512), .A3(new_n499), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n519), .A2(KEYINPUT36), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n427), .B1(new_n518), .B2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT75), .ZN(new_n523));
  INV_X1    g322(.A(G226gat), .ZN(new_n524));
  INV_X1    g323(.A(G233gat), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n526), .B1(new_n490), .B2(new_n395), .ZN(new_n527));
  INV_X1    g326(.A(new_n399), .ZN(new_n528));
  INV_X1    g327(.A(new_n526), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n477), .A2(new_n529), .ZN(new_n530));
  NOR3_X1   g329(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n529), .B1(new_n477), .B2(KEYINPUT29), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n490), .A2(new_n526), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n399), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n523), .B1(new_n531), .B2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G8gat), .B(G36gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(G64gat), .B(G92gat), .ZN(new_n537));
  XOR2_X1   g336(.A(new_n536), .B(new_n537), .Z(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n528), .B1(new_n527), .B2(new_n530), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n532), .A2(new_n533), .A3(new_n399), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n540), .A2(KEYINPUT75), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n535), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n538), .B1(new_n531), .B2(new_n534), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT30), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n540), .A2(new_n541), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n547), .A2(KEYINPUT30), .A3(new_n538), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n543), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n402), .A2(G162gat), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n323), .A2(KEYINPUT77), .ZN(new_n551));
  OAI21_X1  g350(.A(G155gat), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n406), .B1(new_n552), .B2(KEYINPUT2), .ZN(new_n553));
  AND2_X1   g352(.A1(new_n368), .A2(new_n370), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n375), .A2(new_n377), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n372), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(KEYINPUT3), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n557), .A2(new_n407), .A3(new_n491), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n379), .A2(new_n486), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT4), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n379), .A2(KEYINPUT4), .A3(new_n486), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n558), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(G225gat), .A2(G233gat), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  OR2_X1    g365(.A1(new_n566), .A2(KEYINPUT39), .ZN(new_n567));
  XOR2_X1   g366(.A(G1gat), .B(G29gat), .Z(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT0), .ZN(new_n569));
  XNOR2_X1  g368(.A(G57gat), .B(G85gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n485), .B(new_n484), .C1(new_n553), .C2(new_n556), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n572), .A2(new_n559), .A3(new_n564), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n566), .A2(KEYINPUT39), .A3(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n567), .A2(new_n571), .A3(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT40), .ZN(new_n576));
  OR2_X1    g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT5), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n564), .B1(new_n572), .B2(new_n559), .ZN(new_n579));
  OAI22_X1  g378(.A1(new_n563), .A2(new_n565), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n571), .ZN(new_n581));
  AND3_X1   g380(.A1(new_n379), .A2(KEYINPUT4), .A3(new_n486), .ZN(new_n582));
  AOI21_X1  g381(.A(KEYINPUT4), .B1(new_n379), .B2(new_n486), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n584), .A2(KEYINPUT5), .A3(new_n564), .A4(new_n558), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n580), .A2(new_n581), .A3(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n587), .B1(new_n575), .B2(new_n576), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n549), .A2(new_n577), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n581), .B1(new_n580), .B2(new_n585), .ZN(new_n590));
  AOI21_X1  g389(.A(KEYINPUT6), .B1(new_n590), .B2(KEYINPUT78), .ZN(new_n591));
  AND4_X1   g390(.A1(new_n564), .A2(new_n558), .A3(new_n561), .A4(new_n562), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n579), .A2(new_n578), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n585), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(new_n571), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT78), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n591), .A2(new_n597), .A3(new_n586), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n587), .A2(KEYINPUT6), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT37), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n547), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT38), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n540), .A2(KEYINPUT37), .A3(new_n541), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n601), .A2(new_n602), .A3(new_n539), .A4(new_n603), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n598), .A2(new_n599), .A3(new_n544), .A4(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n535), .A2(KEYINPUT37), .A3(new_n542), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n538), .B1(new_n547), .B2(new_n600), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n602), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n589), .B1(new_n605), .B2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT35), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n549), .B1(new_n599), .B2(new_n598), .ZN(new_n611));
  AND2_X1   g410(.A1(new_n422), .A2(new_n426), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n611), .A2(new_n612), .A3(new_n520), .A4(new_n519), .ZN(new_n613));
  AOI22_X1  g412(.A1(new_n522), .A2(new_n609), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(new_n586), .B(KEYINPUT79), .Z(new_n615));
  NAND2_X1  g414(.A1(new_n591), .A2(new_n597), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n599), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n549), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n612), .B1(new_n518), .B2(new_n521), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n519), .A2(new_n520), .ZN(new_n622));
  NOR3_X1   g421(.A1(new_n622), .A2(new_n610), .A3(new_n427), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n620), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT81), .ZN(new_n625));
  AND3_X1   g424(.A1(new_n614), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n625), .B1(new_n614), .B2(new_n624), .ZN(new_n627));
  OAI211_X1 g426(.A(new_n256), .B(new_n356), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(KEYINPUT91), .ZN(new_n629));
  INV_X1    g428(.A(new_n256), .ZN(new_n630));
  NOR3_X1   g429(.A1(new_n511), .A2(new_n517), .A3(new_n428), .ZN(new_n631));
  AOI21_X1  g430(.A(KEYINPUT36), .B1(new_n519), .B2(new_n520), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n427), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n622), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n634), .A2(KEYINPUT35), .A3(new_n612), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n619), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n609), .B(new_n612), .C1(new_n631), .C2(new_n632), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n613), .A2(new_n610), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(KEYINPUT81), .B1(new_n636), .B2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n614), .A2(new_n624), .A3(new_n625), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n630), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT91), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n642), .A2(new_n643), .A3(new_n356), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n617), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g447(.A1(new_n628), .A2(KEYINPUT91), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n643), .B1(new_n642), .B2(new_n356), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n549), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(KEYINPUT92), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT92), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n645), .A2(new_n653), .A3(new_n549), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g454(.A(KEYINPUT16), .B(G8gat), .Z(new_n656));
  AOI21_X1  g455(.A(KEYINPUT42), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n652), .A2(G8gat), .A3(new_n654), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n645), .A2(KEYINPUT42), .A3(new_n549), .A4(new_n656), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(KEYINPUT93), .B1(new_n657), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n653), .B1(new_n645), .B2(new_n549), .ZN(new_n662));
  AOI211_X1 g461(.A(KEYINPUT92), .B(new_n618), .C1(new_n629), .C2(new_n644), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n656), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT42), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT93), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n666), .A2(new_n667), .A3(new_n658), .A4(new_n659), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n661), .A2(new_n668), .ZN(G1325gat));
  INV_X1    g468(.A(new_n645), .ZN(new_n670));
  OR3_X1    g469(.A1(new_n670), .A2(G15gat), .A3(new_n622), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n518), .A2(new_n521), .ZN(new_n672));
  OAI21_X1  g471(.A(G15gat), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n671), .A2(new_n673), .ZN(G1326gat));
  NAND2_X1  g473(.A1(new_n645), .A2(new_n427), .ZN(new_n675));
  XNOR2_X1  g474(.A(KEYINPUT43), .B(G22gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(G1327gat));
  INV_X1    g476(.A(new_n293), .ZN(new_n678));
  INV_X1    g477(.A(new_n355), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n642), .A2(new_n329), .A3(new_n678), .A4(new_n679), .ZN(new_n680));
  OR2_X1    g479(.A1(new_n617), .A2(G29gat), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n682), .B(KEYINPUT94), .Z(new_n683));
  INV_X1    g482(.A(KEYINPUT45), .ZN(new_n684));
  OR2_X1    g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n330), .B1(new_n640), .B2(new_n641), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687));
  OR3_X1    g486(.A1(new_n686), .A2(KEYINPUT95), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n330), .B1(new_n614), .B2(new_n624), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(new_n687), .ZN(new_n690));
  OAI211_X1 g489(.A(KEYINPUT95), .B(new_n690), .C1(new_n686), .C2(new_n687), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n293), .A2(new_n630), .A3(new_n355), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n688), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(G29gat), .B1(new_n693), .B2(new_n617), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n683), .A2(new_n684), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n685), .A2(new_n694), .A3(new_n695), .ZN(G1328gat));
  OR2_X1    g495(.A1(new_n618), .A2(G36gat), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n680), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT46), .ZN(new_n699));
  OAI21_X1  g498(.A(G36gat), .B1(new_n693), .B2(new_n618), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT96), .ZN(G1329gat));
  INV_X1    g501(.A(new_n672), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(G43gat), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n680), .A2(new_n622), .ZN(new_n705));
  OAI22_X1  g504(.A1(new_n693), .A2(new_n704), .B1(G43gat), .B2(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g506(.A1(new_n680), .A2(G50gat), .A3(new_n612), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n688), .A2(new_n427), .A3(new_n691), .A4(new_n692), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n708), .B1(new_n709), .B2(G50gat), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  XOR2_X1   g510(.A(KEYINPUT97), .B(KEYINPUT48), .Z(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(KEYINPUT98), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT98), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n710), .A2(new_n715), .A3(new_n712), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT99), .ZN(new_n717));
  AND3_X1   g516(.A1(new_n710), .A2(new_n717), .A3(KEYINPUT48), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n717), .B1(new_n710), .B2(KEYINPUT48), .ZN(new_n719));
  OAI22_X1  g518(.A1(new_n714), .A2(new_n716), .B1(new_n718), .B2(new_n719), .ZN(G1331gat));
  AOI21_X1  g519(.A(new_n329), .B1(new_n291), .B2(new_n292), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n721), .A2(new_n630), .A3(new_n355), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n722), .B1(new_n624), .B2(new_n614), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(new_n646), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g524(.A(new_n618), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT100), .ZN(new_n728));
  NOR2_X1   g527(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(G1333gat));
  AOI21_X1  g529(.A(new_n260), .B1(new_n723), .B2(new_n703), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n622), .A2(G71gat), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n731), .B1(new_n723), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g533(.A1(new_n723), .A2(new_n427), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT102), .ZN(new_n736));
  XOR2_X1   g535(.A(KEYINPUT101), .B(G78gat), .Z(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(G1335gat));
  NOR3_X1   g537(.A1(new_n293), .A2(new_n256), .A3(new_n679), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n688), .A2(new_n691), .A3(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(G85gat), .B1(new_n740), .B2(new_n617), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n689), .A2(new_n630), .A3(new_n678), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT51), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n743), .A2(new_n679), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n744), .A2(new_n295), .A3(new_n646), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n741), .A2(new_n745), .ZN(new_n746));
  XOR2_X1   g545(.A(new_n746), .B(KEYINPUT103), .Z(G1336gat));
  NAND4_X1  g546(.A1(new_n688), .A2(new_n549), .A3(new_n691), .A4(new_n739), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(G92gat), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n618), .A2(G92gat), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n744), .A2(new_n750), .ZN(new_n751));
  XOR2_X1   g550(.A(KEYINPUT106), .B(KEYINPUT52), .Z(new_n752));
  NAND3_X1  g551(.A1(new_n749), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  AND3_X1   g552(.A1(new_n748), .A2(KEYINPUT104), .A3(G92gat), .ZN(new_n754));
  AOI21_X1  g553(.A(KEYINPUT104), .B1(new_n748), .B2(G92gat), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n742), .A2(KEYINPUT105), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT51), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n757), .A2(new_n355), .A3(new_n750), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n754), .A2(new_n755), .A3(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT52), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n753), .B1(new_n759), .B2(new_n760), .ZN(G1337gat));
  OAI21_X1  g560(.A(G99gat), .B1(new_n740), .B2(new_n672), .ZN(new_n762));
  INV_X1    g561(.A(G99gat), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n744), .A2(new_n763), .A3(new_n634), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n762), .A2(new_n764), .ZN(G1338gat));
  XOR2_X1   g564(.A(KEYINPUT107), .B(KEYINPUT53), .Z(new_n766));
  NOR2_X1   g565(.A1(new_n612), .A2(G106gat), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n766), .B1(new_n744), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(G106gat), .B1(new_n740), .B2(new_n612), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n757), .A2(new_n355), .A3(new_n767), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT53), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n770), .B1(new_n772), .B2(new_n773), .ZN(G1339gat));
  NAND3_X1  g573(.A1(new_n721), .A2(new_n630), .A3(new_n679), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n345), .A2(new_n346), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(new_n332), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n345), .A2(new_n333), .A3(new_n346), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n777), .A2(KEYINPUT54), .A3(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT54), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n352), .B1(new_n347), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n779), .A2(KEYINPUT55), .A3(new_n781), .ZN(new_n782));
  AND3_X1   g581(.A1(new_n329), .A2(new_n782), .A3(new_n354), .ZN(new_n783));
  AND3_X1   g582(.A1(new_n230), .A2(new_n232), .A3(new_n204), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n202), .B1(new_n245), .B2(new_n232), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n239), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n250), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT108), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n779), .A2(new_n781), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT55), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  AOI211_X1 g590(.A(KEYINPUT108), .B(KEYINPUT55), .C1(new_n779), .C2(new_n781), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n783), .B(new_n787), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT109), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OR2_X1    g594(.A1(new_n791), .A2(new_n792), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n796), .A2(KEYINPUT109), .A3(new_n787), .A4(new_n783), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n787), .A2(new_n355), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n791), .A2(new_n792), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n256), .A2(new_n354), .A3(new_n782), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  AOI22_X1  g600(.A1(new_n795), .A2(new_n797), .B1(new_n801), .B2(new_n330), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n775), .B1(new_n802), .B2(new_n293), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n804), .A2(new_n427), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n622), .A2(new_n617), .A3(new_n549), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(G113gat), .B1(new_n807), .B2(new_n630), .ZN(new_n808));
  XOR2_X1   g607(.A(new_n808), .B(KEYINPUT110), .Z(new_n809));
  NAND2_X1  g608(.A1(new_n803), .A2(new_n646), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n634), .A2(new_n612), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n810), .A2(new_n811), .A3(new_n549), .ZN(new_n812));
  INV_X1    g611(.A(G113gat), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n812), .A2(new_n813), .A3(new_n256), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n809), .A2(new_n814), .ZN(G1340gat));
  INV_X1    g614(.A(G120gat), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n807), .A2(new_n816), .A3(new_n679), .ZN(new_n817));
  AOI21_X1  g616(.A(G120gat), .B1(new_n812), .B2(new_n355), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n817), .A2(new_n818), .ZN(G1341gat));
  OAI21_X1  g618(.A(G127gat), .B1(new_n807), .B2(new_n678), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n812), .A2(new_n283), .A3(new_n293), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(G1342gat));
  NAND2_X1  g621(.A1(new_n618), .A2(new_n329), .ZN(new_n823));
  XOR2_X1   g622(.A(new_n823), .B(KEYINPUT111), .Z(new_n824));
  OR4_X1    g623(.A1(G134gat), .A2(new_n810), .A3(new_n811), .A4(new_n824), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n825), .A2(KEYINPUT56), .ZN(new_n826));
  XOR2_X1   g625(.A(new_n826), .B(KEYINPUT112), .Z(new_n827));
  NAND3_X1  g626(.A1(new_n805), .A2(new_n329), .A3(new_n806), .ZN(new_n828));
  AOI22_X1  g627(.A1(new_n825), .A2(KEYINPUT56), .B1(G134gat), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n829), .ZN(G1343gat));
  NAND3_X1  g629(.A1(new_n672), .A2(new_n646), .A3(new_n618), .ZN(new_n831));
  XOR2_X1   g630(.A(new_n831), .B(KEYINPUT113), .Z(new_n832));
  INV_X1    g631(.A(KEYINPUT57), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n612), .A2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(new_n775), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n795), .A2(new_n797), .ZN(new_n837));
  AOI21_X1  g636(.A(KEYINPUT55), .B1(new_n779), .B2(new_n781), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT114), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n838), .B(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n798), .B1(new_n840), .B2(new_n800), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n330), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n293), .B1(new_n837), .B2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT115), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n836), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AOI22_X1  g644(.A1(new_n795), .A2(new_n797), .B1(new_n841), .B2(new_n330), .ZN(new_n846));
  OAI21_X1  g645(.A(KEYINPUT115), .B1(new_n846), .B2(new_n293), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n835), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(KEYINPUT57), .B1(new_n803), .B2(new_n427), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n256), .B(new_n832), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT117), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n837), .A2(new_n842), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n853), .A2(new_n844), .A3(new_n678), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n854), .A2(new_n847), .A3(new_n775), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n834), .ZN(new_n856));
  INV_X1    g655(.A(new_n849), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n858), .A2(KEYINPUT117), .A3(new_n256), .A4(new_n832), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n852), .A2(new_n859), .A3(G141gat), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT58), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT116), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n633), .B1(new_n810), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n803), .A2(KEYINPUT116), .A3(new_n646), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n863), .A2(new_n618), .A3(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n630), .A2(G141gat), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n861), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n860), .A2(new_n869), .ZN(new_n870));
  AND3_X1   g669(.A1(new_n863), .A2(new_n618), .A3(new_n864), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n866), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n850), .A2(G141gat), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(KEYINPUT58), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT118), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n870), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n366), .B1(new_n850), .B2(new_n851), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n868), .B1(new_n878), .B2(new_n859), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n861), .B1(new_n872), .B2(new_n873), .ZN(new_n880));
  OAI21_X1  g679(.A(KEYINPUT118), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n877), .A2(new_n881), .ZN(G1344gat));
  NAND3_X1  g681(.A1(new_n871), .A2(new_n367), .A3(new_n355), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n858), .A2(new_n832), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n884), .A2(new_n679), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n885), .A2(KEYINPUT59), .A3(new_n367), .ZN(new_n886));
  XOR2_X1   g685(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n887));
  NAND3_X1  g686(.A1(new_n796), .A2(KEYINPUT120), .A3(new_n783), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n787), .ZN(new_n889));
  AOI21_X1  g688(.A(KEYINPUT120), .B1(new_n796), .B2(new_n783), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n842), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n836), .B1(new_n891), .B2(new_n678), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n892), .A2(KEYINPUT57), .A3(new_n612), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n833), .B1(new_n803), .B2(new_n427), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n832), .A2(new_n355), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT121), .ZN(new_n897));
  OR2_X1    g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n367), .B1(new_n896), .B2(new_n897), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n887), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n883), .B1(new_n886), .B2(new_n900), .ZN(G1345gat));
  OAI21_X1  g700(.A(G155gat), .B1(new_n884), .B2(new_n678), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n871), .A2(new_n363), .A3(new_n293), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(G1346gat));
  OAI21_X1  g703(.A(new_n404), .B1(new_n884), .B2(new_n330), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n824), .A2(new_n404), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n863), .A2(new_n864), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT122), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n908), .B(new_n909), .ZN(G1347gat));
  NAND2_X1  g709(.A1(new_n617), .A2(new_n549), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n911), .A2(new_n622), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n805), .A2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT123), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n805), .A2(KEYINPUT123), .A3(new_n912), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n917), .A2(new_n441), .A3(new_n630), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n804), .A2(new_n646), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n811), .A2(new_n618), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(G169gat), .B1(new_n922), .B2(new_n256), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n918), .A2(new_n923), .ZN(G1348gat));
  OAI21_X1  g723(.A(G176gat), .B1(new_n917), .B2(new_n679), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n922), .A2(new_n442), .A3(new_n355), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(G1349gat));
  NAND3_X1  g726(.A1(new_n293), .A2(new_n465), .A3(new_n466), .ZN(new_n928));
  OR3_X1    g727(.A1(new_n921), .A2(KEYINPUT124), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g728(.A(KEYINPUT124), .B1(new_n921), .B2(new_n928), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n917), .A2(new_n678), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n931), .B1(new_n932), .B2(new_n447), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(KEYINPUT60), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT60), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n935), .B(new_n931), .C1(new_n932), .C2(new_n447), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n936), .ZN(G1350gat));
  NAND3_X1  g736(.A1(new_n922), .A2(new_n448), .A3(new_n329), .ZN(new_n938));
  OAI21_X1  g737(.A(G190gat), .B1(new_n917), .B2(new_n330), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n939), .A2(KEYINPUT61), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n939), .A2(KEYINPUT61), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n938), .B1(new_n940), .B2(new_n941), .ZN(G1351gat));
  NOR2_X1   g741(.A1(new_n893), .A2(new_n894), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n703), .A2(new_n911), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(G197gat), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n945), .A2(new_n946), .A3(new_n630), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n633), .A2(new_n618), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n919), .A2(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(G197gat), .B1(new_n950), .B2(new_n256), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n947), .A2(new_n951), .ZN(G1352gat));
  NOR3_X1   g751(.A1(new_n949), .A2(G204gat), .A3(new_n679), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(KEYINPUT62), .ZN(new_n954));
  OAI21_X1  g753(.A(G204gat), .B1(new_n945), .B2(new_n679), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(G1353gat));
  NAND3_X1  g755(.A1(new_n950), .A2(new_n382), .A3(new_n293), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n943), .A2(new_n293), .A3(new_n944), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n958), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n959));
  AOI21_X1  g758(.A(KEYINPUT63), .B1(new_n958), .B2(G211gat), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n957), .B1(new_n959), .B2(new_n960), .ZN(G1354gat));
  INV_X1    g760(.A(G218gat), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n962), .B1(new_n949), .B2(new_n330), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n963), .A2(KEYINPUT125), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n963), .A2(KEYINPUT125), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n330), .A2(new_n381), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n966), .B(KEYINPUT126), .ZN(new_n967));
  INV_X1    g766(.A(new_n967), .ZN(new_n968));
  OAI22_X1  g767(.A1(new_n964), .A2(new_n965), .B1(new_n945), .B2(new_n968), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT127), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OAI221_X1 g770(.A(KEYINPUT127), .B1(new_n945), .B2(new_n968), .C1(new_n964), .C2(new_n965), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(G1355gat));
endmodule


