

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730;

  AND2_X1 U366 ( .A1(n594), .A2(n591), .ZN(n345) );
  NOR2_X1 U367 ( .A1(n728), .A2(n730), .ZN(n563) );
  NAND2_X1 U368 ( .A1(n580), .A2(n661), .ZN(n369) );
  AND2_X1 U369 ( .A1(n347), .A2(n552), .ZN(n580) );
  NAND2_X1 U370 ( .A1(n344), .A2(n343), .ZN(n547) );
  INV_X1 U371 ( .A(n545), .ZN(n344) );
  INV_X1 U372 ( .A(n492), .ZN(n671) );
  INV_X1 U373 ( .A(n544), .ZN(n343) );
  BUF_X1 U374 ( .A(n490), .Z(n676) );
  BUF_X1 U375 ( .A(G116), .Z(n346) );
  XNOR2_X1 U376 ( .A(n719), .B(G146), .ZN(n464) );
  INV_X1 U377 ( .A(G125), .ZN(n379) );
  XNOR2_X1 U378 ( .A(KEYINPUT3), .B(G116), .ZN(n386) );
  XNOR2_X2 U379 ( .A(n468), .B(n467), .ZN(n545) );
  NAND2_X1 U380 ( .A1(n592), .A2(n345), .ZN(n596) );
  INV_X2 U381 ( .A(n704), .ZN(n371) );
  AND2_X1 U382 ( .A1(n550), .A2(n549), .ZN(n347) );
  XNOR2_X1 U383 ( .A(n463), .B(n464), .ZN(n600) );
  NOR2_X1 U384 ( .A1(n642), .A2(n665), .ZN(n574) );
  NOR2_X1 U385 ( .A1(n548), .A2(n676), .ZN(n475) );
  INV_X1 U386 ( .A(G953), .ZN(n720) );
  XNOR2_X1 U387 ( .A(n488), .B(KEYINPUT32), .ZN(n510) );
  OR2_X2 U388 ( .A1(n558), .A2(n513), .ZN(n571) );
  XNOR2_X2 U389 ( .A(n441), .B(n440), .ZN(n513) );
  XNOR2_X2 U390 ( .A(n370), .B(n348), .ZN(n490) );
  NOR2_X2 U391 ( .A1(n502), .A2(n501), .ZN(n503) );
  NOR2_X1 U392 ( .A1(n359), .A2(n356), .ZN(n355) );
  AND2_X1 U393 ( .A1(n510), .A2(n608), .ZN(n373) );
  XNOR2_X1 U394 ( .A(n509), .B(n508), .ZN(n608) );
  XNOR2_X1 U395 ( .A(n496), .B(n495), .ZN(n518) );
  OR2_X1 U396 ( .A1(n682), .A2(n515), .ZN(n496) );
  XNOR2_X1 U397 ( .A(n464), .B(n365), .ZN(n701) );
  INV_X2 U398 ( .A(G143), .ZN(n383) );
  NOR2_X1 U399 ( .A1(n360), .A2(n362), .ZN(n359) );
  NAND2_X1 U400 ( .A1(n358), .A2(KEYINPUT65), .ZN(n357) );
  INV_X1 U401 ( .A(n350), .ZN(n358) );
  BUF_X1 U402 ( .A(n543), .Z(n597) );
  XNOR2_X1 U403 ( .A(KEYINPUT103), .B(KEYINPUT30), .ZN(n546) );
  XNOR2_X1 U404 ( .A(n395), .B(n394), .ZN(n481) );
  OR2_X1 U405 ( .A1(n620), .A2(n542), .ZN(n395) );
  NOR2_X1 U406 ( .A1(n513), .A2(n672), .ZN(n514) );
  AND2_X1 U407 ( .A1(n350), .A2(n362), .ZN(n354) );
  OR2_X2 U408 ( .A1(n481), .A2(n544), .ZN(n565) );
  NAND2_X1 U409 ( .A1(n490), .A2(n677), .ZN(n672) );
  XOR2_X1 U410 ( .A(KEYINPUT75), .B(G119), .Z(n460) );
  XNOR2_X1 U411 ( .A(G137), .B(G113), .ZN(n459) );
  XNOR2_X1 U412 ( .A(n438), .B(n376), .ZN(n719) );
  XNOR2_X1 U413 ( .A(n352), .B(n351), .ZN(n364) );
  INV_X1 U414 ( .A(n652), .ZN(n363) );
  INV_X1 U415 ( .A(KEYINPUT78), .ZN(n351) );
  XNOR2_X1 U416 ( .A(G101), .B(G104), .ZN(n439) );
  XNOR2_X1 U417 ( .A(n367), .B(n366), .ZN(n365) );
  XNOR2_X1 U418 ( .A(n349), .B(n439), .ZN(n366) );
  XNOR2_X1 U419 ( .A(n377), .B(n448), .ZN(n367) );
  NAND2_X1 U420 ( .A1(n598), .A2(n597), .ZN(n656) );
  INV_X1 U421 ( .A(n548), .ZN(n549) );
  XNOR2_X1 U422 ( .A(n547), .B(n546), .ZN(n550) );
  BUF_X1 U423 ( .A(n481), .Z(n577) );
  INV_X1 U424 ( .A(KEYINPUT28), .ZN(n556) );
  BUF_X1 U425 ( .A(n500), .Z(n484) );
  AND2_X1 U426 ( .A1(n603), .A2(G953), .ZN(n715) );
  XNOR2_X1 U427 ( .A(n567), .B(KEYINPUT36), .ZN(n568) );
  NAND2_X1 U428 ( .A1(n374), .A2(n375), .ZN(n511) );
  XNOR2_X1 U429 ( .A(n498), .B(KEYINPUT101), .ZN(n374) );
  XOR2_X1 U430 ( .A(n452), .B(KEYINPUT25), .Z(n348) );
  XNOR2_X1 U431 ( .A(n531), .B(n530), .ZN(n543) );
  AND2_X1 U432 ( .A1(G227), .A2(n720), .ZN(n349) );
  OR2_X1 U433 ( .A1(n590), .A2(n654), .ZN(n350) );
  INV_X1 U434 ( .A(KEYINPUT65), .ZN(n362) );
  NAND2_X1 U435 ( .A1(n543), .A2(n542), .ZN(n352) );
  NAND2_X1 U436 ( .A1(n355), .A2(n353), .ZN(n704) );
  NAND2_X1 U437 ( .A1(n360), .A2(n354), .ZN(n353) );
  NAND2_X1 U438 ( .A1(n656), .A2(n357), .ZN(n356) );
  NAND2_X1 U439 ( .A1(n364), .A2(n363), .ZN(n360) );
  XNOR2_X2 U440 ( .A(n361), .B(n384), .ZN(n438) );
  XNOR2_X1 U441 ( .A(n361), .B(n346), .ZN(n428) );
  XNOR2_X2 U442 ( .A(n383), .B(G128), .ZN(n361) );
  XNOR2_X1 U443 ( .A(n443), .B(n421), .ZN(n390) );
  XNOR2_X2 U444 ( .A(G122), .B(G107), .ZN(n421) );
  XNOR2_X2 U445 ( .A(G119), .B(G110), .ZN(n443) );
  NAND2_X1 U446 ( .A1(n572), .A2(n402), .ZN(n403) );
  XNOR2_X2 U447 ( .A(n565), .B(KEYINPUT19), .ZN(n572) );
  NAND2_X1 U448 ( .A1(n368), .A2(n487), .ZN(n488) );
  NAND2_X1 U449 ( .A1(n368), .A2(n673), .ZN(n498) );
  NAND2_X1 U450 ( .A1(n368), .A2(n470), .ZN(n524) );
  XNOR2_X2 U451 ( .A(n437), .B(n436), .ZN(n368) );
  NAND2_X1 U452 ( .A1(n587), .A2(n626), .ZN(n554) );
  XNOR2_X2 U453 ( .A(n369), .B(KEYINPUT39), .ZN(n587) );
  OR2_X2 U454 ( .A1(n712), .A2(G902), .ZN(n370) );
  NAND2_X1 U455 ( .A1(n371), .A2(G475), .ZN(n614) );
  NAND2_X1 U456 ( .A1(n371), .A2(G210), .ZN(n622) );
  XNOR2_X1 U457 ( .A(n372), .B(n512), .ZN(n529) );
  NAND2_X1 U458 ( .A1(n373), .A2(n511), .ZN(n372) );
  XNOR2_X2 U459 ( .A(G113), .B(G104), .ZN(n412) );
  AND2_X1 U460 ( .A1(n671), .A2(n499), .ZN(n375) );
  XOR2_X1 U461 ( .A(G131), .B(G134), .Z(n376) );
  XOR2_X1 U462 ( .A(G110), .B(G107), .Z(n377) );
  INV_X1 U463 ( .A(KEYINPUT47), .ZN(n575) );
  XNOR2_X1 U464 ( .A(n576), .B(n575), .ZN(n581) );
  XNOR2_X1 U465 ( .A(G469), .B(KEYINPUT70), .ZN(n440) );
  BUF_X1 U466 ( .A(n659), .Z(n693) );
  INV_X1 U467 ( .A(KEYINPUT106), .ZN(n567) );
  XNOR2_X1 U468 ( .A(n545), .B(KEYINPUT6), .ZN(n500) );
  XNOR2_X1 U469 ( .A(n569), .B(n568), .ZN(n570) );
  BUF_X1 U470 ( .A(n518), .Z(n646) );
  NAND2_X1 U471 ( .A1(n720), .A2(G224), .ZN(n378) );
  XNOR2_X1 U472 ( .A(n378), .B(KEYINPUT85), .ZN(n382) );
  XNOR2_X2 U473 ( .A(n379), .B(G146), .ZN(n404) );
  XNOR2_X1 U474 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n380) );
  XNOR2_X1 U475 ( .A(n404), .B(n380), .ZN(n381) );
  XNOR2_X1 U476 ( .A(n382), .B(n381), .ZN(n385) );
  INV_X1 U477 ( .A(KEYINPUT4), .ZN(n384) );
  XNOR2_X1 U478 ( .A(n385), .B(n438), .ZN(n392) );
  XNOR2_X1 U479 ( .A(n386), .B(KEYINPUT72), .ZN(n388) );
  XOR2_X1 U480 ( .A(G101), .B(KEYINPUT71), .Z(n387) );
  XNOR2_X1 U481 ( .A(n388), .B(n387), .ZN(n453) );
  XNOR2_X1 U482 ( .A(n412), .B(KEYINPUT16), .ZN(n389) );
  XNOR2_X1 U483 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U484 ( .A(n453), .B(n391), .ZN(n537) );
  XNOR2_X1 U485 ( .A(n392), .B(n537), .ZN(n620) );
  XNOR2_X1 U486 ( .A(G902), .B(KEYINPUT15), .ZN(n590) );
  INV_X1 U487 ( .A(n590), .ZN(n542) );
  INV_X1 U488 ( .A(G902), .ZN(n465) );
  INV_X1 U489 ( .A(G237), .ZN(n393) );
  NAND2_X1 U490 ( .A1(n465), .A2(n393), .ZN(n396) );
  NAND2_X1 U491 ( .A1(n396), .A2(G210), .ZN(n394) );
  NAND2_X1 U492 ( .A1(n396), .A2(G214), .ZN(n660) );
  INV_X1 U493 ( .A(n660), .ZN(n544) );
  NAND2_X1 U494 ( .A1(G234), .A2(G237), .ZN(n397) );
  XNOR2_X1 U495 ( .A(n397), .B(KEYINPUT14), .ZN(n399) );
  NAND2_X1 U496 ( .A1(n399), .A2(G902), .ZN(n398) );
  XOR2_X1 U497 ( .A(KEYINPUT87), .B(n398), .Z(n471) );
  XOR2_X1 U498 ( .A(G898), .B(KEYINPUT86), .Z(n534) );
  NAND2_X1 U499 ( .A1(G953), .A2(n534), .ZN(n538) );
  OR2_X1 U500 ( .A1(n471), .A2(n538), .ZN(n401) );
  NAND2_X1 U501 ( .A1(G952), .A2(n399), .ZN(n692) );
  NOR2_X1 U502 ( .A1(n692), .A2(G953), .ZN(n474) );
  INV_X1 U503 ( .A(n474), .ZN(n400) );
  NAND2_X1 U504 ( .A1(n401), .A2(n400), .ZN(n402) );
  XNOR2_X2 U505 ( .A(n403), .B(KEYINPUT0), .ZN(n515) );
  XOR2_X1 U506 ( .A(KEYINPUT10), .B(n404), .Z(n449) );
  XOR2_X1 U507 ( .A(KEYINPUT11), .B(KEYINPUT95), .Z(n406) );
  XNOR2_X1 U508 ( .A(G131), .B(KEYINPUT97), .ZN(n405) );
  XNOR2_X1 U509 ( .A(n406), .B(n405), .ZN(n408) );
  XOR2_X1 U510 ( .A(G122), .B(G140), .Z(n407) );
  XNOR2_X1 U511 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U512 ( .A(n449), .B(n409), .ZN(n416) );
  NOR2_X1 U513 ( .A1(G953), .A2(G237), .ZN(n454) );
  NAND2_X1 U514 ( .A1(G214), .A2(n454), .ZN(n410) );
  XNOR2_X1 U515 ( .A(n410), .B(KEYINPUT96), .ZN(n414) );
  XNOR2_X1 U516 ( .A(G143), .B(KEYINPUT12), .ZN(n411) );
  XNOR2_X1 U517 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U518 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U519 ( .A(n416), .B(n415), .ZN(n612) );
  NAND2_X1 U520 ( .A1(n612), .A2(n465), .ZN(n418) );
  XNOR2_X1 U521 ( .A(KEYINPUT13), .B(G475), .ZN(n417) );
  XNOR2_X1 U522 ( .A(n418), .B(n417), .ZN(n521) );
  NAND2_X1 U523 ( .A1(n720), .A2(G234), .ZN(n420) );
  XNOR2_X1 U524 ( .A(KEYINPUT8), .B(KEYINPUT69), .ZN(n419) );
  XNOR2_X1 U525 ( .A(n420), .B(n419), .ZN(n442) );
  NAND2_X1 U526 ( .A1(n442), .A2(G217), .ZN(n426) );
  XNOR2_X1 U527 ( .A(KEYINPUT98), .B(KEYINPUT7), .ZN(n422) );
  XNOR2_X1 U528 ( .A(n422), .B(n421), .ZN(n424) );
  XNOR2_X1 U529 ( .A(G134), .B(KEYINPUT9), .ZN(n423) );
  XOR2_X1 U530 ( .A(n424), .B(n423), .Z(n425) );
  XNOR2_X1 U531 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U532 ( .A(n428), .B(n427), .ZN(n708) );
  NOR2_X1 U533 ( .A1(G902), .A2(n708), .ZN(n429) );
  XNOR2_X1 U534 ( .A(G478), .B(n429), .ZN(n505) );
  NAND2_X1 U535 ( .A1(n521), .A2(n505), .ZN(n430) );
  XNOR2_X1 U536 ( .A(n430), .B(KEYINPUT99), .ZN(n559) );
  NAND2_X1 U537 ( .A1(n590), .A2(G234), .ZN(n431) );
  XNOR2_X1 U538 ( .A(n431), .B(KEYINPUT20), .ZN(n451) );
  NAND2_X1 U539 ( .A1(n451), .A2(G221), .ZN(n433) );
  XOR2_X1 U540 ( .A(KEYINPUT88), .B(KEYINPUT21), .Z(n432) );
  XNOR2_X1 U541 ( .A(n433), .B(n432), .ZN(n677) );
  NAND2_X1 U542 ( .A1(n559), .A2(n677), .ZN(n434) );
  OR2_X2 U543 ( .A1(n515), .A2(n434), .ZN(n437) );
  INV_X1 U544 ( .A(KEYINPUT74), .ZN(n435) );
  XNOR2_X1 U545 ( .A(n435), .B(KEYINPUT22), .ZN(n436) );
  XNOR2_X1 U546 ( .A(G137), .B(G140), .ZN(n448) );
  NOR2_X1 U547 ( .A1(n701), .A2(G902), .ZN(n441) );
  XNOR2_X1 U548 ( .A(n513), .B(KEYINPUT1), .ZN(n491) );
  BUF_X1 U549 ( .A(n491), .Z(n673) );
  NAND2_X1 U550 ( .A1(n442), .A2(G221), .ZN(n447) );
  XOR2_X1 U551 ( .A(G128), .B(n443), .Z(n445) );
  XOR2_X1 U552 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n444) );
  XNOR2_X1 U553 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U554 ( .A(n447), .B(n446), .ZN(n450) );
  XNOR2_X1 U555 ( .A(n449), .B(n448), .ZN(n716) );
  XNOR2_X1 U556 ( .A(n450), .B(n716), .ZN(n712) );
  NAND2_X1 U557 ( .A1(n451), .A2(G217), .ZN(n452) );
  NAND2_X1 U558 ( .A1(n673), .A2(n676), .ZN(n469) );
  INV_X1 U559 ( .A(n453), .ZN(n458) );
  XOR2_X1 U560 ( .A(KEYINPUT5), .B(KEYINPUT90), .Z(n456) );
  NAND2_X1 U561 ( .A1(G210), .A2(n454), .ZN(n455) );
  XNOR2_X1 U562 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U563 ( .A(n458), .B(n457), .ZN(n462) );
  XNOR2_X1 U564 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U565 ( .A(n462), .B(n461), .ZN(n463) );
  NAND2_X1 U566 ( .A1(n600), .A2(n465), .ZN(n468) );
  XNOR2_X1 U567 ( .A(KEYINPUT73), .B(KEYINPUT91), .ZN(n466) );
  INV_X1 U568 ( .A(G472), .ZN(n599) );
  XNOR2_X1 U569 ( .A(n466), .B(n599), .ZN(n467) );
  NOR2_X1 U570 ( .A1(n469), .A2(n484), .ZN(n470) );
  XNOR2_X1 U571 ( .A(n524), .B(G101), .ZN(G3) );
  INV_X1 U572 ( .A(n673), .ZN(n477) );
  INV_X1 U573 ( .A(n505), .ZN(n520) );
  OR2_X1 U574 ( .A1(n521), .A2(n520), .ZN(n641) );
  OR2_X1 U575 ( .A1(n720), .A2(n471), .ZN(n472) );
  NOR2_X1 U576 ( .A1(G900), .A2(n472), .ZN(n473) );
  NOR2_X1 U577 ( .A1(n474), .A2(n473), .ZN(n548) );
  NAND2_X1 U578 ( .A1(n677), .A2(n475), .ZN(n555) );
  NOR2_X1 U579 ( .A1(n641), .A2(n555), .ZN(n476) );
  NAND2_X1 U580 ( .A1(n484), .A2(n476), .ZN(n564) );
  NOR2_X1 U581 ( .A1(n477), .A2(n564), .ZN(n478) );
  NAND2_X1 U582 ( .A1(n478), .A2(n660), .ZN(n480) );
  XNOR2_X1 U583 ( .A(KEYINPUT102), .B(KEYINPUT43), .ZN(n479) );
  XNOR2_X1 U584 ( .A(n480), .B(n479), .ZN(n482) );
  NAND2_X1 U585 ( .A1(n482), .A2(n577), .ZN(n591) );
  XOR2_X1 U586 ( .A(G140), .B(KEYINPUT115), .Z(n483) );
  XNOR2_X1 U587 ( .A(n591), .B(n483), .ZN(G42) );
  OR2_X1 U588 ( .A1(n673), .A2(n676), .ZN(n485) );
  NOR2_X1 U589 ( .A1(n485), .A2(n484), .ZN(n486) );
  XNOR2_X1 U590 ( .A(n486), .B(KEYINPUT76), .ZN(n487) );
  XOR2_X1 U591 ( .A(G119), .B(KEYINPUT127), .Z(n489) );
  XNOR2_X1 U592 ( .A(n510), .B(n489), .ZN(G21) );
  OR2_X2 U593 ( .A1(n491), .A2(n672), .ZN(n501) );
  INV_X1 U594 ( .A(n545), .ZN(n492) );
  NOR2_X1 U595 ( .A1(n501), .A2(n671), .ZN(n494) );
  INV_X1 U596 ( .A(KEYINPUT92), .ZN(n493) );
  XNOR2_X1 U597 ( .A(n494), .B(n493), .ZN(n682) );
  XNOR2_X1 U598 ( .A(KEYINPUT93), .B(KEYINPUT31), .ZN(n495) );
  NOR2_X1 U599 ( .A1(n646), .A2(n641), .ZN(n497) );
  XOR2_X1 U600 ( .A(G113), .B(n497), .Z(G15) );
  INV_X1 U601 ( .A(n676), .ZN(n499) );
  XNOR2_X1 U602 ( .A(n511), .B(G110), .ZN(G12) );
  INV_X1 U603 ( .A(n500), .ZN(n502) );
  XNOR2_X1 U604 ( .A(n503), .B(KEYINPUT33), .ZN(n659) );
  NOR2_X1 U605 ( .A1(n659), .A2(n515), .ZN(n504) );
  XNOR2_X1 U606 ( .A(n504), .B(KEYINPUT34), .ZN(n507) );
  OR2_X1 U607 ( .A1(n521), .A2(n505), .ZN(n578) );
  INV_X1 U608 ( .A(n578), .ZN(n506) );
  NAND2_X1 U609 ( .A1(n507), .A2(n506), .ZN(n509) );
  INV_X1 U610 ( .A(KEYINPUT35), .ZN(n508) );
  INV_X1 U611 ( .A(KEYINPUT44), .ZN(n512) );
  XOR2_X1 U612 ( .A(KEYINPUT89), .B(n514), .Z(n552) );
  AND2_X1 U613 ( .A1(n552), .A2(n671), .ZN(n517) );
  INV_X1 U614 ( .A(n515), .ZN(n516) );
  NAND2_X1 U615 ( .A1(n517), .A2(n516), .ZN(n625) );
  NAND2_X1 U616 ( .A1(n518), .A2(n625), .ZN(n519) );
  XNOR2_X1 U617 ( .A(n519), .B(KEYINPUT94), .ZN(n523) );
  NAND2_X1 U618 ( .A1(n521), .A2(n520), .ZN(n645) );
  AND2_X1 U619 ( .A1(n641), .A2(n645), .ZN(n665) );
  INV_X1 U620 ( .A(n665), .ZN(n522) );
  NAND2_X1 U621 ( .A1(n523), .A2(n522), .ZN(n525) );
  NAND2_X1 U622 ( .A1(n525), .A2(n524), .ZN(n527) );
  INV_X1 U623 ( .A(KEYINPUT100), .ZN(n526) );
  XNOR2_X1 U624 ( .A(n527), .B(n526), .ZN(n528) );
  NAND2_X1 U625 ( .A1(n529), .A2(n528), .ZN(n531) );
  XNOR2_X1 U626 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n530) );
  INV_X1 U627 ( .A(n597), .ZN(n653) );
  NOR2_X1 U628 ( .A1(n653), .A2(G953), .ZN(n536) );
  NAND2_X1 U629 ( .A1(G953), .A2(G224), .ZN(n532) );
  XOR2_X1 U630 ( .A(KEYINPUT61), .B(n532), .Z(n533) );
  NOR2_X1 U631 ( .A1(n534), .A2(n533), .ZN(n535) );
  NOR2_X1 U632 ( .A1(n536), .A2(n535), .ZN(n541) );
  INV_X1 U633 ( .A(n537), .ZN(n539) );
  NAND2_X1 U634 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U635 ( .A(n541), .B(n540), .ZN(G69) );
  INV_X1 U636 ( .A(n641), .ZN(n626) );
  XNOR2_X1 U637 ( .A(n577), .B(KEYINPUT38), .ZN(n661) );
  XOR2_X1 U638 ( .A(KEYINPUT40), .B(KEYINPUT104), .Z(n553) );
  XNOR2_X1 U639 ( .A(n554), .B(n553), .ZN(n728) );
  NOR2_X1 U640 ( .A1(n555), .A2(n671), .ZN(n557) );
  XNOR2_X1 U641 ( .A(n557), .B(n556), .ZN(n558) );
  NAND2_X1 U642 ( .A1(n661), .A2(n660), .ZN(n664) );
  INV_X1 U643 ( .A(n559), .ZN(n663) );
  NOR2_X1 U644 ( .A1(n664), .A2(n663), .ZN(n560) );
  XNOR2_X1 U645 ( .A(n560), .B(KEYINPUT41), .ZN(n694) );
  NOR2_X1 U646 ( .A1(n571), .A2(n694), .ZN(n561) );
  XNOR2_X1 U647 ( .A(n561), .B(KEYINPUT42), .ZN(n730) );
  XNOR2_X1 U648 ( .A(KEYINPUT46), .B(KEYINPUT82), .ZN(n562) );
  XNOR2_X1 U649 ( .A(n563), .B(n562), .ZN(n584) );
  XOR2_X1 U650 ( .A(n564), .B(KEYINPUT105), .Z(n566) );
  NOR2_X1 U651 ( .A1(n566), .A2(n565), .ZN(n569) );
  NOR2_X1 U652 ( .A1(n673), .A2(n570), .ZN(n649) );
  INV_X1 U653 ( .A(n571), .ZN(n573) );
  NAND2_X1 U654 ( .A1(n573), .A2(n572), .ZN(n642) );
  NAND2_X1 U655 ( .A1(KEYINPUT68), .A2(n574), .ZN(n576) );
  NOR2_X1 U656 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U657 ( .A1(n580), .A2(n579), .ZN(n639) );
  NAND2_X1 U658 ( .A1(n581), .A2(n639), .ZN(n582) );
  NOR2_X1 U659 ( .A1(n649), .A2(n582), .ZN(n583) );
  NAND2_X1 U660 ( .A1(n584), .A2(n583), .ZN(n586) );
  INV_X1 U661 ( .A(KEYINPUT48), .ZN(n585) );
  XNOR2_X1 U662 ( .A(n586), .B(n585), .ZN(n592) );
  INV_X1 U663 ( .A(n645), .ZN(n631) );
  NAND2_X1 U664 ( .A1(n587), .A2(n631), .ZN(n651) );
  AND2_X1 U665 ( .A1(n591), .A2(n651), .ZN(n588) );
  NAND2_X1 U666 ( .A1(n592), .A2(n588), .ZN(n589) );
  XNOR2_X2 U667 ( .A(n589), .B(KEYINPUT80), .ZN(n652) );
  INV_X1 U668 ( .A(KEYINPUT2), .ZN(n654) );
  NAND2_X1 U669 ( .A1(KEYINPUT2), .A2(n651), .ZN(n593) );
  XNOR2_X1 U670 ( .A(KEYINPUT77), .B(n593), .ZN(n594) );
  XNOR2_X1 U671 ( .A(n596), .B(KEYINPUT81), .ZN(n598) );
  NOR2_X1 U672 ( .A1(n704), .A2(n599), .ZN(n602) );
  XNOR2_X1 U673 ( .A(n600), .B(KEYINPUT62), .ZN(n601) );
  XNOR2_X1 U674 ( .A(n602), .B(n601), .ZN(n604) );
  INV_X1 U675 ( .A(G952), .ZN(n603) );
  NOR2_X1 U676 ( .A1(n604), .A2(n715), .ZN(n607) );
  XNOR2_X1 U677 ( .A(KEYINPUT107), .B(KEYINPUT63), .ZN(n605) );
  XOR2_X1 U678 ( .A(n605), .B(KEYINPUT83), .Z(n606) );
  XNOR2_X1 U679 ( .A(n607), .B(n606), .ZN(G57) );
  XNOR2_X1 U680 ( .A(n608), .B(G122), .ZN(G24) );
  XNOR2_X1 U681 ( .A(KEYINPUT84), .B(KEYINPUT122), .ZN(n610) );
  XNOR2_X1 U682 ( .A(KEYINPUT59), .B(KEYINPUT66), .ZN(n609) );
  XNOR2_X1 U683 ( .A(n610), .B(n609), .ZN(n611) );
  XNOR2_X1 U684 ( .A(n612), .B(n611), .ZN(n613) );
  XNOR2_X1 U685 ( .A(n614), .B(n613), .ZN(n615) );
  NOR2_X2 U686 ( .A1(n615), .A2(n715), .ZN(n618) );
  XNOR2_X1 U687 ( .A(KEYINPUT123), .B(KEYINPUT60), .ZN(n616) );
  XNOR2_X1 U688 ( .A(n616), .B(KEYINPUT67), .ZN(n617) );
  XNOR2_X1 U689 ( .A(n618), .B(n617), .ZN(G60) );
  XOR2_X1 U690 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n619) );
  XNOR2_X1 U691 ( .A(n620), .B(n619), .ZN(n621) );
  XNOR2_X1 U692 ( .A(n622), .B(n621), .ZN(n623) );
  NOR2_X2 U693 ( .A1(n623), .A2(n715), .ZN(n624) );
  XNOR2_X1 U694 ( .A(n624), .B(KEYINPUT56), .ZN(G51) );
  INV_X1 U695 ( .A(n625), .ZN(n632) );
  NAND2_X1 U696 ( .A1(n632), .A2(n626), .ZN(n627) );
  XNOR2_X1 U697 ( .A(n627), .B(G104), .ZN(G6) );
  XOR2_X1 U698 ( .A(KEYINPUT27), .B(KEYINPUT109), .Z(n629) );
  XNOR2_X1 U699 ( .A(G107), .B(KEYINPUT26), .ZN(n628) );
  XNOR2_X1 U700 ( .A(n629), .B(n628), .ZN(n630) );
  XOR2_X1 U701 ( .A(KEYINPUT108), .B(n630), .Z(n634) );
  NAND2_X1 U702 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U703 ( .A(n634), .B(n633), .ZN(G9) );
  NOR2_X1 U704 ( .A1(n642), .A2(n645), .ZN(n638) );
  XOR2_X1 U705 ( .A(KEYINPUT110), .B(KEYINPUT29), .Z(n636) );
  XNOR2_X1 U706 ( .A(G128), .B(KEYINPUT111), .ZN(n635) );
  XNOR2_X1 U707 ( .A(n636), .B(n635), .ZN(n637) );
  XNOR2_X1 U708 ( .A(n638), .B(n637), .ZN(G30) );
  XNOR2_X1 U709 ( .A(G143), .B(KEYINPUT112), .ZN(n640) );
  XNOR2_X1 U710 ( .A(n640), .B(n639), .ZN(G45) );
  NOR2_X1 U711 ( .A1(n642), .A2(n641), .ZN(n644) );
  XNOR2_X1 U712 ( .A(G146), .B(KEYINPUT113), .ZN(n643) );
  XNOR2_X1 U713 ( .A(n644), .B(n643), .ZN(G48) );
  NOR2_X1 U714 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U715 ( .A(KEYINPUT114), .B(n647), .Z(n648) );
  XNOR2_X1 U716 ( .A(n346), .B(n648), .ZN(G18) );
  XNOR2_X1 U717 ( .A(G125), .B(n649), .ZN(n650) );
  XNOR2_X1 U718 ( .A(n650), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U719 ( .A(G134), .B(n651), .ZN(G36) );
  OR2_X1 U720 ( .A1(n652), .A2(n653), .ZN(n655) );
  NAND2_X1 U721 ( .A1(n655), .A2(n654), .ZN(n657) );
  AND2_X1 U722 ( .A1(n656), .A2(n657), .ZN(n658) );
  XNOR2_X1 U723 ( .A(KEYINPUT79), .B(n658), .ZN(n698) );
  NOR2_X1 U724 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U725 ( .A1(n663), .A2(n662), .ZN(n668) );
  NOR2_X1 U726 ( .A1(n665), .A2(n664), .ZN(n666) );
  XOR2_X1 U727 ( .A(KEYINPUT119), .B(n666), .Z(n667) );
  NOR2_X1 U728 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U729 ( .A(n669), .B(KEYINPUT120), .ZN(n670) );
  NOR2_X1 U730 ( .A1(n693), .A2(n670), .ZN(n689) );
  NAND2_X1 U731 ( .A1(n673), .A2(n672), .ZN(n674) );
  XOR2_X1 U732 ( .A(KEYINPUT50), .B(n674), .Z(n675) );
  NOR2_X1 U733 ( .A1(n492), .A2(n675), .ZN(n681) );
  NOR2_X1 U734 ( .A1(n677), .A2(n676), .ZN(n679) );
  XNOR2_X1 U735 ( .A(KEYINPUT49), .B(KEYINPUT116), .ZN(n678) );
  XNOR2_X1 U736 ( .A(n679), .B(n678), .ZN(n680) );
  NAND2_X1 U737 ( .A1(n681), .A2(n680), .ZN(n683) );
  NAND2_X1 U738 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U739 ( .A(n684), .B(KEYINPUT51), .ZN(n686) );
  XOR2_X1 U740 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n685) );
  XNOR2_X1 U741 ( .A(n686), .B(n685), .ZN(n687) );
  NOR2_X1 U742 ( .A1(n694), .A2(n687), .ZN(n688) );
  NOR2_X1 U743 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U744 ( .A(n690), .B(KEYINPUT52), .ZN(n691) );
  NOR2_X1 U745 ( .A1(n692), .A2(n691), .ZN(n696) );
  NOR2_X1 U746 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U747 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U748 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U749 ( .A1(n699), .A2(G953), .ZN(n700) );
  XNOR2_X1 U750 ( .A(n700), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U751 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n703) );
  XNOR2_X1 U752 ( .A(n701), .B(KEYINPUT121), .ZN(n702) );
  XNOR2_X1 U753 ( .A(n703), .B(n702), .ZN(n706) );
  INV_X1 U754 ( .A(n704), .ZN(n711) );
  NAND2_X1 U755 ( .A1(n711), .A2(G469), .ZN(n705) );
  XOR2_X1 U756 ( .A(n706), .B(n705), .Z(n707) );
  NOR2_X1 U757 ( .A1(n715), .A2(n707), .ZN(G54) );
  NAND2_X1 U758 ( .A1(n711), .A2(G478), .ZN(n709) );
  XNOR2_X1 U759 ( .A(n709), .B(n708), .ZN(n710) );
  NOR2_X1 U760 ( .A1(n715), .A2(n710), .ZN(G63) );
  NAND2_X1 U761 ( .A1(n711), .A2(G217), .ZN(n713) );
  XNOR2_X1 U762 ( .A(n713), .B(n712), .ZN(n714) );
  NOR2_X1 U763 ( .A1(n715), .A2(n714), .ZN(G66) );
  XOR2_X1 U764 ( .A(n716), .B(KEYINPUT125), .Z(n717) );
  XNOR2_X1 U765 ( .A(KEYINPUT124), .B(n717), .ZN(n718) );
  XNOR2_X1 U766 ( .A(n719), .B(n718), .ZN(n722) );
  XNOR2_X1 U767 ( .A(n722), .B(n652), .ZN(n721) );
  NAND2_X1 U768 ( .A1(n721), .A2(n720), .ZN(n727) );
  XNOR2_X1 U769 ( .A(n722), .B(G227), .ZN(n723) );
  XNOR2_X1 U770 ( .A(n723), .B(KEYINPUT126), .ZN(n724) );
  NAND2_X1 U771 ( .A1(n724), .A2(G900), .ZN(n725) );
  NAND2_X1 U772 ( .A1(n725), .A2(G953), .ZN(n726) );
  NAND2_X1 U773 ( .A1(n727), .A2(n726), .ZN(G72) );
  BUF_X1 U774 ( .A(n728), .Z(n729) );
  XOR2_X1 U775 ( .A(G131), .B(n729), .Z(G33) );
  XOR2_X1 U776 ( .A(G137), .B(n730), .Z(G39) );
endmodule

