//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 0 0 1 1 0 1 0 1 1 0 0 0 1 1 1 1 0 1 0 0 0 0 1 1 1 1 0 1 1 0 0 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:10 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370, new_n1371;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT64), .Z(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  AND2_X1   g0015(.A1(KEYINPUT65), .A2(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(KEYINPUT65), .A2(G20), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n203), .A2(G50), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  INV_X1    g0024(.A(G238), .ZN(new_n225));
  INV_X1    g0025(.A(G77), .ZN(new_n226));
  INV_X1    g0026(.A(G244), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n224), .B1(new_n202), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(KEYINPUT66), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n230));
  AOI22_X1  g0030(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n228), .A2(KEYINPUT66), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n212), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  OAI211_X1 g0034(.A(new_n215), .B(new_n223), .C1(new_n234), .C2(KEYINPUT1), .ZN(new_n235));
  AOI21_X1  g0035(.A(new_n235), .B1(KEYINPUT1), .B2(new_n234), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  INV_X1    g0037(.A(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G264), .B(G270), .Z(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G358));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G50), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G68), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n202), .A2(G50), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G58), .B(G77), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n248), .B(new_n254), .ZN(G351));
  OAI21_X1  g0055(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n256));
  INV_X1    g0056(.A(G150), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n210), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT8), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(G58), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n201), .A2(KEYINPUT8), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  OR2_X1    g0063(.A1(KEYINPUT65), .A2(G20), .ZN(new_n264));
  NAND2_X1  g0064(.A1(KEYINPUT65), .A2(G20), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n264), .A2(G33), .A3(new_n265), .ZN(new_n266));
  OAI221_X1 g0066(.A(new_n256), .B1(new_n257), .B2(new_n259), .C1(new_n263), .C2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n268));
  AND2_X1   g0068(.A1(new_n268), .A2(new_n219), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n267), .A2(new_n270), .B1(new_n249), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n269), .A2(new_n271), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT68), .ZN(new_n275));
  AND3_X1   g0075(.A1(new_n271), .A2(new_n219), .A3(new_n268), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT68), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI22_X1  g0078(.A1(new_n275), .A2(new_n278), .B1(new_n209), .B2(G20), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n273), .B1(new_n280), .B2(new_n249), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT3), .B(G33), .ZN(new_n282));
  INV_X1    g0082(.A(G1698), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n282), .A2(G222), .A3(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n282), .A2(G223), .A3(G1698), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n284), .B(new_n285), .C1(new_n226), .C2(new_n282), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G33), .A2(G41), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n287), .A2(G1), .A3(G13), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G179), .ZN(new_n291));
  INV_X1    g0091(.A(G274), .ZN(new_n292));
  AND2_X1   g0092(.A1(G1), .A2(G13), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n292), .B1(new_n293), .B2(new_n287), .ZN(new_n294));
  XNOR2_X1  g0094(.A(KEYINPUT67), .B(G45), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n294), .B(new_n209), .C1(new_n295), .C2(G41), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n288), .A2(G226), .A3(new_n297), .ZN(new_n298));
  AND2_X1   g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n290), .A2(new_n291), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n290), .A2(new_n299), .ZN(new_n301));
  INV_X1    g0101(.A(G169), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AND3_X1   g0103(.A1(new_n281), .A2(new_n300), .A3(new_n303), .ZN(new_n304));
  XNOR2_X1  g0104(.A(new_n281), .B(KEYINPUT9), .ZN(new_n305));
  INV_X1    g0105(.A(G190), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n307), .B1(G200), .B2(new_n301), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(KEYINPUT10), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT10), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n305), .A2(new_n311), .A3(new_n308), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n304), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  NOR2_X1   g0113(.A1(G20), .A2(G33), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n314), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n315), .B1(new_n266), .B2(new_n226), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n270), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT11), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n316), .A2(KEYINPUT11), .A3(new_n270), .ZN(new_n320));
  OR3_X1    g0120(.A1(new_n271), .A2(KEYINPUT12), .A3(G68), .ZN(new_n321));
  OAI21_X1  g0121(.A(KEYINPUT12), .B1(new_n271), .B2(G68), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n202), .B1(new_n209), .B2(G20), .ZN(new_n323));
  AOI22_X1  g0123(.A1(new_n321), .A2(new_n322), .B1(new_n276), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n319), .A2(new_n320), .A3(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n288), .A2(G238), .A3(new_n297), .ZN(new_n327));
  NAND2_X1  g0127(.A1(G33), .A2(G97), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  NOR2_X1   g0129(.A1(G226), .A2(G1698), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n330), .B1(new_n238), .B2(G1698), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n329), .B1(new_n331), .B2(new_n282), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n296), .B(new_n327), .C1(new_n332), .C2(new_n288), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(KEYINPUT13), .ZN(new_n334));
  AND3_X1   g0134(.A1(new_n288), .A2(G238), .A3(new_n297), .ZN(new_n335));
  INV_X1    g0135(.A(G226), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n283), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n238), .A2(G1698), .ZN(new_n338));
  AND2_X1   g0138(.A1(KEYINPUT3), .A2(G33), .ZN(new_n339));
  NOR2_X1   g0139(.A1(KEYINPUT3), .A2(G33), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n337), .B(new_n338), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n328), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n335), .B1(new_n342), .B2(new_n289), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT13), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n343), .A2(new_n344), .A3(new_n296), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n334), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n326), .B1(new_n346), .B2(new_n306), .ZN(new_n347));
  INV_X1    g0147(.A(G200), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n348), .B1(new_n334), .B2(new_n345), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n333), .A2(KEYINPUT13), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n344), .B1(new_n343), .B2(new_n296), .ZN(new_n352));
  OAI21_X1  g0152(.A(G169), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(KEYINPUT14), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n334), .A2(new_n345), .A3(G179), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT14), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n356), .B(G169), .C1(new_n351), .C2(new_n352), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n354), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n350), .B1(new_n358), .B2(new_n325), .ZN(new_n359));
  OAI211_X1 g0159(.A(G232), .B(new_n283), .C1(new_n339), .C2(new_n340), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(KEYINPUT69), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT69), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n282), .A2(new_n362), .A3(G232), .A4(new_n283), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n282), .A2(G238), .A3(G1698), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n339), .A2(new_n340), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(G107), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n361), .A2(new_n363), .A3(new_n364), .A4(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n289), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n288), .A2(G244), .A3(new_n297), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n296), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n368), .A2(new_n291), .A3(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(KEYINPUT70), .B1(new_n261), .B2(new_n262), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n201), .A2(KEYINPUT8), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n260), .A2(G58), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT70), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n259), .B1(new_n373), .B2(new_n377), .ZN(new_n378));
  XNOR2_X1  g0178(.A(KEYINPUT15), .B(G87), .ZN(new_n379));
  OAI22_X1  g0179(.A1(new_n266), .A2(new_n379), .B1(new_n218), .B2(new_n226), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n270), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n226), .B1(new_n209), .B2(G20), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n276), .A2(new_n382), .B1(new_n226), .B2(new_n272), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n370), .B1(new_n367), .B2(new_n289), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n372), .B(new_n384), .C1(G169), .C2(new_n385), .ZN(new_n386));
  AND2_X1   g0186(.A1(new_n381), .A2(new_n383), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n368), .A2(G190), .A3(new_n371), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n387), .B(new_n388), .C1(new_n348), .C2(new_n385), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n313), .A2(new_n359), .A3(new_n386), .A4(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT18), .ZN(new_n391));
  OR2_X1    g0191(.A1(new_n391), .A2(KEYINPUT72), .ZN(new_n392));
  INV_X1    g0192(.A(new_n263), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n393), .A2(new_n272), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(new_n279), .B2(new_n263), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT7), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n218), .A2(new_n365), .A3(new_n397), .ZN(new_n398));
  OR2_X1    g0198(.A1(KEYINPUT3), .A2(G33), .ZN(new_n399));
  NAND2_X1  g0199(.A1(KEYINPUT3), .A2(G33), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n399), .A2(new_n210), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(KEYINPUT7), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n398), .A2(new_n402), .A3(G68), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT71), .ZN(new_n404));
  NAND2_X1  g0204(.A1(G58), .A2(G68), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n210), .B1(new_n203), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n314), .A2(G159), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n404), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  AND2_X1   g0209(.A1(G58), .A2(G68), .ZN(new_n410));
  NOR2_X1   g0210(.A1(G58), .A2(G68), .ZN(new_n411));
  OAI21_X1  g0211(.A(G20), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n412), .A2(KEYINPUT71), .A3(new_n407), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n403), .A2(KEYINPUT16), .A3(new_n409), .A4(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n270), .ZN(new_n415));
  AND3_X1   g0215(.A1(new_n412), .A2(KEYINPUT71), .A3(new_n407), .ZN(new_n416));
  AOI21_X1  g0216(.A(KEYINPUT71), .B1(new_n412), .B2(new_n407), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n264), .A2(new_n265), .ZN(new_n419));
  OAI21_X1  g0219(.A(KEYINPUT7), .B1(new_n419), .B2(new_n282), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n365), .A2(new_n397), .A3(new_n210), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n420), .A2(G68), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT16), .B1(new_n418), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n396), .B1(new_n415), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n288), .A2(G232), .A3(new_n297), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n296), .A2(new_n425), .ZN(new_n426));
  OR2_X1    g0226(.A1(G223), .A2(G1698), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n336), .A2(G1698), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n282), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(G33), .A2(G87), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n288), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(G169), .B1(new_n426), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n427), .A2(new_n428), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n430), .B1(new_n433), .B2(new_n365), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n289), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n435), .A2(G179), .A3(new_n296), .A4(new_n425), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n392), .B1(new_n424), .B2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n437), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT16), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n420), .A2(G68), .A3(new_n421), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n409), .A2(new_n413), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n440), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n443), .A2(new_n270), .A3(new_n414), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n439), .B1(new_n444), .B2(new_n396), .ZN(new_n445));
  XNOR2_X1  g0245(.A(KEYINPUT72), .B(KEYINPUT18), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n438), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n348), .B1(new_n426), .B2(new_n431), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n435), .A2(new_n306), .A3(new_n296), .A4(new_n425), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n450), .B(new_n396), .C1(new_n415), .C2(new_n423), .ZN(new_n451));
  XNOR2_X1  g0251(.A(new_n451), .B(KEYINPUT17), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n447), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g0253(.A(new_n453), .B(KEYINPUT73), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n390), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n258), .A2(G97), .ZN(new_n456));
  NAND2_X1  g0256(.A1(G33), .A2(G283), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n264), .A2(new_n456), .A3(new_n265), .A4(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(G116), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n268), .A2(new_n219), .B1(G20), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT20), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n458), .A2(KEYINPUT20), .A3(new_n460), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n209), .A2(G33), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n276), .A2(KEYINPUT78), .A3(G116), .A4(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT78), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n271), .A2(new_n466), .A3(new_n219), .A4(new_n268), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n468), .B1(new_n469), .B2(new_n459), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n272), .A2(new_n459), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n465), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  OAI211_X1 g0273(.A(G264), .B(G1698), .C1(new_n339), .C2(new_n340), .ZN(new_n474));
  OAI211_X1 g0274(.A(G257), .B(new_n283), .C1(new_n339), .C2(new_n340), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n399), .A2(G303), .A3(new_n400), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n289), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n209), .A2(G45), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT5), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n479), .B1(new_n480), .B2(G41), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT75), .ZN(new_n482));
  INV_X1    g0282(.A(G41), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n482), .A2(new_n483), .A3(KEYINPUT5), .ZN(new_n484));
  OAI21_X1  g0284(.A(KEYINPUT75), .B1(new_n480), .B2(G41), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n481), .A2(new_n294), .A3(new_n484), .A4(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n480), .A2(G41), .ZN(new_n487));
  INV_X1    g0287(.A(G45), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n488), .A2(G1), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n485), .A2(new_n484), .A3(new_n487), .A4(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n490), .A2(G270), .A3(new_n288), .ZN(new_n491));
  AND3_X1   g0291(.A1(new_n478), .A2(new_n486), .A3(new_n491), .ZN(new_n492));
  AND3_X1   g0292(.A1(new_n473), .A2(new_n492), .A3(G179), .ZN(new_n493));
  INV_X1    g0293(.A(new_n471), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n458), .A2(KEYINPUT20), .A3(new_n460), .ZN(new_n495));
  AOI21_X1  g0295(.A(KEYINPUT20), .B1(new_n458), .B2(new_n460), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n472), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n478), .A2(new_n486), .A3(new_n491), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT21), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n500), .A2(new_n302), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(KEYINPUT79), .B1(new_n498), .B2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n501), .ZN(new_n504));
  AND2_X1   g0304(.A1(new_n491), .A2(new_n486), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n504), .B1(new_n505), .B2(new_n478), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT79), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n506), .A2(new_n507), .A3(new_n473), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n493), .B1(new_n503), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n492), .A2(G190), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n499), .A2(G200), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n510), .A2(new_n498), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n302), .B1(new_n505), .B2(new_n478), .ZN(new_n513));
  AOI211_X1 g0313(.A(KEYINPUT80), .B(KEYINPUT21), .C1(new_n513), .C2(new_n473), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT80), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n499), .B(G169), .C1(new_n494), .C2(new_n497), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n515), .B1(new_n516), .B2(new_n500), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n509), .B(new_n512), .C1(new_n514), .C2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(G250), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n283), .ZN(new_n520));
  INV_X1    g0320(.A(G257), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(G1698), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n520), .B(new_n522), .C1(new_n339), .C2(new_n340), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G33), .A2(G294), .ZN(new_n524));
  AND3_X1   g0324(.A1(new_n523), .A2(KEYINPUT83), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(KEYINPUT83), .B1(new_n523), .B2(new_n524), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n289), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n490), .A2(G264), .A3(new_n288), .ZN(new_n528));
  AND2_X1   g0328(.A1(new_n528), .A2(new_n486), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n527), .A2(new_n529), .A3(KEYINPUT84), .A4(new_n306), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT84), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n527), .A2(new_n529), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n531), .B1(new_n532), .B2(new_n348), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n532), .A2(G190), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n530), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  OR2_X1    g0335(.A1(new_n469), .A2(KEYINPUT74), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n469), .A2(KEYINPUT74), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n536), .A2(G107), .A3(new_n537), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n271), .A2(G107), .ZN(new_n539));
  XNOR2_X1  g0339(.A(KEYINPUT82), .B(KEYINPUT25), .ZN(new_n540));
  XNOR2_X1  g0340(.A(new_n539), .B(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n218), .A2(new_n282), .A3(G87), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT22), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n544), .A2(KEYINPUT81), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(new_n545), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n218), .A2(new_n282), .A3(new_n547), .A4(G87), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT23), .ZN(new_n550));
  INV_X1    g0350(.A(G107), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(G33), .A2(G116), .ZN(new_n553));
  AOI21_X1  g0353(.A(G20), .B1(new_n553), .B2(new_n550), .ZN(new_n554));
  NOR2_X1   g0354(.A1(KEYINPUT23), .A2(G107), .ZN(new_n555));
  AOI211_X1 g0355(.A(new_n552), .B(new_n554), .C1(new_n419), .C2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n549), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(KEYINPUT24), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT24), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n549), .A2(new_n559), .A3(new_n556), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n542), .B1(new_n561), .B2(new_n270), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n535), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n527), .A2(new_n529), .A3(new_n291), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n523), .A2(new_n524), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT83), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n523), .A2(KEYINPUT83), .A3(new_n524), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n288), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n528), .A2(new_n486), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n302), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n269), .B1(new_n558), .B2(new_n560), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n564), .B(new_n571), .C1(new_n572), .C2(new_n542), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n563), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n518), .A2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT77), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n271), .A2(G97), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT6), .ZN(new_n578));
  AND2_X1   g0378(.A1(G97), .A2(G107), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n578), .B1(new_n579), .B2(new_n205), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n551), .A2(KEYINPUT6), .A3(G97), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n582), .A2(new_n419), .B1(G77), .B2(new_n314), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n420), .A2(G107), .A3(new_n421), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n577), .B1(new_n585), .B2(new_n270), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n536), .A2(G97), .A3(new_n537), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n490), .A2(G257), .A3(new_n288), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n486), .ZN(new_n589));
  OAI211_X1 g0389(.A(G244), .B(new_n283), .C1(new_n339), .C2(new_n340), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT4), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n282), .A2(KEYINPUT4), .A3(G244), .A4(new_n283), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n282), .A2(G250), .A3(G1698), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n592), .A2(new_n593), .A3(new_n457), .A4(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n589), .B1(new_n289), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n586), .A2(new_n587), .B1(new_n596), .B2(new_n291), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n595), .A2(new_n289), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n588), .A2(new_n486), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n302), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n598), .A2(new_n306), .A3(new_n599), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(new_n596), .B2(G200), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n269), .B1(new_n583), .B2(new_n584), .ZN(new_n604));
  INV_X1    g0404(.A(new_n587), .ZN(new_n605));
  NOR3_X1   g0405(.A1(new_n604), .A2(new_n605), .A3(new_n577), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n597), .A2(new_n601), .B1(new_n603), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n264), .A2(G33), .A3(G97), .A4(new_n265), .ZN(new_n609));
  XOR2_X1   g0409(.A(KEYINPUT76), .B(KEYINPUT19), .Z(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n218), .A2(new_n282), .A3(G68), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n206), .A2(G87), .ZN(new_n614));
  XNOR2_X1  g0414(.A(KEYINPUT76), .B(KEYINPUT19), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n329), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n614), .B1(new_n616), .B2(new_n218), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n270), .B1(new_n613), .B2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n379), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n619), .A2(new_n271), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n536), .A2(new_n619), .A3(new_n537), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n618), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n479), .A2(new_n519), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n209), .A2(new_n292), .A3(G45), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n624), .A2(new_n288), .A3(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(G238), .A2(G1698), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n627), .B1(new_n227), .B2(G1698), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n628), .A2(new_n282), .B1(G33), .B2(G116), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n291), .B(new_n626), .C1(new_n629), .C2(new_n288), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n225), .A2(new_n283), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n227), .A2(G1698), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n631), .B(new_n632), .C1(new_n339), .C2(new_n340), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n288), .B1(new_n633), .B2(new_n553), .ZN(new_n634));
  INV_X1    g0434(.A(new_n626), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n302), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n630), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n623), .A2(new_n637), .ZN(new_n638));
  OR2_X1    g0438(.A1(KEYINPUT76), .A2(KEYINPUT19), .ZN(new_n639));
  NAND2_X1  g0439(.A1(KEYINPUT76), .A2(KEYINPUT19), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n328), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI22_X1  g0441(.A1(new_n641), .A2(new_n419), .B1(G87), .B2(new_n206), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n642), .A2(new_n612), .A3(new_n611), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n620), .B1(new_n643), .B2(new_n270), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n626), .B1(new_n629), .B2(new_n288), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(G200), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n536), .A2(G87), .A3(new_n537), .ZN(new_n647));
  OAI211_X1 g0447(.A(G190), .B(new_n626), .C1(new_n629), .C2(new_n288), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n644), .A2(new_n646), .A3(new_n647), .A4(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n638), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n576), .B1(new_n608), .B2(new_n650), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n607), .A2(KEYINPUT77), .A3(new_n638), .A4(new_n649), .ZN(new_n652));
  AND4_X1   g0452(.A1(new_n455), .A2(new_n575), .A3(new_n651), .A4(new_n652), .ZN(G372));
  AND3_X1   g0453(.A1(new_n424), .A2(new_n437), .A3(KEYINPUT86), .ZN(new_n654));
  AOI21_X1  g0454(.A(KEYINPUT86), .B1(new_n424), .B2(new_n437), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n391), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n424), .A2(new_n437), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT86), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n424), .A2(new_n437), .A3(KEYINPUT86), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(KEYINPUT18), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n656), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT17), .ZN(new_n664));
  XNOR2_X1  g0464(.A(new_n451), .B(new_n664), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n347), .A2(new_n349), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT87), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n384), .B1(new_n385), .B2(G169), .ZN(new_n668));
  AOI211_X1 g0468(.A(G179), .B(new_n370), .C1(new_n289), .C2(new_n367), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n368), .A2(new_n371), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(new_n302), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n672), .A2(KEYINPUT87), .A3(new_n372), .A4(new_n384), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n666), .A2(new_n670), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n357), .A2(new_n355), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n356), .B1(new_n346), .B2(G169), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n325), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n665), .B1(new_n674), .B2(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n663), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n679), .B1(new_n310), .B2(new_n312), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(new_n304), .ZN(new_n681));
  AND4_X1   g0481(.A1(new_n618), .A2(new_n621), .A3(new_n647), .A4(new_n648), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n634), .A2(new_n635), .ZN(new_n683));
  OAI21_X1  g0483(.A(KEYINPUT85), .B1(new_n683), .B2(new_n348), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT85), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n645), .A2(new_n685), .A3(G200), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  AOI22_X1  g0487(.A1(new_n682), .A2(new_n687), .B1(new_n623), .B2(new_n637), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT26), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n688), .A2(new_n689), .A3(new_n601), .A4(new_n597), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n585), .A2(new_n270), .ZN(new_n691));
  INV_X1    g0491(.A(new_n577), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(new_n587), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n596), .A2(new_n291), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n693), .A2(new_n694), .A3(new_n601), .ZN(new_n695));
  OAI21_X1  g0495(.A(KEYINPUT26), .B1(new_n695), .B2(new_n650), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n690), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n514), .A2(new_n517), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n499), .A2(new_n291), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(new_n473), .ZN(new_n700));
  AND4_X1   g0500(.A1(new_n507), .A2(new_n473), .A3(new_n499), .A4(new_n501), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n507), .B1(new_n506), .B2(new_n473), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n700), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n571), .A2(new_n564), .ZN(new_n704));
  INV_X1    g0504(.A(new_n560), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n559), .B1(new_n549), .B2(new_n556), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n270), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n542), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n704), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NOR3_X1   g0509(.A1(new_n698), .A2(new_n703), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n682), .A2(new_n687), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n563), .A2(new_n607), .A3(new_n711), .ZN(new_n712));
  OAI211_X1 g0512(.A(new_n697), .B(new_n638), .C1(new_n710), .C2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n455), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n681), .A2(new_n714), .ZN(G369));
  INV_X1    g0515(.A(G330), .ZN(new_n716));
  OR2_X1    g0516(.A1(new_n514), .A2(new_n517), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n218), .A2(new_n209), .A3(G13), .ZN(new_n718));
  OR2_X1    g0518(.A1(new_n718), .A2(KEYINPUT27), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(KEYINPUT27), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n719), .A2(G213), .A3(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(G343), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(new_n473), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n717), .A2(new_n509), .A3(new_n512), .A4(new_n724), .ZN(new_n725));
  OAI211_X1 g0525(.A(new_n473), .B(new_n723), .C1(new_n698), .C2(new_n703), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n716), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n723), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n562), .A2(new_n728), .ZN(new_n729));
  OAI22_X1  g0529(.A1(new_n574), .A2(new_n729), .B1(new_n573), .B2(new_n728), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n727), .A2(KEYINPUT88), .A3(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(KEYINPUT88), .B1(new_n727), .B2(new_n730), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n723), .B1(new_n717), .B2(new_n509), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n709), .B1(new_n562), .B2(new_n535), .ZN(new_n736));
  AOI22_X1  g0536(.A1(new_n735), .A2(new_n736), .B1(new_n709), .B2(new_n728), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n734), .A2(new_n737), .ZN(G399));
  INV_X1    g0538(.A(new_n213), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(G41), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(new_n209), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n614), .A2(new_n459), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI22_X1  g0543(.A1(new_n741), .A2(new_n743), .B1(new_n222), .B2(new_n740), .ZN(new_n744));
  XOR2_X1   g0544(.A(new_n744), .B(KEYINPUT28), .Z(new_n745));
  NAND4_X1  g0545(.A1(new_n575), .A2(new_n651), .A3(new_n652), .A4(new_n728), .ZN(new_n746));
  AND3_X1   g0546(.A1(new_n527), .A2(new_n528), .A3(new_n683), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n747), .A2(new_n699), .A3(new_n596), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT30), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(KEYINPUT89), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n683), .A2(G179), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n600), .A2(new_n532), .A3(new_n499), .A4(new_n753), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n747), .A2(new_n699), .A3(new_n596), .A4(new_n750), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n752), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n756), .A2(KEYINPUT31), .A3(new_n723), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(KEYINPUT31), .B1(new_n756), .B2(new_n723), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n716), .B1(new_n746), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n689), .B1(new_n695), .B2(new_n650), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n688), .A2(new_n601), .A3(new_n597), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n762), .B1(new_n763), .B2(new_n689), .ZN(new_n764));
  OAI211_X1 g0564(.A(new_n638), .B(new_n764), .C1(new_n710), .C2(new_n712), .ZN(new_n765));
  AND3_X1   g0565(.A1(new_n765), .A2(KEYINPUT90), .A3(new_n728), .ZN(new_n766));
  AOI21_X1  g0566(.A(KEYINPUT90), .B1(new_n765), .B2(new_n728), .ZN(new_n767));
  OAI21_X1  g0567(.A(KEYINPUT29), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n713), .A2(new_n728), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT29), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n761), .B1(new_n768), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n745), .B1(new_n772), .B2(G1), .ZN(G364));
  INV_X1    g0573(.A(G13), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n419), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G45), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n741), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n727), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n725), .A2(new_n716), .A3(new_n726), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n778), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n774), .A2(new_n258), .A3(KEYINPUT91), .ZN(new_n782));
  INV_X1    g0582(.A(KEYINPUT91), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n783), .B1(G13), .B2(G33), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(G20), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n219), .B1(G20), .B2(new_n302), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n739), .A2(new_n282), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n791), .B1(new_n221), .B2(new_n295), .C1(new_n254), .C2(new_n488), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n739), .A2(new_n365), .ZN(new_n793));
  AOI22_X1  g0593(.A1(G355), .A2(new_n793), .B1(new_n459), .B2(new_n739), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n790), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n218), .A2(new_n291), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G200), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G190), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT92), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(G326), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n306), .A2(G200), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n218), .B1(new_n291), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(G179), .A2(G200), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n419), .A2(new_n306), .A3(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n805), .A2(G294), .B1(new_n808), .B2(G329), .ZN(new_n809));
  NOR2_X1   g0609(.A1(G190), .A2(G200), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n796), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n796), .A2(new_n803), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n812), .A2(G311), .B1(new_n814), .B2(G322), .ZN(new_n815));
  INV_X1    g0615(.A(G303), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n348), .A2(G179), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n817), .A2(G20), .A3(G190), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n419), .A2(new_n306), .A3(new_n817), .ZN(new_n819));
  INV_X1    g0619(.A(G283), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n365), .B1(new_n816), .B2(new_n818), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n798), .A2(new_n306), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  XNOR2_X1  g0623(.A(KEYINPUT33), .B(G317), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n821), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n802), .A2(new_n809), .A3(new_n815), .A4(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT32), .ZN(new_n827));
  INV_X1    g0627(.A(G159), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n807), .A2(new_n828), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n822), .A2(new_n202), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(new_n827), .B2(new_n829), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n805), .A2(G97), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n812), .A2(G77), .B1(new_n814), .B2(G58), .ZN(new_n833));
  INV_X1    g0633(.A(G87), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n282), .B1(new_n834), .B2(new_n818), .C1(new_n819), .C2(new_n551), .ZN(new_n835));
  INV_X1    g0635(.A(new_n799), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n835), .B1(new_n836), .B2(G50), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n831), .A2(new_n832), .A3(new_n833), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n826), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n795), .B1(new_n839), .B2(new_n788), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n787), .B(KEYINPUT93), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n725), .A2(new_n726), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n777), .B1(new_n840), .B2(new_n843), .ZN(new_n844));
  OR2_X1    g0644(.A1(new_n781), .A2(new_n844), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n845), .A2(KEYINPUT94), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n845), .A2(KEYINPUT94), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n846), .A2(new_n847), .ZN(G396));
  NAND2_X1  g0648(.A1(new_n723), .A2(new_n384), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  AND4_X1   g0650(.A1(KEYINPUT95), .A2(new_n670), .A3(new_n673), .A4(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n670), .A2(new_n673), .A3(new_n850), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n389), .A2(new_n386), .A3(new_n849), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT95), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n851), .B1(new_n852), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n769), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n713), .A2(new_n728), .A3(new_n856), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n761), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(new_n741), .B2(new_n776), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n858), .A2(new_n761), .A3(new_n859), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n788), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n786), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n818), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n282), .B1(new_n866), .B2(G107), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n832), .B(new_n867), .C1(new_n799), .C2(new_n816), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n819), .A2(new_n834), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n869), .B1(new_n812), .B2(G116), .ZN(new_n870));
  INV_X1    g0670(.A(G294), .ZN(new_n871));
  INV_X1    g0671(.A(G311), .ZN(new_n872));
  OAI221_X1 g0672(.A(new_n870), .B1(new_n871), .B2(new_n813), .C1(new_n872), .C2(new_n807), .ZN(new_n873));
  AOI211_X1 g0673(.A(new_n868), .B(new_n873), .C1(G283), .C2(new_n823), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n812), .A2(G159), .B1(new_n814), .B2(G143), .ZN(new_n875));
  INV_X1    g0675(.A(G137), .ZN(new_n876));
  OAI221_X1 g0676(.A(new_n875), .B1(new_n822), .B2(new_n257), .C1(new_n876), .C2(new_n799), .ZN(new_n877));
  XNOR2_X1  g0677(.A(new_n877), .B(KEYINPUT34), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n282), .B1(new_n818), .B2(new_n249), .ZN(new_n879));
  INV_X1    g0679(.A(G132), .ZN(new_n880));
  OAI22_X1  g0680(.A1(new_n202), .A2(new_n819), .B1(new_n807), .B2(new_n880), .ZN(new_n881));
  AOI211_X1 g0681(.A(new_n879), .B(new_n881), .C1(G58), .C2(new_n805), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n874), .B1(new_n878), .B2(new_n882), .ZN(new_n883));
  OAI221_X1 g0683(.A(new_n778), .B1(G77), .B2(new_n865), .C1(new_n883), .C2(new_n864), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(new_n785), .B2(new_n857), .ZN(new_n885));
  XOR2_X1   g0685(.A(new_n885), .B(KEYINPUT96), .Z(new_n886));
  NOR2_X1   g0686(.A1(new_n863), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(G384));
  NOR2_X1   g0688(.A1(new_n775), .A2(new_n209), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT38), .ZN(new_n890));
  INV_X1    g0690(.A(new_n721), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n424), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT37), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n657), .A2(new_n892), .A3(new_n893), .A4(new_n451), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT98), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT37), .B1(new_n424), .B2(new_n437), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n897), .A2(KEYINPUT98), .A3(new_n451), .A4(new_n892), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n403), .A2(new_n409), .A3(new_n413), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT16), .B1(new_n899), .B2(KEYINPUT97), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT97), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n418), .A2(new_n901), .A3(new_n403), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n415), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n396), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n437), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n891), .B1(new_n903), .B2(new_n904), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n905), .A2(new_n906), .A3(new_n451), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n896), .A2(new_n898), .B1(new_n907), .B2(KEYINPUT37), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n906), .B1(new_n447), .B2(new_n452), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n890), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n899), .A2(KEYINPUT97), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n911), .A2(new_n440), .A3(new_n902), .ZN(new_n912));
  INV_X1    g0712(.A(new_n415), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n904), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n451), .B1(new_n914), .B2(new_n721), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n914), .A2(new_n439), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT37), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n451), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n721), .B1(new_n444), .B2(new_n396), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT98), .B1(new_n920), .B2(new_n897), .ZN(new_n921));
  INV_X1    g0721(.A(new_n898), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n917), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n906), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n453), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n923), .A2(KEYINPUT38), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n910), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n723), .A2(new_n325), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n677), .A2(new_n666), .A3(new_n928), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n325), .B(new_n723), .C1(new_n358), .C2(new_n350), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n856), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(new_n746), .B2(new_n760), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n927), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT40), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(KEYINPUT99), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT99), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n934), .A2(new_n938), .A3(new_n935), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  AOI211_X1 g0740(.A(new_n935), .B(new_n932), .C1(new_n746), .C2(new_n760), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n892), .B1(new_n662), .B2(new_n452), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n451), .B(new_n892), .C1(new_n654), .C2(new_n655), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n896), .A2(new_n898), .B1(new_n943), .B2(KEYINPUT37), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n890), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n926), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n941), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n940), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n746), .A2(new_n760), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n455), .A2(new_n949), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n948), .A2(new_n950), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n951), .A2(G330), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(KEYINPUT39), .B1(new_n945), .B2(new_n926), .ZN(new_n954));
  AND3_X1   g0754(.A1(new_n910), .A2(new_n926), .A3(KEYINPUT39), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n358), .A2(new_n325), .A3(new_n728), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n931), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n386), .A2(new_n723), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n960), .B1(new_n859), .B2(new_n962), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n963), .A2(new_n927), .B1(new_n663), .B2(new_n721), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n959), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n768), .A2(new_n455), .A3(new_n771), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n681), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n965), .B(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n889), .B1(new_n953), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n968), .B2(new_n953), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n582), .A2(KEYINPUT35), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n582), .A2(KEYINPUT35), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n971), .A2(G116), .A3(new_n220), .A4(new_n972), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT36), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n405), .A2(G77), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n250), .B1(new_n221), .B2(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n976), .A2(G1), .A3(new_n774), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n970), .A2(new_n974), .A3(new_n977), .ZN(G367));
  OAI21_X1  g0778(.A(new_n607), .B1(new_n606), .B2(new_n728), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n597), .A2(new_n601), .A3(new_n723), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n981), .A2(new_n736), .A3(new_n735), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n982), .A2(KEYINPUT42), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n695), .B1(new_n979), .B2(new_n573), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n982), .A2(KEYINPUT42), .B1(new_n728), .B2(new_n984), .ZN(new_n985));
  AND2_X1   g0785(.A1(new_n644), .A2(new_n647), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n688), .B1(new_n986), .B2(new_n728), .ZN(new_n987));
  OR3_X1    g0787(.A1(new_n986), .A2(new_n638), .A3(new_n728), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n983), .A2(new_n985), .B1(KEYINPUT43), .B2(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n989), .A2(KEYINPUT43), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n990), .B(new_n991), .Z(new_n992));
  INV_X1    g0792(.A(new_n981), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n734), .A2(new_n993), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n992), .B(new_n994), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n740), .B(KEYINPUT41), .Z(new_n996));
  NAND2_X1  g0796(.A1(new_n735), .A2(new_n736), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n730), .B2(new_n735), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT102), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT103), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n997), .B(KEYINPUT102), .C1(new_n730), .C2(new_n735), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n1000), .A2(new_n1001), .A3(new_n779), .A4(new_n1002), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n998), .A2(new_n779), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n727), .B1(new_n998), .B2(new_n999), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1001), .B1(new_n1006), .B2(new_n1002), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT45), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n709), .A2(new_n728), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n997), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1009), .B1(new_n1011), .B2(new_n993), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n737), .A2(KEYINPUT45), .A3(new_n981), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1011), .A2(KEYINPUT44), .A3(new_n993), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT44), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n737), .B2(new_n981), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1014), .A2(new_n1018), .A3(KEYINPUT100), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n734), .B1(new_n1019), .B2(KEYINPUT101), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n1013), .A2(new_n1012), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1021));
  OAI21_X1  g0821(.A(KEYINPUT101), .B1(new_n732), .B2(new_n733), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1021), .B1(new_n1022), .B2(KEYINPUT100), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n772), .B(new_n1008), .C1(new_n1020), .C2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n996), .B1(new_n1024), .B2(new_n772), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n776), .A2(G1), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n995), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n791), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1028), .A2(new_n244), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n789), .B1(new_n213), .B2(new_n379), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n282), .B1(new_n813), .B2(new_n257), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n805), .A2(G68), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1032), .B1(new_n226), .B2(new_n819), .C1(new_n811), .C2(new_n249), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n1031), .B(new_n1033), .C1(G159), .C2(new_n823), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n801), .A2(G143), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n807), .A2(new_n876), .B1(new_n201), .B2(new_n818), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT105), .Z(new_n1037));
  NAND3_X1  g0837(.A1(new_n1034), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT106), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n800), .A2(new_n872), .B1(new_n816), .B2(new_n813), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n1040), .A2(KEYINPUT104), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1040), .A2(KEYINPUT104), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n819), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n805), .A2(G107), .B1(new_n1043), .B2(G97), .ZN(new_n1044));
  INV_X1    g0844(.A(G317), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1044), .B1(new_n820), .B2(new_n811), .C1(new_n1045), .C2(new_n807), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n866), .A2(G116), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT46), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n282), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1049), .B1(new_n1048), .B2(new_n1047), .C1(new_n822), .C2(new_n871), .ZN(new_n1050));
  NOR4_X1   g0850(.A1(new_n1041), .A2(new_n1042), .A3(new_n1046), .A4(new_n1050), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n1039), .A2(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT47), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n778), .B1(new_n1029), .B2(new_n1030), .C1(new_n1053), .C2(new_n864), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT107), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1056), .B(new_n1057), .C1(new_n841), .C2(new_n989), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1027), .A2(new_n1058), .ZN(G387));
  INV_X1    g0859(.A(new_n772), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n1007), .B2(new_n1005), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1008), .A2(new_n772), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1061), .A2(new_n740), .A3(new_n1062), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n730), .A2(new_n841), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n793), .A2(new_n742), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(G107), .B2(new_n213), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1028), .B1(new_n241), .B2(new_n295), .ZN(new_n1067));
  AOI21_X1  g0867(.A(G50), .B1(new_n373), .B2(new_n377), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1071));
  AOI21_X1  g0871(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1070), .A2(new_n743), .A3(new_n1071), .A4(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1066), .B1(new_n1067), .B2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n778), .B1(new_n1074), .B2(new_n790), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n804), .A2(new_n379), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n811), .A2(new_n202), .B1(new_n257), .B2(new_n807), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n1076), .B(new_n1077), .C1(G50), .C2(new_n814), .ZN(new_n1078));
  INV_X1    g0878(.A(G97), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n282), .B1(new_n226), .B2(new_n818), .C1(new_n819), .C2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n823), .B2(new_n393), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1078), .B(new_n1081), .C1(new_n828), .C2(new_n799), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n282), .B1(new_n808), .B2(G326), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n804), .A2(new_n820), .B1(new_n871), .B2(new_n818), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n812), .A2(G303), .B1(new_n814), .B2(G317), .ZN(new_n1085));
  INV_X1    g0885(.A(G322), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n1085), .B1(new_n872), .B2(new_n822), .C1(new_n800), .C2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT48), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1084), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n1088), .B2(new_n1087), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT49), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n1083), .B1(new_n459), .B2(new_n819), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1082), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1075), .B1(new_n1094), .B2(new_n788), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n1008), .A2(new_n1026), .B1(new_n1064), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1063), .A2(new_n1096), .ZN(G393));
  NAND2_X1  g0897(.A1(new_n1021), .A2(new_n734), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT109), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  OR2_X1    g0900(.A1(new_n1021), .A2(new_n734), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1021), .A2(new_n734), .A3(KEYINPUT109), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1100), .A2(new_n1101), .A3(new_n1026), .A4(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n789), .B1(new_n1079), .B2(new_n213), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1028), .A2(new_n248), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n778), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n799), .A2(new_n1045), .B1(new_n872), .B2(new_n813), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT52), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n812), .A2(G294), .B1(new_n805), .B2(G116), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1108), .B(new_n1109), .C1(new_n816), .C2(new_n822), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n282), .B1(new_n866), .B2(G283), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n1111), .B1(new_n551), .B2(new_n819), .C1(new_n1086), .C2(new_n807), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT110), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n799), .A2(new_n257), .B1(new_n828), .B2(new_n813), .ZN(new_n1114));
  XOR2_X1   g0914(.A(new_n1114), .B(KEYINPUT51), .Z(new_n1115));
  NAND2_X1  g0915(.A1(new_n823), .A2(G50), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n365), .B(new_n869), .C1(G68), .C2(new_n866), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n808), .A2(G143), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n804), .A2(new_n226), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n373), .A2(new_n377), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1119), .B1(new_n1120), .B2(new_n812), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1116), .A2(new_n1117), .A3(new_n1118), .A4(new_n1121), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n1110), .A2(new_n1113), .B1(new_n1115), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1106), .B1(new_n1123), .B2(new_n788), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n787), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1124), .B1(new_n1125), .B2(new_n981), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1103), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n740), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n1019), .A2(KEYINPUT101), .ZN(new_n1129));
  AND2_X1   g0929(.A1(new_n1022), .A2(KEYINPUT100), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n1129), .A2(new_n734), .B1(new_n1130), .B2(new_n1021), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1062), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1128), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n1062), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1127), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(G390));
  NAND2_X1  g0937(.A1(new_n859), .A2(new_n962), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n761), .A2(new_n856), .A3(new_n931), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n931), .B1(new_n761), .B2(new_n856), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1138), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n949), .A2(G330), .A3(new_n856), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n960), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n856), .B1(new_n766), .B2(new_n767), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1144), .A2(new_n962), .A3(new_n1145), .A4(new_n1139), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1142), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n455), .A2(new_n761), .ZN(new_n1148));
  AND3_X1   g0948(.A1(new_n966), .A2(new_n681), .A3(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n946), .A2(new_n957), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n765), .A2(new_n728), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT90), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n765), .A2(KEYINPUT90), .A3(new_n728), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n961), .B1(new_n1157), .B2(new_n856), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1152), .B1(new_n1158), .B2(new_n960), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n954), .A2(new_n955), .B1(new_n963), .B2(new_n958), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1139), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n960), .B1(new_n1145), .B2(new_n962), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1160), .B(new_n1139), .C1(new_n1162), .C2(new_n1151), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1150), .B1(new_n1161), .B2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1160), .B1(new_n1162), .B2(new_n1151), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(new_n1140), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1167), .A2(new_n1163), .A3(new_n1149), .A4(new_n1147), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1165), .A2(new_n740), .A3(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1167), .A2(new_n1026), .A3(new_n1163), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n778), .B1(new_n393), .B2(new_n865), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n813), .A2(new_n459), .B1(new_n871), .B2(new_n807), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1119), .B(new_n1172), .C1(G97), .C2(new_n812), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n365), .B1(new_n834), .B2(new_n818), .C1(new_n819), .C2(new_n202), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(new_n823), .B2(G107), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1173), .B(new_n1175), .C1(new_n820), .C2(new_n799), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(G128), .A2(new_n836), .B1(new_n823), .B2(G137), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n804), .A2(new_n828), .B1(new_n819), .B2(new_n249), .ZN(new_n1178));
  XOR2_X1   g0978(.A(KEYINPUT54), .B(G143), .Z(new_n1179));
  AOI21_X1  g0979(.A(new_n1178), .B1(new_n812), .B2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n365), .B1(new_n808), .B2(G125), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n818), .A2(new_n257), .ZN(new_n1182));
  XOR2_X1   g0982(.A(KEYINPUT111), .B(KEYINPUT53), .Z(new_n1183));
  XNOR2_X1  g0983(.A(new_n1182), .B(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(G132), .B2(new_n814), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n1177), .A2(new_n1180), .A3(new_n1181), .A4(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1176), .A2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1171), .B1(new_n1187), .B2(new_n788), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(new_n956), .B2(new_n786), .ZN(new_n1189));
  AND2_X1   g0989(.A1(new_n1170), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1169), .A2(new_n1190), .ZN(G378));
  INV_X1    g0991(.A(KEYINPUT57), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(new_n1168), .B2(new_n1149), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT114), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n965), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n281), .A2(new_n891), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n313), .B(new_n1196), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1197), .B(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n716), .B1(new_n941), .B2(new_n946), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1199), .B1(new_n940), .B2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n938), .B1(new_n934), .B2(new_n935), .ZN(new_n1202));
  AOI211_X1 g1002(.A(KEYINPUT99), .B(KEYINPUT40), .C1(new_n927), .C2(new_n933), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1199), .B(new_n1200), .C1(new_n1202), .C2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1195), .B1(new_n1201), .B2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1200), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1199), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1209), .A2(new_n965), .A3(new_n1204), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1194), .B1(new_n1206), .B2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n965), .B1(new_n1209), .B2(new_n1204), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1212), .A2(KEYINPUT114), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1193), .B1(new_n1211), .B2(new_n1213), .ZN(new_n1214));
  AND3_X1   g1014(.A1(new_n1209), .A2(new_n965), .A3(new_n1204), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1215), .A2(new_n1212), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n966), .A2(new_n681), .A3(new_n1148), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1161), .A2(new_n1164), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1150), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1217), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1192), .B1(new_n1216), .B2(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1214), .A2(new_n1221), .A3(new_n740), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1206), .A2(new_n1210), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(new_n1026), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n778), .B1(G50), .B2(new_n865), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n814), .A2(G128), .B1(new_n866), .B2(new_n1179), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(new_n1226), .B(KEYINPUT112), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n812), .A2(G137), .B1(new_n805), .B2(G150), .ZN(new_n1228));
  INV_X1    g1028(.A(G125), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n1228), .B1(new_n822), .B2(new_n880), .C1(new_n1229), .C2(new_n799), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1227), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  OR2_X1    g1032(.A1(new_n1232), .A2(KEYINPUT59), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(KEYINPUT59), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n258), .B(new_n483), .C1(new_n819), .C2(new_n828), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(G124), .B2(new_n808), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1233), .A2(new_n1234), .A3(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n808), .A2(G283), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1043), .A2(G58), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  OAI221_X1 g1040(.A(new_n1240), .B1(new_n551), .B2(new_n813), .C1(new_n379), .C2(new_n811), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n823), .A2(G97), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n365), .A2(new_n483), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(new_n866), .B2(G77), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1242), .A2(new_n1032), .A3(new_n1244), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n1241), .B(new_n1245), .C1(G116), .C2(new_n836), .ZN(new_n1246));
  OR2_X1    g1046(.A1(new_n1246), .A2(KEYINPUT58), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(KEYINPUT58), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1243), .B(new_n249), .C1(G33), .C2(G41), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1237), .A2(new_n1247), .A3(new_n1248), .A4(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1225), .B1(new_n1250), .B2(new_n788), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(new_n1208), .B2(new_n786), .ZN(new_n1252));
  XNOR2_X1  g1052(.A(new_n1252), .B(KEYINPUT113), .ZN(new_n1253));
  AND2_X1   g1053(.A1(new_n1224), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1222), .A2(new_n1254), .ZN(G375));
  NAND2_X1  g1055(.A1(new_n1147), .A2(new_n1026), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n551), .A2(new_n811), .B1(new_n813), .B2(new_n820), .ZN(new_n1257));
  AOI211_X1 g1057(.A(new_n1076), .B(new_n1257), .C1(G303), .C2(new_n808), .ZN(new_n1258));
  OAI221_X1 g1058(.A(new_n365), .B1(new_n1079), .B2(new_n818), .C1(new_n819), .C2(new_n226), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(new_n836), .B2(G294), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1258), .B(new_n1260), .C1(new_n459), .C2(new_n822), .ZN(new_n1261));
  XOR2_X1   g1061(.A(new_n1261), .B(KEYINPUT115), .Z(new_n1262));
  AOI21_X1  g1062(.A(new_n365), .B1(new_n866), .B2(G159), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n1239), .B(new_n1263), .C1(new_n799), .C2(new_n880), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(new_n805), .A2(G50), .B1(new_n808), .B2(G128), .ZN(new_n1265));
  OAI221_X1 g1065(.A(new_n1265), .B1(new_n876), .B2(new_n813), .C1(new_n257), .C2(new_n811), .ZN(new_n1266));
  AOI211_X1 g1066(.A(new_n1264), .B(new_n1266), .C1(new_n823), .C2(new_n1179), .ZN(new_n1267));
  OAI21_X1  g1067(.A(KEYINPUT116), .B1(new_n1262), .B2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n788), .ZN(new_n1269));
  NOR3_X1   g1069(.A1(new_n1262), .A2(KEYINPUT116), .A3(new_n1267), .ZN(new_n1270));
  OAI221_X1 g1070(.A(new_n778), .B1(G68), .B2(new_n865), .C1(new_n1269), .C2(new_n1270), .ZN(new_n1271));
  XOR2_X1   g1071(.A(new_n1271), .B(KEYINPUT117), .Z(new_n1272));
  NOR2_X1   g1072(.A1(new_n931), .A2(new_n786), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1256), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1219), .A2(new_n996), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1217), .A2(new_n1142), .A3(new_n1146), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1274), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(G381));
  INV_X1    g1078(.A(G396), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1063), .A2(new_n1279), .A3(new_n1096), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1136), .A2(new_n887), .A3(new_n1281), .ZN(new_n1282));
  NOR3_X1   g1082(.A1(G381), .A2(new_n1282), .A3(G387), .ZN(new_n1283));
  XNOR2_X1  g1083(.A(new_n1283), .B(KEYINPUT118), .ZN(new_n1284));
  AND3_X1   g1084(.A1(new_n1169), .A2(KEYINPUT119), .A3(new_n1190), .ZN(new_n1285));
  AOI21_X1  g1085(.A(KEYINPUT119), .B1(new_n1169), .B2(new_n1190), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1222), .A2(new_n1287), .A3(new_n1254), .ZN(new_n1288));
  OR2_X1    g1088(.A1(new_n1284), .A2(new_n1288), .ZN(G407));
  OAI211_X1 g1089(.A(G407), .B(G213), .C1(G343), .C2(new_n1288), .ZN(G409));
  INV_X1    g1090(.A(KEYINPUT123), .ZN(new_n1291));
  AND3_X1   g1091(.A1(new_n1027), .A2(new_n1136), .A3(new_n1058), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1136), .B1(new_n1027), .B2(new_n1058), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT121), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1279), .B1(new_n1063), .B2(new_n1096), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1295), .B1(new_n1281), .B2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1296), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1298), .A2(KEYINPUT121), .A3(new_n1280), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1297), .A2(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1291), .B1(new_n1294), .B2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(G387), .A2(G390), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1027), .A2(new_n1136), .A3(new_n1058), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  AND2_X1   g1104(.A1(new_n1297), .A2(new_n1299), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1304), .A2(KEYINPUT123), .A3(new_n1305), .ZN(new_n1306));
  OAI21_X1  g1106(.A(KEYINPUT122), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT122), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1294), .A2(new_n1308), .A3(new_n1300), .ZN(new_n1309));
  AOI22_X1  g1109(.A1(new_n1301), .A2(new_n1306), .B1(new_n1307), .B2(new_n1309), .ZN(new_n1310));
  XNOR2_X1  g1110(.A(new_n1310), .B(KEYINPUT126), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n722), .A2(G213), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1222), .A2(G378), .A3(new_n1254), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1026), .B1(new_n1211), .B2(new_n1213), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n996), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1168), .A2(new_n1149), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1223), .A2(new_n1316), .A3(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1315), .A2(new_n1253), .A3(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1319), .A2(new_n1287), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1313), .B1(new_n1314), .B2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1150), .A2(KEYINPUT60), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1322), .A2(new_n1276), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1323), .A2(new_n1128), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1322), .A2(new_n1276), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1274), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1326));
  XNOR2_X1  g1126(.A(new_n1326), .B(new_n887), .ZN(new_n1327));
  AOI21_X1  g1127(.A(KEYINPUT62), .B1(new_n1321), .B2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT125), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1314), .A2(new_n1320), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1329), .B1(new_n1330), .B2(new_n1312), .ZN(new_n1331));
  AOI211_X1 g1131(.A(KEYINPUT125), .B(new_n1313), .C1(new_n1314), .C2(new_n1320), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  AND2_X1   g1133(.A1(new_n1327), .A2(KEYINPUT62), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1328), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  XNOR2_X1  g1135(.A(new_n1326), .B(G384), .ZN(new_n1336));
  INV_X1    g1136(.A(G2897), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1336), .B1(new_n1337), .B2(new_n1312), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(new_n1312), .A2(new_n1337), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1327), .A2(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1338), .A2(new_n1340), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1341), .B1(new_n1331), .B2(new_n1332), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT61), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1342), .A2(new_n1343), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1311), .B1(new_n1335), .B2(new_n1344), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1321), .B1(new_n1338), .B2(new_n1340), .ZN(new_n1346));
  OAI21_X1  g1146(.A(KEYINPUT124), .B1(new_n1310), .B2(KEYINPUT61), .ZN(new_n1347));
  NOR3_X1   g1147(.A1(new_n1294), .A2(new_n1291), .A3(new_n1300), .ZN(new_n1348));
  AOI21_X1  g1148(.A(KEYINPUT123), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1308), .B1(new_n1294), .B2(new_n1300), .ZN(new_n1350));
  AND4_X1   g1150(.A1(new_n1308), .A2(new_n1300), .A3(new_n1302), .A4(new_n1303), .ZN(new_n1351));
  OAI22_X1  g1151(.A1(new_n1348), .A2(new_n1349), .B1(new_n1350), .B2(new_n1351), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT124), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1352), .A2(new_n1353), .A3(new_n1343), .ZN(new_n1354));
  AOI21_X1  g1154(.A(new_n1346), .B1(new_n1347), .B2(new_n1354), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1333), .A2(KEYINPUT63), .A3(new_n1327), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1321), .A2(new_n1327), .ZN(new_n1357));
  XNOR2_X1  g1157(.A(KEYINPUT120), .B(KEYINPUT63), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1357), .A2(new_n1358), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1355), .A2(new_n1356), .A3(new_n1359), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1345), .A2(new_n1360), .ZN(G405));
  AND2_X1   g1161(.A1(G375), .A2(new_n1287), .ZN(new_n1362));
  INV_X1    g1162(.A(new_n1314), .ZN(new_n1363));
  NOR2_X1   g1163(.A1(new_n1362), .A2(new_n1363), .ZN(new_n1364));
  NOR2_X1   g1164(.A1(new_n1364), .A2(new_n1336), .ZN(new_n1365));
  NOR3_X1   g1165(.A1(new_n1362), .A2(new_n1363), .A3(new_n1327), .ZN(new_n1366));
  NOR2_X1   g1166(.A1(new_n1365), .A2(new_n1366), .ZN(new_n1367));
  NAND3_X1  g1167(.A1(new_n1367), .A2(KEYINPUT127), .A3(new_n1352), .ZN(new_n1368));
  OR2_X1    g1168(.A1(new_n1352), .A2(KEYINPUT127), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1352), .A2(KEYINPUT127), .ZN(new_n1370));
  OAI211_X1 g1170(.A(new_n1369), .B(new_n1370), .C1(new_n1365), .C2(new_n1366), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1368), .A2(new_n1371), .ZN(G402));
endmodule


