//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 1 0 1 1 0 0 0 0 0 0 1 1 1 1 1 1 1 0 0 0 1 0 0 1 0 1 0 0 1 1 0 1 1 0 0 0 0 0 1 1 1 0 0 0 1 0 1 1 0 1 0 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n796, new_n797, new_n798, new_n799,
    new_n801, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n907, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n990,
    new_n991, new_n992, new_n994, new_n995, new_n996, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1011, new_n1012, new_n1013,
    new_n1015, new_n1016;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  INV_X1    g001(.A(G113gat), .ZN(new_n203));
  INV_X1    g002(.A(G120gat), .ZN(new_n204));
  AOI21_X1  g003(.A(KEYINPUT1), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(new_n203), .B2(new_n204), .ZN(new_n206));
  INV_X1    g005(.A(G134gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G127gat), .ZN(new_n208));
  INV_X1    g007(.A(G127gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G134gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT70), .ZN(new_n211));
  AND3_X1   g010(.A1(new_n208), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n211), .B1(new_n208), .B2(new_n210), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n206), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G127gat), .B(G134gat), .ZN(new_n215));
  XNOR2_X1  g014(.A(KEYINPUT71), .B(G113gat), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n205), .B(new_n215), .C1(new_n216), .C2(new_n204), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT23), .ZN(new_n220));
  NAND2_X1  g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT23), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n222), .B1(G169gat), .B2(G176gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n220), .A2(new_n221), .A3(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G183gat), .A2(G190gat), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n220), .A2(new_n228), .A3(new_n223), .A4(new_n221), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT65), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n220), .A2(new_n230), .A3(new_n223), .A4(new_n221), .ZN(new_n231));
  AND3_X1   g030(.A1(new_n229), .A2(new_n231), .A3(KEYINPUT25), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n229), .B1(KEYINPUT25), .B2(new_n231), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n227), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  AND3_X1   g033(.A1(new_n220), .A2(new_n221), .A3(new_n223), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT25), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n235), .B(new_n228), .C1(new_n230), .C2(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n229), .A2(new_n231), .A3(KEYINPUT25), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n237), .A2(new_n226), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n234), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(KEYINPUT66), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n234), .A2(new_n242), .A3(new_n239), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n245));
  INV_X1    g044(.A(G183gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(KEYINPUT27), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT27), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(G183gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(KEYINPUT67), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT67), .ZN(new_n252));
  AOI21_X1  g051(.A(G190gat), .B1(new_n247), .B2(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT28), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT28), .ZN(new_n255));
  NOR3_X1   g054(.A1(new_n250), .A2(new_n255), .A3(G190gat), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n245), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT27), .B(G183gat), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n258), .A2(new_n252), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n247), .A2(new_n252), .ZN(new_n260));
  INV_X1    g059(.A(G190gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n255), .B1(new_n259), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n256), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n263), .A2(new_n264), .A3(KEYINPUT68), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n257), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n267));
  OR3_X1    g066(.A1(new_n267), .A2(new_n219), .A3(KEYINPUT69), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT69), .B1(new_n267), .B2(new_n219), .ZN(new_n269));
  INV_X1    g068(.A(G169gat), .ZN(new_n270));
  INV_X1    g069(.A(G176gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OAI211_X1 g071(.A(new_n268), .B(new_n269), .C1(KEYINPUT26), .C2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(new_n228), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n266), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n218), .B1(new_n244), .B2(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n274), .B1(new_n257), .B2(new_n265), .ZN(new_n278));
  INV_X1    g077(.A(new_n218), .ZN(new_n279));
  AOI211_X1 g078(.A(new_n278), .B(new_n279), .C1(new_n241), .C2(new_n243), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(G227gat), .A2(G233gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n282), .B(KEYINPUT64), .ZN(new_n283));
  OAI21_X1  g082(.A(KEYINPUT34), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n278), .B1(new_n241), .B2(new_n243), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(new_n218), .ZN(new_n286));
  AND3_X1   g085(.A1(new_n234), .A2(new_n242), .A3(new_n239), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n242), .B1(new_n234), .B2(new_n239), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n276), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(new_n279), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT34), .ZN(new_n292));
  INV_X1    g091(.A(new_n283), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT33), .B1(new_n281), .B2(new_n283), .ZN(new_n295));
  XNOR2_X1  g094(.A(G15gat), .B(G43gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(G71gat), .B(G99gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n296), .B(new_n297), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n284), .B(new_n294), .C1(new_n295), .C2(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n286), .A2(new_n290), .A3(new_n283), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT32), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT33), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n298), .B1(new_n300), .B2(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n292), .B1(new_n291), .B2(new_n293), .ZN(new_n305));
  AOI211_X1 g104(.A(KEYINPUT34), .B(new_n283), .C1(new_n286), .C2(new_n290), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AND3_X1   g106(.A1(new_n299), .A2(new_n302), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n302), .B1(new_n299), .B2(new_n307), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n202), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(KEYINPUT73), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT73), .ZN(new_n312));
  OAI211_X1 g111(.A(new_n312), .B(new_n202), .C1(new_n308), .C2(new_n309), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n299), .A2(new_n307), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(new_n301), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n299), .A2(new_n302), .A3(new_n307), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n316), .A2(KEYINPUT36), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT72), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT72), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n316), .A2(new_n320), .A3(KEYINPUT36), .A4(new_n317), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n314), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(G228gat), .ZN(new_n324));
  INV_X1    g123(.A(G233gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT81), .ZN(new_n327));
  INV_X1    g126(.A(G141gat), .ZN(new_n328));
  INV_X1    g127(.A(G148gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT2), .ZN(new_n331));
  NAND2_X1  g130(.A1(G141gat), .A2(G148gat), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT79), .ZN(new_n334));
  INV_X1    g133(.A(G155gat), .ZN(new_n335));
  INV_X1    g134(.A(G162gat), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(G155gat), .A2(G162gat), .ZN(new_n338));
  OAI21_X1  g137(.A(KEYINPUT79), .B1(G155gat), .B2(G162gat), .ZN(new_n339));
  AND4_X1   g138(.A1(new_n333), .A2(new_n337), .A3(new_n338), .A4(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n331), .A2(new_n335), .A3(new_n336), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(new_n338), .ZN(new_n342));
  AND2_X1   g141(.A1(G141gat), .A2(G148gat), .ZN(new_n343));
  NOR2_X1   g142(.A1(G141gat), .A2(G148gat), .ZN(new_n344));
  OAI21_X1  g143(.A(KEYINPUT80), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT80), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n330), .A2(new_n346), .A3(new_n332), .ZN(new_n347));
  AND3_X1   g146(.A1(new_n342), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n327), .B1(new_n340), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n330), .A2(new_n332), .ZN(new_n350));
  AOI22_X1  g149(.A1(new_n350), .A2(KEYINPUT80), .B1(new_n341), .B2(new_n338), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(new_n347), .ZN(new_n352));
  AND3_X1   g151(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(new_n333), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n352), .A2(new_n354), .A3(KEYINPUT81), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n349), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(G197gat), .B(G204gat), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT22), .ZN(new_n358));
  INV_X1    g157(.A(G211gat), .ZN(new_n359));
  INV_X1    g158(.A(G218gat), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n357), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  XOR2_X1   g162(.A(G211gat), .B(G218gat), .Z(new_n364));
  INV_X1    g163(.A(KEYINPUT74), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n363), .B(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT29), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT3), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n366), .B(new_n362), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n370), .B(KEYINPUT75), .ZN(new_n371));
  AOI22_X1  g170(.A1(new_n351), .A2(new_n347), .B1(new_n353), .B2(new_n333), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT3), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT29), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  OAI221_X1 g173(.A(new_n326), .B1(new_n356), .B2(new_n369), .C1(new_n371), .C2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(G22gat), .ZN(new_n376));
  OR2_X1    g175(.A1(new_n363), .A2(new_n364), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n363), .A2(new_n364), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n377), .A2(new_n368), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n372), .B1(new_n379), .B2(new_n373), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n374), .A2(new_n367), .ZN(new_n381));
  OAI22_X1  g180(.A1(new_n380), .A2(new_n381), .B1(new_n324), .B2(new_n325), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n375), .A2(new_n376), .A3(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n376), .B1(new_n375), .B2(new_n382), .ZN(new_n385));
  OAI21_X1  g184(.A(G78gat), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n385), .ZN(new_n387));
  INV_X1    g186(.A(G78gat), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n387), .A2(new_n388), .A3(new_n383), .ZN(new_n389));
  XNOR2_X1  g188(.A(KEYINPUT31), .B(G50gat), .ZN(new_n390));
  INV_X1    g189(.A(G106gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n390), .B(new_n391), .ZN(new_n392));
  AND3_X1   g191(.A1(new_n386), .A2(new_n389), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n392), .B1(new_n386), .B2(new_n389), .ZN(new_n394));
  OR2_X1    g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(G226gat), .A2(G233gat), .ZN(new_n396));
  XOR2_X1   g195(.A(new_n396), .B(KEYINPUT76), .Z(new_n397));
  OAI21_X1  g196(.A(new_n397), .B1(new_n285), .B2(KEYINPUT29), .ZN(new_n398));
  AND2_X1   g197(.A1(new_n234), .A2(new_n239), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(new_n276), .ZN(new_n400));
  INV_X1    g199(.A(new_n396), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n371), .B1(new_n398), .B2(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n397), .B1(new_n244), .B2(new_n276), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n401), .B1(new_n400), .B2(new_n368), .ZN(new_n405));
  NOR3_X1   g204(.A1(new_n404), .A2(new_n405), .A3(new_n370), .ZN(new_n406));
  OAI21_X1  g205(.A(KEYINPUT77), .B1(new_n403), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT29), .B1(new_n399), .B2(new_n276), .ZN(new_n408));
  OAI221_X1 g207(.A(new_n367), .B1(new_n408), .B2(new_n401), .C1(new_n285), .C2(new_n397), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT77), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n289), .A2(new_n368), .ZN(new_n411));
  AOI22_X1  g210(.A1(new_n411), .A2(new_n397), .B1(new_n401), .B2(new_n400), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n409), .B(new_n410), .C1(new_n412), .C2(new_n371), .ZN(new_n413));
  XOR2_X1   g212(.A(G8gat), .B(G36gat), .Z(new_n414));
  XNOR2_X1  g213(.A(new_n414), .B(KEYINPUT78), .ZN(new_n415));
  XNOR2_X1  g214(.A(G64gat), .B(G92gat), .ZN(new_n416));
  XOR2_X1   g215(.A(new_n415), .B(new_n416), .Z(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n407), .A2(new_n413), .A3(new_n418), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n409), .B(new_n417), .C1(new_n412), .C2(new_n371), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT30), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n403), .A2(new_n406), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n423), .A2(KEYINPUT30), .A3(new_n417), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n419), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT82), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n352), .A2(new_n354), .A3(new_n214), .A4(new_n217), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n426), .B1(new_n427), .B2(KEYINPUT4), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT4), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n279), .A2(KEYINPUT82), .A3(new_n429), .A4(new_n372), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n427), .A2(KEYINPUT4), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n428), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(G225gat), .A2(G233gat), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n349), .A2(new_n355), .A3(KEYINPUT3), .ZN(new_n435));
  AOI22_X1  g234(.A1(new_n372), .A2(new_n373), .B1(new_n214), .B2(new_n217), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n432), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT5), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n349), .A2(new_n355), .A3(new_n218), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n427), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n439), .B1(new_n441), .B2(new_n434), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n279), .A2(new_n429), .A3(new_n372), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n431), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n437), .A2(new_n439), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  XOR2_X1   g246(.A(G1gat), .B(G29gat), .Z(new_n448));
  XNOR2_X1  g247(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n448), .B(new_n449), .ZN(new_n450));
  XNOR2_X1  g249(.A(G57gat), .B(G85gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n450), .B(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n447), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT6), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n443), .A2(KEYINPUT84), .A3(new_n452), .A4(new_n446), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n457), .A2(new_n455), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n443), .A2(new_n452), .A3(new_n446), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT84), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AND2_X1   g260(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n454), .B(KEYINPUT85), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n456), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n395), .B1(new_n425), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT38), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n407), .A2(KEYINPUT37), .A3(new_n413), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT37), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n417), .B1(new_n423), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n466), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  OAI22_X1  g269(.A1(new_n285), .A2(new_n397), .B1(new_n408), .B2(new_n401), .ZN(new_n471));
  AOI22_X1  g270(.A1(new_n412), .A2(new_n371), .B1(new_n370), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n466), .B1(new_n472), .B2(new_n468), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n409), .B1(new_n412), .B2(new_n371), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n418), .B1(new_n474), .B2(KEYINPUT37), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n420), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n461), .A2(new_n454), .A3(new_n455), .A4(new_n457), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT87), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT87), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n458), .A2(new_n479), .A3(new_n454), .A4(new_n461), .ZN(new_n480));
  INV_X1    g279(.A(new_n456), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n478), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NOR3_X1   g281(.A1(new_n470), .A2(new_n476), .A3(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT86), .ZN(new_n484));
  AOI22_X1  g283(.A1(new_n444), .A2(new_n431), .B1(new_n435), .B2(new_n436), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n484), .B1(new_n485), .B2(new_n433), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n435), .A2(new_n436), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n445), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n488), .A2(KEYINPUT86), .A3(new_n434), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT39), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n440), .A2(new_n433), .A3(new_n427), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n486), .A2(new_n489), .A3(KEYINPUT39), .A4(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n492), .A2(new_n452), .A3(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT40), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n492), .A2(KEYINPUT40), .A3(new_n452), .A4(new_n494), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n497), .A2(new_n454), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n425), .A2(new_n499), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n393), .A2(new_n394), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n465), .B1(new_n483), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n323), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n308), .A2(new_n309), .ZN(new_n506));
  INV_X1    g305(.A(new_n425), .ZN(new_n507));
  INV_X1    g306(.A(new_n464), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n506), .A2(new_n507), .A3(new_n508), .A4(new_n501), .ZN(new_n509));
  AND4_X1   g308(.A1(new_n507), .A2(new_n501), .A3(new_n316), .A4(new_n317), .ZN(new_n510));
  INV_X1    g309(.A(new_n482), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n511), .A2(KEYINPUT35), .ZN(new_n512));
  AOI22_X1  g311(.A1(new_n509), .A2(KEYINPUT35), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(KEYINPUT88), .B1(new_n505), .B2(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n503), .B1(new_n322), .B2(new_n314), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT88), .ZN(new_n517));
  NOR3_X1   g316(.A1(new_n516), .A2(new_n517), .A3(new_n513), .ZN(new_n518));
  OR2_X1    g317(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(G29gat), .ZN(new_n520));
  INV_X1    g319(.A(G36gat), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n520), .A2(new_n521), .A3(KEYINPUT14), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT14), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n523), .B1(G29gat), .B2(G36gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(G29gat), .A2(G36gat), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n522), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT15), .ZN(new_n527));
  OR2_X1    g326(.A1(G43gat), .A2(G50gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(G43gat), .A2(G50gat), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n528), .A2(new_n527), .A3(new_n529), .ZN(new_n532));
  AND2_X1   g331(.A1(G43gat), .A2(G50gat), .ZN(new_n533));
  NOR2_X1   g332(.A1(G43gat), .A2(G50gat), .ZN(new_n534));
  OAI21_X1  g333(.A(KEYINPUT15), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n531), .B(KEYINPUT90), .C1(new_n536), .C2(new_n526), .ZN(new_n537));
  INV_X1    g336(.A(new_n526), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT90), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n538), .A2(new_n539), .A3(new_n535), .A4(new_n532), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT93), .ZN(new_n543));
  XNOR2_X1  g342(.A(G15gat), .B(G22gat), .ZN(new_n544));
  INV_X1    g343(.A(G1gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(KEYINPUT16), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n544), .A2(G1gat), .ZN(new_n549));
  NOR3_X1   g348(.A1(new_n548), .A2(new_n549), .A3(G8gat), .ZN(new_n550));
  INV_X1    g349(.A(G8gat), .ZN(new_n551));
  OR2_X1    g350(.A1(new_n544), .A2(G1gat), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n551), .B1(new_n552), .B2(new_n547), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n543), .B1(new_n550), .B2(new_n553), .ZN(new_n554));
  OAI21_X1  g353(.A(G8gat), .B1(new_n548), .B2(new_n549), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n552), .A2(new_n551), .A3(new_n547), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n555), .A2(new_n556), .A3(KEYINPUT93), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n542), .A2(new_n554), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(G229gat), .A2(G233gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(KEYINPUT92), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n541), .A2(KEYINPUT17), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n550), .A2(new_n553), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT17), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n537), .A2(new_n565), .A3(new_n540), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n563), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT91), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n563), .A2(KEYINPUT91), .A3(new_n564), .A4(new_n566), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n562), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n554), .A2(new_n557), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(new_n541), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(new_n558), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n560), .B(KEYINPUT13), .ZN(new_n575));
  AOI22_X1  g374(.A1(new_n571), .A2(KEYINPUT18), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT18), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT94), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n577), .B1(new_n571), .B2(new_n578), .ZN(new_n579));
  AOI211_X1 g378(.A(KEYINPUT94), .B(new_n562), .C1(new_n569), .C2(new_n570), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n576), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  AND2_X1   g380(.A1(new_n558), .A2(new_n561), .ZN(new_n582));
  AND3_X1   g381(.A1(new_n537), .A2(new_n565), .A3(new_n540), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n565), .B1(new_n537), .B2(new_n540), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(KEYINPUT91), .B1(new_n585), .B2(new_n564), .ZN(new_n586));
  INV_X1    g385(.A(new_n570), .ZN(new_n587));
  OAI211_X1 g386(.A(KEYINPUT18), .B(new_n582), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT95), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n575), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G113gat), .B(G141gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(G197gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(KEYINPUT11), .B(G169gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(KEYINPUT89), .B(KEYINPUT12), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n581), .A2(new_n591), .A3(new_n598), .ZN(new_n599));
  OAI221_X1 g398(.A(new_n576), .B1(new_n589), .B2(new_n597), .C1(new_n579), .C2(new_n580), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AND2_X1   g400(.A1(new_n519), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(G71gat), .A2(G78gat), .ZN(new_n603));
  OR2_X1    g402(.A1(G71gat), .A2(G78gat), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT9), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(G64gat), .ZN(new_n607));
  OAI21_X1  g406(.A(KEYINPUT96), .B1(new_n607), .B2(G57gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(G57gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NOR3_X1   g409(.A1(new_n607), .A2(KEYINPUT96), .A3(G57gat), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n606), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(G57gat), .B(G64gat), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n603), .B(new_n604), .C1(new_n613), .C2(new_n605), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT21), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(G231gat), .A2(G233gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  OR2_X1    g418(.A1(new_n619), .A2(new_n209), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n209), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n572), .B1(new_n616), .B2(new_n615), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n620), .A2(new_n623), .A3(new_n621), .ZN(new_n626));
  XNOR2_X1  g425(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(KEYINPUT97), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(G155gat), .ZN(new_n629));
  XOR2_X1   g428(.A(G183gat), .B(G211gat), .Z(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  AND3_X1   g430(.A1(new_n625), .A2(new_n626), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n631), .B1(new_n625), .B2(new_n626), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT100), .ZN(new_n635));
  NAND2_X1  g434(.A1(G85gat), .A2(G92gat), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT98), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n638), .A2(KEYINPUT7), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT7), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n640), .A2(KEYINPUT98), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n637), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(KEYINPUT98), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n638), .A2(KEYINPUT7), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n643), .A2(new_n644), .A3(new_n636), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(G99gat), .B(G106gat), .ZN(new_n647));
  AND2_X1   g446(.A1(KEYINPUT99), .A2(G85gat), .ZN(new_n648));
  NOR2_X1   g447(.A1(KEYINPUT99), .A2(G85gat), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(G92gat), .ZN(new_n651));
  NAND2_X1  g450(.A1(G99gat), .A2(G106gat), .ZN(new_n652));
  AOI22_X1  g451(.A1(new_n650), .A2(new_n651), .B1(KEYINPUT8), .B2(new_n652), .ZN(new_n653));
  AND3_X1   g452(.A1(new_n646), .A2(new_n647), .A3(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n647), .B1(new_n646), .B2(new_n653), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n635), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n647), .ZN(new_n657));
  AND3_X1   g456(.A1(new_n643), .A2(new_n644), .A3(new_n636), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n636), .B1(new_n643), .B2(new_n644), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n652), .A2(KEYINPUT8), .ZN(new_n661));
  XNOR2_X1  g460(.A(KEYINPUT99), .B(G85gat), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n661), .B1(new_n662), .B2(G92gat), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n657), .B1(new_n660), .B2(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n646), .A2(new_n647), .A3(new_n653), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n664), .A2(KEYINPUT100), .A3(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n656), .A2(new_n542), .A3(new_n666), .ZN(new_n667));
  AND2_X1   g466(.A1(G232gat), .A2(G233gat), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(KEYINPUT41), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n656), .A2(new_n666), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n671), .A2(new_n563), .A3(new_n566), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g472(.A(G190gat), .B(G218gat), .Z(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n674), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n670), .A2(new_n676), .A3(new_n672), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n668), .A2(KEYINPUT41), .ZN(new_n678));
  XNOR2_X1  g477(.A(G134gat), .B(G162gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n675), .A2(new_n677), .A3(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n680), .B1(new_n675), .B2(new_n677), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n634), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(G230gat), .A2(G233gat), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  OR2_X1    g485(.A1(new_n647), .A2(KEYINPUT101), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n612), .A2(new_n614), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n688), .B1(new_n654), .B2(new_n655), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n612), .A2(new_n614), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n664), .A2(new_n690), .A3(new_n665), .A4(new_n687), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT10), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n689), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n615), .A2(new_n692), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n656), .A2(new_n666), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n686), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT102), .ZN(new_n698));
  XNOR2_X1  g497(.A(G120gat), .B(G148gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(G176gat), .B(G204gat), .ZN(new_n700));
  XOR2_X1   g499(.A(new_n699), .B(new_n700), .Z(new_n701));
  NAND2_X1  g500(.A1(new_n689), .A2(new_n691), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(new_n686), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n697), .A2(new_n698), .A3(new_n701), .A4(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n701), .ZN(new_n705));
  OAI21_X1  g504(.A(KEYINPUT102), .B1(new_n705), .B2(new_n696), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n701), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n685), .B(KEYINPUT103), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n709), .B1(new_n693), .B2(new_n695), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n685), .B1(new_n689), .B2(new_n691), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n708), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n707), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n684), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  OR2_X1    g515(.A1(new_n464), .A2(KEYINPUT104), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n464), .A2(KEYINPUT104), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n602), .A2(new_n716), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(G1gat), .ZN(G1324gat));
  AND3_X1   g521(.A1(new_n602), .A2(new_n425), .A3(new_n716), .ZN(new_n723));
  OR2_X1    g522(.A1(new_n723), .A2(new_n551), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT42), .ZN(new_n725));
  XOR2_X1   g524(.A(KEYINPUT16), .B(G8gat), .Z(new_n726));
  AOI21_X1  g525(.A(new_n725), .B1(new_n723), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(KEYINPUT105), .A2(KEYINPUT42), .ZN(new_n728));
  MUX2_X1   g527(.A(KEYINPUT105), .B(new_n728), .S(new_n726), .Z(new_n729));
  AOI22_X1  g528(.A1(new_n724), .A2(new_n727), .B1(new_n723), .B2(new_n729), .ZN(G1325gat));
  NAND2_X1  g529(.A1(new_n602), .A2(new_n716), .ZN(new_n731));
  OAI21_X1  g530(.A(G15gat), .B1(new_n731), .B2(new_n323), .ZN(new_n732));
  INV_X1    g531(.A(new_n506), .ZN(new_n733));
  OR2_X1    g532(.A1(new_n733), .A2(G15gat), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n732), .B1(new_n731), .B2(new_n734), .ZN(G1326gat));
  NOR2_X1   g534(.A1(new_n731), .A2(new_n501), .ZN(new_n736));
  XOR2_X1   g535(.A(KEYINPUT43), .B(G22gat), .Z(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(G1327gat));
  NAND3_X1  g537(.A1(new_n601), .A2(new_n634), .A3(new_n714), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n719), .A2(G29gat), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n519), .A2(new_n683), .A3(new_n740), .A4(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT45), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n742), .B(new_n743), .ZN(new_n744));
  OAI211_X1 g543(.A(KEYINPUT44), .B(new_n683), .C1(new_n515), .C2(new_n518), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n505), .A2(new_n514), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n683), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT44), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n745), .A2(new_n740), .A3(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n750), .A2(new_n719), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n751), .A2(new_n520), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT106), .ZN(new_n753));
  OR3_X1    g552(.A1(new_n744), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n753), .B1(new_n744), .B2(new_n752), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(G1328gat));
  NAND3_X1  g555(.A1(new_n519), .A2(new_n683), .A3(new_n740), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n757), .A2(G36gat), .A3(new_n507), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT46), .ZN(new_n759));
  OR2_X1    g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(G36gat), .B1(new_n750), .B2(new_n507), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n758), .A2(new_n759), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(G1329gat));
  INV_X1    g562(.A(new_n323), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n745), .A2(new_n749), .A3(new_n764), .A4(new_n740), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(G43gat), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n733), .A2(G43gat), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n766), .B1(new_n757), .B2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT47), .ZN(new_n770));
  AND3_X1   g569(.A1(new_n769), .A2(KEYINPUT107), .A3(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(KEYINPUT107), .B1(new_n769), .B2(new_n770), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n769), .A2(KEYINPUT108), .A3(new_n770), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT108), .ZN(new_n774));
  INV_X1    g573(.A(new_n757), .ZN(new_n775));
  AOI22_X1  g574(.A1(new_n775), .A2(new_n767), .B1(new_n765), .B2(G43gat), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n774), .B1(new_n776), .B2(KEYINPUT47), .ZN(new_n777));
  OAI22_X1  g576(.A1(new_n771), .A2(new_n772), .B1(new_n773), .B2(new_n777), .ZN(G1330gat));
  OAI21_X1  g577(.A(G50gat), .B1(new_n750), .B2(new_n501), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n501), .A2(G50gat), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n775), .A2(new_n780), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n779), .B(new_n781), .C1(KEYINPUT109), .C2(KEYINPUT48), .ZN(new_n782));
  NAND2_X1  g581(.A1(KEYINPUT109), .A2(KEYINPUT48), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n782), .B(new_n783), .ZN(G1331gat));
  NAND2_X1  g583(.A1(new_n591), .A2(new_n598), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n581), .B(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n786), .A2(new_n684), .A3(new_n713), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n787), .B1(new_n505), .B2(new_n514), .ZN(new_n788));
  XOR2_X1   g587(.A(new_n719), .B(KEYINPUT110), .Z(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g590(.A1(new_n788), .A2(new_n425), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n792), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n793));
  XOR2_X1   g592(.A(KEYINPUT49), .B(G64gat), .Z(new_n794));
  OAI21_X1  g593(.A(new_n793), .B1(new_n792), .B2(new_n794), .ZN(G1333gat));
  NAND3_X1  g594(.A1(new_n788), .A2(G71gat), .A3(new_n764), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT111), .ZN(new_n797));
  AOI21_X1  g596(.A(G71gat), .B1(new_n788), .B2(new_n506), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  XOR2_X1   g598(.A(new_n799), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g599(.A1(new_n788), .A2(new_n395), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(G78gat), .ZN(G1335gat));
  INV_X1    g601(.A(new_n634), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n601), .A2(new_n803), .A3(new_n714), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n745), .A2(new_n749), .A3(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT112), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n745), .A2(new_n749), .A3(KEYINPUT112), .A4(new_n804), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n807), .A2(new_n720), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n662), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n601), .A2(new_n803), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n746), .A2(KEYINPUT51), .A3(new_n683), .A4(new_n811), .ZN(new_n812));
  OR2_X1    g611(.A1(new_n812), .A2(KEYINPUT113), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(KEYINPUT113), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n683), .B(new_n811), .C1(new_n516), .C2(new_n513), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT51), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n813), .A2(new_n814), .A3(new_n817), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n818), .A2(new_n650), .A3(new_n713), .A4(new_n720), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n810), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(KEYINPUT114), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT114), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n810), .A2(new_n822), .A3(new_n819), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(G1336gat));
  NOR3_X1   g623(.A1(new_n507), .A2(G92gat), .A3(new_n714), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n818), .A2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT52), .ZN(new_n827));
  OAI21_X1  g626(.A(G92gat), .B1(new_n805), .B2(new_n507), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n812), .A2(new_n817), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n825), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n831), .B(KEYINPUT115), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n807), .A2(new_n425), .A3(new_n808), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n832), .B1(G92gat), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n829), .B1(new_n834), .B2(new_n827), .ZN(G1337gat));
  NAND3_X1  g634(.A1(new_n807), .A2(new_n764), .A3(new_n808), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT116), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(G99gat), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n836), .A2(new_n837), .ZN(new_n840));
  INV_X1    g639(.A(new_n818), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n733), .A2(G99gat), .A3(new_n714), .ZN(new_n842));
  XOR2_X1   g641(.A(new_n842), .B(KEYINPUT117), .Z(new_n843));
  OAI22_X1  g642(.A1(new_n839), .A2(new_n840), .B1(new_n841), .B2(new_n843), .ZN(G1338gat));
  OAI21_X1  g643(.A(G106gat), .B1(new_n805), .B2(new_n501), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n395), .A2(new_n391), .A3(new_n713), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n845), .B(new_n846), .C1(new_n841), .C2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n807), .A2(new_n395), .A3(new_n808), .ZN(new_n849));
  INV_X1    g648(.A(new_n847), .ZN(new_n850));
  AOI22_X1  g649(.A1(new_n849), .A2(G106gat), .B1(new_n830), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n848), .B1(new_n851), .B2(new_n846), .ZN(G1339gat));
  NOR2_X1   g651(.A1(new_n715), .A2(new_n601), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(new_n595), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n569), .A2(new_n570), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n561), .B1(new_n856), .B2(new_n558), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n574), .A2(new_n575), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n855), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n576), .B(new_n597), .C1(new_n579), .C2(new_n580), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n683), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n693), .A2(new_n695), .ZN(new_n862));
  INV_X1    g661(.A(new_n709), .ZN(new_n863));
  OAI211_X1 g662(.A(new_n697), .B(KEYINPUT54), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n865));
  AOI211_X1 g664(.A(KEYINPUT118), .B(new_n701), .C1(new_n710), .C2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT118), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n862), .A2(new_n865), .A3(new_n863), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n867), .B1(new_n868), .B2(new_n708), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n864), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT55), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OAI211_X1 g671(.A(KEYINPUT55), .B(new_n864), .C1(new_n866), .C2(new_n869), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n872), .A2(new_n707), .A3(new_n873), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n861), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n860), .A2(new_n713), .A3(new_n859), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n876), .B1(new_n786), .B2(new_n874), .ZN(new_n877));
  INV_X1    g676(.A(new_n683), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n875), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n854), .B1(new_n879), .B2(new_n803), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(KEYINPUT119), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n873), .A2(new_n707), .ZN(new_n882));
  AOI211_X1 g681(.A(KEYINPUT54), .B(new_n709), .C1(new_n693), .C2(new_n695), .ZN(new_n883));
  OAI21_X1  g682(.A(KEYINPUT118), .B1(new_n883), .B2(new_n701), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n868), .A2(new_n867), .A3(new_n708), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(KEYINPUT55), .B1(new_n886), .B2(new_n864), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n882), .A2(new_n887), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n888), .A2(new_n683), .A3(new_n859), .A4(new_n860), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n860), .A2(new_n713), .A3(new_n859), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n890), .B1(new_n888), .B2(new_n601), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n889), .B1(new_n891), .B2(new_n683), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n853), .B1(new_n892), .B2(new_n634), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT119), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n395), .B1(new_n881), .B2(new_n895), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n896), .A2(new_n507), .A3(new_n506), .A4(new_n720), .ZN(new_n897));
  OAI21_X1  g696(.A(G113gat), .B1(new_n897), .B2(new_n786), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n881), .A2(new_n895), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n899), .A2(new_n789), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n510), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n601), .A2(new_n216), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n898), .B1(new_n901), .B2(new_n902), .ZN(G1340gat));
  NOR3_X1   g702(.A1(new_n897), .A2(new_n204), .A3(new_n714), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n900), .A2(new_n510), .A3(new_n713), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n904), .B1(new_n905), .B2(new_n204), .ZN(G1341gat));
  OAI21_X1  g705(.A(G127gat), .B1(new_n897), .B2(new_n634), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n803), .A2(new_n209), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n907), .B1(new_n901), .B2(new_n908), .ZN(G1342gat));
  NOR3_X1   g708(.A1(new_n901), .A2(G134gat), .A3(new_n878), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT56), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT120), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n910), .A2(new_n911), .ZN(new_n914));
  OAI21_X1  g713(.A(G134gat), .B1(new_n897), .B2(new_n878), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(G1343gat));
  NOR3_X1   g715(.A1(new_n764), .A2(new_n425), .A3(new_n719), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n892), .A2(new_n634), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n894), .B1(new_n918), .B2(new_n854), .ZN(new_n919));
  AOI211_X1 g718(.A(KEYINPUT119), .B(new_n853), .C1(new_n892), .C2(new_n634), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n395), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT57), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n921), .A2(KEYINPUT121), .A3(new_n922), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n880), .A2(KEYINPUT57), .A3(new_n395), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(KEYINPUT121), .B1(new_n921), .B2(new_n922), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n917), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(G141gat), .B1(new_n927), .B2(new_n786), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT58), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n764), .A2(new_n501), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n900), .A2(new_n930), .ZN(new_n931));
  OR2_X1    g730(.A1(new_n931), .A2(KEYINPUT123), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(KEYINPUT123), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n932), .A2(new_n507), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n601), .A2(new_n328), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n928), .B(new_n929), .C1(new_n934), .C2(new_n935), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n931), .A2(new_n425), .A3(new_n935), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT121), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n501), .B1(new_n881), .B2(new_n895), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n938), .B1(new_n939), .B2(KEYINPUT57), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n940), .A2(new_n924), .A3(new_n923), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT122), .ZN(new_n942));
  AND3_X1   g741(.A1(new_n941), .A2(new_n942), .A3(new_n917), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n942), .B1(new_n941), .B2(new_n917), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(new_n601), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n937), .B1(new_n946), .B2(G141gat), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n936), .B1(new_n947), .B2(new_n929), .ZN(G1344gat));
  OAI21_X1  g747(.A(new_n922), .B1(new_n893), .B2(new_n501), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n949), .B1(new_n921), .B2(new_n922), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n950), .A2(new_n713), .A3(new_n917), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(G148gat), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n952), .A2(KEYINPUT59), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n943), .A2(new_n944), .A3(new_n714), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n329), .A2(KEYINPUT59), .ZN(new_n956));
  INV_X1    g755(.A(new_n956), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n954), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT124), .ZN(new_n959));
  NOR3_X1   g758(.A1(new_n934), .A2(G148gat), .A3(new_n714), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n958), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n927), .A2(KEYINPUT122), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n941), .A2(new_n942), .A3(new_n917), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n963), .A2(new_n713), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n953), .B1(new_n965), .B2(new_n956), .ZN(new_n966));
  OAI21_X1  g765(.A(KEYINPUT124), .B1(new_n966), .B2(new_n960), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n962), .A2(new_n967), .ZN(G1345gat));
  OAI21_X1  g767(.A(new_n335), .B1(new_n934), .B2(new_n634), .ZN(new_n969));
  NAND4_X1  g768(.A1(new_n963), .A2(G155gat), .A3(new_n803), .A4(new_n964), .ZN(new_n970));
  AND3_X1   g769(.A1(new_n969), .A2(KEYINPUT125), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g770(.A(KEYINPUT125), .B1(new_n969), .B2(new_n970), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n971), .A2(new_n972), .ZN(G1346gat));
  INV_X1    g772(.A(new_n934), .ZN(new_n974));
  AOI21_X1  g773(.A(G162gat), .B1(new_n974), .B2(new_n683), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n878), .A2(new_n336), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n975), .B1(new_n945), .B2(new_n976), .ZN(G1347gat));
  OR2_X1    g776(.A1(new_n789), .A2(new_n507), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n978), .A2(new_n733), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(new_n896), .ZN(new_n980));
  OAI21_X1  g779(.A(G169gat), .B1(new_n980), .B2(new_n786), .ZN(new_n981));
  XNOR2_X1  g780(.A(new_n981), .B(KEYINPUT126), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n720), .B1(new_n881), .B2(new_n895), .ZN(new_n983));
  AND4_X1   g782(.A1(new_n425), .A2(new_n983), .A3(new_n501), .A4(new_n506), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n984), .A2(new_n270), .A3(new_n601), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n982), .A2(new_n985), .ZN(G1348gat));
  OAI21_X1  g785(.A(G176gat), .B1(new_n980), .B2(new_n714), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n984), .A2(new_n271), .A3(new_n713), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n987), .A2(new_n988), .ZN(G1349gat));
  OAI21_X1  g788(.A(G183gat), .B1(new_n980), .B2(new_n634), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n984), .A2(new_n258), .A3(new_n803), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  XNOR2_X1  g791(.A(new_n992), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g792(.A(G190gat), .B1(new_n980), .B2(new_n878), .ZN(new_n994));
  XNOR2_X1  g793(.A(new_n994), .B(KEYINPUT61), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n984), .A2(new_n261), .A3(new_n683), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n995), .A2(new_n996), .ZN(G1351gat));
  AND3_X1   g796(.A1(new_n930), .A2(new_n983), .A3(new_n425), .ZN(new_n998));
  AOI21_X1  g797(.A(G197gat), .B1(new_n998), .B2(new_n601), .ZN(new_n999));
  NOR2_X1   g798(.A1(new_n978), .A2(new_n764), .ZN(new_n1000));
  AND2_X1   g799(.A1(new_n1000), .A2(new_n950), .ZN(new_n1001));
  AND2_X1   g800(.A1(new_n601), .A2(G197gat), .ZN(new_n1002));
  AOI21_X1  g801(.A(new_n999), .B1(new_n1001), .B2(new_n1002), .ZN(G1352gat));
  INV_X1    g802(.A(G204gat), .ZN(new_n1004));
  NAND3_X1  g803(.A1(new_n998), .A2(new_n1004), .A3(new_n713), .ZN(new_n1005));
  XNOR2_X1  g804(.A(new_n1005), .B(KEYINPUT62), .ZN(new_n1006));
  AOI21_X1  g805(.A(new_n1004), .B1(new_n1001), .B2(new_n713), .ZN(new_n1007));
  NOR2_X1   g806(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g807(.A(KEYINPUT127), .ZN(new_n1009));
  XNOR2_X1  g808(.A(new_n1008), .B(new_n1009), .ZN(G1353gat));
  AOI21_X1  g809(.A(new_n359), .B1(new_n1001), .B2(new_n803), .ZN(new_n1011));
  XNOR2_X1  g810(.A(new_n1011), .B(KEYINPUT63), .ZN(new_n1012));
  NAND3_X1  g811(.A1(new_n998), .A2(new_n359), .A3(new_n803), .ZN(new_n1013));
  NAND2_X1  g812(.A1(new_n1012), .A2(new_n1013), .ZN(G1354gat));
  NAND3_X1  g813(.A1(new_n998), .A2(new_n360), .A3(new_n683), .ZN(new_n1015));
  AND2_X1   g814(.A1(new_n1001), .A2(new_n683), .ZN(new_n1016));
  OAI21_X1  g815(.A(new_n1015), .B1(new_n1016), .B2(new_n360), .ZN(G1355gat));
endmodule


