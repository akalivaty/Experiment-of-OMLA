

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575;

  INV_X1 U318 ( .A(KEYINPUT114), .ZN(n388) );
  XNOR2_X1 U319 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n356) );
  XNOR2_X1 U320 ( .A(n357), .B(n356), .ZN(n379) );
  XNOR2_X1 U321 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U322 ( .A(n329), .B(n328), .ZN(n333) );
  NOR2_X1 U323 ( .A1(n503), .A2(n409), .ZN(n558) );
  XOR2_X1 U324 ( .A(n450), .B(KEYINPUT28), .Z(n520) );
  XNOR2_X1 U325 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n441) );
  XNOR2_X1 U326 ( .A(n442), .B(n441), .ZN(G1351GAT) );
  XOR2_X1 U327 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n287) );
  XNOR2_X1 U328 ( .A(G36GAT), .B(KEYINPUT64), .ZN(n286) );
  XNOR2_X1 U329 ( .A(n287), .B(n286), .ZN(n288) );
  XOR2_X1 U330 ( .A(G50GAT), .B(G162GAT), .Z(n411) );
  XOR2_X1 U331 ( .A(n288), .B(n411), .Z(n291) );
  XNOR2_X1 U332 ( .A(G29GAT), .B(KEYINPUT7), .ZN(n289) );
  XNOR2_X1 U333 ( .A(n289), .B(KEYINPUT8), .ZN(n348) );
  XOR2_X1 U334 ( .A(G43GAT), .B(G134GAT), .Z(n435) );
  XNOR2_X1 U335 ( .A(n348), .B(n435), .ZN(n290) );
  XNOR2_X1 U336 ( .A(n291), .B(n290), .ZN(n292) );
  XOR2_X1 U337 ( .A(n292), .B(KEYINPUT10), .Z(n294) );
  XOR2_X1 U338 ( .A(G99GAT), .B(G85GAT), .Z(n321) );
  XNOR2_X1 U339 ( .A(G218GAT), .B(n321), .ZN(n293) );
  XOR2_X1 U340 ( .A(n294), .B(n293), .Z(n299) );
  XOR2_X1 U341 ( .A(G92GAT), .B(G106GAT), .Z(n296) );
  NAND2_X1 U342 ( .A1(G232GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U343 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U344 ( .A(G190GAT), .B(n297), .Z(n298) );
  XNOR2_X1 U345 ( .A(n299), .B(n298), .ZN(n544) );
  INV_X1 U346 ( .A(n544), .ZN(n529) );
  XOR2_X1 U347 ( .A(KEYINPUT55), .B(KEYINPUT122), .Z(n426) );
  XOR2_X1 U348 ( .A(G85GAT), .B(G162GAT), .Z(n301) );
  XNOR2_X1 U349 ( .A(G29GAT), .B(G134GAT), .ZN(n300) );
  XNOR2_X1 U350 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U351 ( .A(KEYINPUT91), .B(G155GAT), .Z(n303) );
  XNOR2_X1 U352 ( .A(G127GAT), .B(G148GAT), .ZN(n302) );
  XNOR2_X1 U353 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U354 ( .A(n305), .B(n304), .Z(n310) );
  XOR2_X1 U355 ( .A(KEYINPUT90), .B(KEYINPUT4), .Z(n307) );
  NAND2_X1 U356 ( .A1(G225GAT), .A2(G233GAT), .ZN(n306) );
  XNOR2_X1 U357 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U358 ( .A(KEYINPUT5), .B(n308), .ZN(n309) );
  XNOR2_X1 U359 ( .A(n310), .B(n309), .ZN(n314) );
  XOR2_X1 U360 ( .A(G57GAT), .B(KEYINPUT1), .Z(n312) );
  XNOR2_X1 U361 ( .A(G1GAT), .B(KEYINPUT6), .ZN(n311) );
  XNOR2_X1 U362 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U363 ( .A(n314), .B(n313), .Z(n320) );
  XOR2_X1 U364 ( .A(G120GAT), .B(KEYINPUT79), .Z(n316) );
  XNOR2_X1 U365 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n315) );
  XNOR2_X1 U366 ( .A(n316), .B(n315), .ZN(n427) );
  XOR2_X1 U367 ( .A(KEYINPUT2), .B(KEYINPUT88), .Z(n318) );
  XNOR2_X1 U368 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n317) );
  XNOR2_X1 U369 ( .A(n318), .B(n317), .ZN(n414) );
  XNOR2_X1 U370 ( .A(n427), .B(n414), .ZN(n319) );
  XNOR2_X1 U371 ( .A(n320), .B(n319), .ZN(n503) );
  XOR2_X1 U372 ( .A(G92GAT), .B(G64GAT), .Z(n403) );
  XNOR2_X1 U373 ( .A(n403), .B(n321), .ZN(n323) );
  XOR2_X1 U374 ( .A(G176GAT), .B(G204GAT), .Z(n322) );
  XNOR2_X1 U375 ( .A(n323), .B(n322), .ZN(n329) );
  XOR2_X1 U376 ( .A(KEYINPUT32), .B(KEYINPUT69), .Z(n325) );
  XNOR2_X1 U377 ( .A(KEYINPUT33), .B(KEYINPUT73), .ZN(n324) );
  XOR2_X1 U378 ( .A(n325), .B(n324), .Z(n327) );
  NAND2_X1 U379 ( .A1(G230GAT), .A2(G233GAT), .ZN(n326) );
  XOR2_X1 U380 ( .A(KEYINPUT72), .B(KEYINPUT70), .Z(n331) );
  XNOR2_X1 U381 ( .A(G120GAT), .B(KEYINPUT31), .ZN(n330) );
  XOR2_X1 U382 ( .A(n331), .B(n330), .Z(n332) );
  XNOR2_X1 U383 ( .A(n333), .B(n332), .ZN(n338) );
  XOR2_X1 U384 ( .A(G78GAT), .B(G148GAT), .Z(n335) );
  XNOR2_X1 U385 ( .A(G106GAT), .B(KEYINPUT71), .ZN(n334) );
  XNOR2_X1 U386 ( .A(n335), .B(n334), .ZN(n410) );
  XNOR2_X1 U387 ( .A(G71GAT), .B(G57GAT), .ZN(n336) );
  XNOR2_X1 U388 ( .A(n336), .B(KEYINPUT13), .ZN(n364) );
  XNOR2_X1 U389 ( .A(n410), .B(n364), .ZN(n337) );
  XNOR2_X1 U390 ( .A(n338), .B(n337), .ZN(n564) );
  XNOR2_X1 U391 ( .A(n564), .B(KEYINPUT41), .ZN(n549) );
  XOR2_X1 U392 ( .A(G15GAT), .B(G113GAT), .Z(n340) );
  XNOR2_X1 U393 ( .A(G169GAT), .B(G197GAT), .ZN(n339) );
  XNOR2_X1 U394 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U395 ( .A(KEYINPUT68), .B(KEYINPUT67), .Z(n342) );
  XNOR2_X1 U396 ( .A(KEYINPUT65), .B(KEYINPUT30), .ZN(n341) );
  XNOR2_X1 U397 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U398 ( .A(n344), .B(n343), .ZN(n355) );
  XOR2_X1 U399 ( .A(G22GAT), .B(G141GAT), .Z(n346) );
  XOR2_X1 U400 ( .A(G36GAT), .B(G8GAT), .Z(n398) );
  XOR2_X1 U401 ( .A(G1GAT), .B(KEYINPUT66), .Z(n361) );
  XNOR2_X1 U402 ( .A(n398), .B(n361), .ZN(n345) );
  XNOR2_X1 U403 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U404 ( .A(n347), .B(G43GAT), .Z(n353) );
  XOR2_X1 U405 ( .A(n348), .B(KEYINPUT29), .Z(n350) );
  NAND2_X1 U406 ( .A1(G229GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U407 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U408 ( .A(n351), .B(G50GAT), .ZN(n352) );
  XNOR2_X1 U409 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U410 ( .A(n355), .B(n354), .ZN(n547) );
  NAND2_X1 U411 ( .A1(n549), .A2(n547), .ZN(n357) );
  XOR2_X1 U412 ( .A(G64GAT), .B(G78GAT), .Z(n359) );
  XNOR2_X1 U413 ( .A(G183GAT), .B(G211GAT), .ZN(n358) );
  XNOR2_X1 U414 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U415 ( .A(n360), .B(KEYINPUT12), .Z(n363) );
  XNOR2_X1 U416 ( .A(G8GAT), .B(n361), .ZN(n362) );
  XNOR2_X1 U417 ( .A(n363), .B(n362), .ZN(n365) );
  XOR2_X1 U418 ( .A(n365), .B(n364), .Z(n367) );
  XOR2_X1 U419 ( .A(G15GAT), .B(G127GAT), .Z(n434) );
  XOR2_X1 U420 ( .A(G22GAT), .B(G155GAT), .Z(n412) );
  XNOR2_X1 U421 ( .A(n434), .B(n412), .ZN(n366) );
  XNOR2_X1 U422 ( .A(n367), .B(n366), .ZN(n371) );
  XOR2_X1 U423 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n369) );
  NAND2_X1 U424 ( .A1(G231GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U425 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U426 ( .A(n371), .B(n370), .ZN(n376) );
  XOR2_X1 U427 ( .A(KEYINPUT77), .B(KEYINPUT78), .Z(n373) );
  XNOR2_X1 U428 ( .A(KEYINPUT74), .B(KEYINPUT75), .ZN(n372) );
  XNOR2_X1 U429 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U430 ( .A(n374), .B(KEYINPUT76), .ZN(n375) );
  XNOR2_X1 U431 ( .A(n376), .B(n375), .ZN(n568) );
  INV_X1 U432 ( .A(KEYINPUT111), .ZN(n377) );
  XNOR2_X1 U433 ( .A(n568), .B(n377), .ZN(n555) );
  AND2_X1 U434 ( .A1(n555), .A2(n544), .ZN(n378) );
  AND2_X1 U435 ( .A1(n379), .A2(n378), .ZN(n380) );
  XNOR2_X1 U436 ( .A(n380), .B(KEYINPUT47), .ZN(n386) );
  XNOR2_X1 U437 ( .A(KEYINPUT36), .B(n544), .ZN(n572) );
  NOR2_X1 U438 ( .A1(n572), .A2(n568), .ZN(n381) );
  XNOR2_X1 U439 ( .A(KEYINPUT45), .B(n381), .ZN(n382) );
  NAND2_X1 U440 ( .A1(n382), .A2(n564), .ZN(n383) );
  XNOR2_X1 U441 ( .A(n383), .B(KEYINPUT113), .ZN(n384) );
  INV_X1 U442 ( .A(n547), .ZN(n559) );
  NAND2_X1 U443 ( .A1(n384), .A2(n559), .ZN(n385) );
  NAND2_X1 U444 ( .A1(n386), .A2(n385), .ZN(n387) );
  XNOR2_X1 U445 ( .A(n387), .B(KEYINPUT48), .ZN(n389) );
  XNOR2_X1 U446 ( .A(n389), .B(n388), .ZN(n516) );
  XOR2_X1 U447 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n391) );
  XNOR2_X1 U448 ( .A(G176GAT), .B(KEYINPUT82), .ZN(n390) );
  XNOR2_X1 U449 ( .A(n391), .B(n390), .ZN(n395) );
  XOR2_X1 U450 ( .A(KEYINPUT83), .B(KEYINPUT84), .Z(n393) );
  XNOR2_X1 U451 ( .A(G190GAT), .B(KEYINPUT17), .ZN(n392) );
  XNOR2_X1 U452 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U453 ( .A(n395), .B(n394), .Z(n397) );
  XNOR2_X1 U454 ( .A(G169GAT), .B(G183GAT), .ZN(n396) );
  XNOR2_X1 U455 ( .A(n397), .B(n396), .ZN(n439) );
  XNOR2_X1 U456 ( .A(n398), .B(n439), .ZN(n407) );
  XNOR2_X1 U457 ( .A(G211GAT), .B(G218GAT), .ZN(n399) );
  XNOR2_X1 U458 ( .A(n399), .B(KEYINPUT21), .ZN(n400) );
  XOR2_X1 U459 ( .A(n400), .B(KEYINPUT87), .Z(n402) );
  XNOR2_X1 U460 ( .A(G197GAT), .B(G204GAT), .ZN(n401) );
  XNOR2_X1 U461 ( .A(n402), .B(n401), .ZN(n422) );
  XOR2_X1 U462 ( .A(n403), .B(n422), .Z(n405) );
  NAND2_X1 U463 ( .A1(G226GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U464 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U465 ( .A(n407), .B(n406), .ZN(n446) );
  NOR2_X1 U466 ( .A1(n516), .A2(n446), .ZN(n408) );
  XOR2_X1 U467 ( .A(KEYINPUT54), .B(n408), .Z(n409) );
  XNOR2_X1 U468 ( .A(n411), .B(n410), .ZN(n413) );
  XNOR2_X1 U469 ( .A(n413), .B(n412), .ZN(n418) );
  XOR2_X1 U470 ( .A(n414), .B(KEYINPUT89), .Z(n416) );
  NAND2_X1 U471 ( .A1(G228GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U472 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U473 ( .A(n418), .B(n417), .Z(n424) );
  XOR2_X1 U474 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n420) );
  XNOR2_X1 U475 ( .A(KEYINPUT23), .B(KEYINPUT86), .ZN(n419) );
  XNOR2_X1 U476 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U477 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U478 ( .A(n424), .B(n423), .ZN(n450) );
  NAND2_X1 U479 ( .A1(n558), .A2(n450), .ZN(n425) );
  XOR2_X1 U480 ( .A(n426), .B(n425), .Z(n440) );
  XOR2_X1 U481 ( .A(KEYINPUT20), .B(n427), .Z(n429) );
  NAND2_X1 U482 ( .A1(G227GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U483 ( .A(n429), .B(n428), .ZN(n433) );
  XOR2_X1 U484 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n431) );
  XNOR2_X1 U485 ( .A(G99GAT), .B(G71GAT), .ZN(n430) );
  XNOR2_X1 U486 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U487 ( .A(n433), .B(n432), .Z(n437) );
  XNOR2_X1 U488 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U489 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X2 U490 ( .A(n439), .B(n438), .Z(n517) );
  NAND2_X1 U491 ( .A1(n440), .A2(n517), .ZN(n554) );
  INV_X1 U492 ( .A(n554), .ZN(n550) );
  NAND2_X1 U493 ( .A1(n529), .A2(n550), .ZN(n442) );
  XOR2_X1 U494 ( .A(KEYINPUT94), .B(KEYINPUT34), .Z(n462) );
  NAND2_X1 U495 ( .A1(n547), .A2(n564), .ZN(n475) );
  NOR2_X1 U496 ( .A1(n529), .A2(n568), .ZN(n443) );
  XNOR2_X1 U497 ( .A(n443), .B(KEYINPUT16), .ZN(n460) );
  XNOR2_X1 U498 ( .A(n517), .B(KEYINPUT85), .ZN(n445) );
  XOR2_X1 U499 ( .A(n446), .B(KEYINPUT27), .Z(n452) );
  NAND2_X1 U500 ( .A1(n503), .A2(n452), .ZN(n515) );
  NOR2_X1 U501 ( .A1(n520), .A2(n515), .ZN(n444) );
  NAND2_X1 U502 ( .A1(n445), .A2(n444), .ZN(n459) );
  INV_X1 U503 ( .A(n503), .ZN(n457) );
  INV_X1 U504 ( .A(n446), .ZN(n507) );
  NAND2_X1 U505 ( .A1(n507), .A2(n517), .ZN(n447) );
  NAND2_X1 U506 ( .A1(n447), .A2(n450), .ZN(n448) );
  XNOR2_X1 U507 ( .A(n448), .B(KEYINPUT93), .ZN(n449) );
  XNOR2_X1 U508 ( .A(KEYINPUT25), .B(n449), .ZN(n455) );
  NOR2_X1 U509 ( .A1(n450), .A2(n517), .ZN(n451) );
  XNOR2_X1 U510 ( .A(n451), .B(KEYINPUT26), .ZN(n557) );
  NAND2_X1 U511 ( .A1(n452), .A2(n557), .ZN(n453) );
  XNOR2_X1 U512 ( .A(KEYINPUT92), .B(n453), .ZN(n454) );
  NAND2_X1 U513 ( .A1(n455), .A2(n454), .ZN(n456) );
  NAND2_X1 U514 ( .A1(n457), .A2(n456), .ZN(n458) );
  NAND2_X1 U515 ( .A1(n459), .A2(n458), .ZN(n471) );
  NAND2_X1 U516 ( .A1(n460), .A2(n471), .ZN(n488) );
  NOR2_X1 U517 ( .A1(n475), .A2(n488), .ZN(n469) );
  NAND2_X1 U518 ( .A1(n469), .A2(n503), .ZN(n461) );
  XNOR2_X1 U519 ( .A(n462), .B(n461), .ZN(n463) );
  XOR2_X1 U520 ( .A(G1GAT), .B(n463), .Z(G1324GAT) );
  NAND2_X1 U521 ( .A1(n507), .A2(n469), .ZN(n464) );
  XNOR2_X1 U522 ( .A(n464), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U523 ( .A(KEYINPUT96), .B(KEYINPUT35), .Z(n466) );
  NAND2_X1 U524 ( .A1(n469), .A2(n517), .ZN(n465) );
  XNOR2_X1 U525 ( .A(n466), .B(n465), .ZN(n468) );
  XOR2_X1 U526 ( .A(G15GAT), .B(KEYINPUT95), .Z(n467) );
  XNOR2_X1 U527 ( .A(n468), .B(n467), .ZN(G1326GAT) );
  NAND2_X1 U528 ( .A1(n469), .A2(n520), .ZN(n470) );
  XNOR2_X1 U529 ( .A(n470), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U530 ( .A(KEYINPUT97), .B(KEYINPUT39), .Z(n479) );
  NAND2_X1 U531 ( .A1(n568), .A2(n471), .ZN(n472) );
  NOR2_X1 U532 ( .A1(n572), .A2(n472), .ZN(n474) );
  XNOR2_X1 U533 ( .A(KEYINPUT37), .B(KEYINPUT98), .ZN(n473) );
  XNOR2_X1 U534 ( .A(n474), .B(n473), .ZN(n502) );
  NOR2_X1 U535 ( .A1(n502), .A2(n475), .ZN(n476) );
  XOR2_X1 U536 ( .A(KEYINPUT38), .B(n476), .Z(n477) );
  XNOR2_X1 U537 ( .A(KEYINPUT99), .B(n477), .ZN(n484) );
  NAND2_X1 U538 ( .A1(n503), .A2(n484), .ZN(n478) );
  XNOR2_X1 U539 ( .A(n479), .B(n478), .ZN(n480) );
  XOR2_X1 U540 ( .A(G29GAT), .B(n480), .Z(G1328GAT) );
  NAND2_X1 U541 ( .A1(n484), .A2(n507), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n481), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U543 ( .A1(n484), .A2(n517), .ZN(n482) );
  XNOR2_X1 U544 ( .A(n482), .B(KEYINPUT40), .ZN(n483) );
  XNOR2_X1 U545 ( .A(G43GAT), .B(n483), .ZN(G1330GAT) );
  XOR2_X1 U546 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n486) );
  NAND2_X1 U547 ( .A1(n520), .A2(n484), .ZN(n485) );
  XNOR2_X1 U548 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U549 ( .A(G50GAT), .B(n487), .ZN(G1331GAT) );
  XOR2_X1 U550 ( .A(KEYINPUT102), .B(KEYINPUT42), .Z(n490) );
  NAND2_X1 U551 ( .A1(n559), .A2(n549), .ZN(n501) );
  NOR2_X1 U552 ( .A1(n501), .A2(n488), .ZN(n496) );
  NAND2_X1 U553 ( .A1(n496), .A2(n503), .ZN(n489) );
  XNOR2_X1 U554 ( .A(n490), .B(n489), .ZN(n491) );
  XOR2_X1 U555 ( .A(G57GAT), .B(n491), .Z(G1332GAT) );
  XOR2_X1 U556 ( .A(G64GAT), .B(KEYINPUT103), .Z(n493) );
  NAND2_X1 U557 ( .A1(n496), .A2(n507), .ZN(n492) );
  XNOR2_X1 U558 ( .A(n493), .B(n492), .ZN(G1333GAT) );
  NAND2_X1 U559 ( .A1(n496), .A2(n517), .ZN(n494) );
  XNOR2_X1 U560 ( .A(n494), .B(KEYINPUT104), .ZN(n495) );
  XNOR2_X1 U561 ( .A(G71GAT), .B(n495), .ZN(G1334GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT106), .B(KEYINPUT43), .Z(n498) );
  NAND2_X1 U563 ( .A1(n496), .A2(n520), .ZN(n497) );
  XNOR2_X1 U564 ( .A(n498), .B(n497), .ZN(n500) );
  XOR2_X1 U565 ( .A(G78GAT), .B(KEYINPUT105), .Z(n499) );
  XNOR2_X1 U566 ( .A(n500), .B(n499), .ZN(G1335GAT) );
  XOR2_X1 U567 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n505) );
  NOR2_X1 U568 ( .A1(n502), .A2(n501), .ZN(n510) );
  NAND2_X1 U569 ( .A1(n510), .A2(n503), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U571 ( .A(G85GAT), .B(n506), .ZN(G1336GAT) );
  NAND2_X1 U572 ( .A1(n507), .A2(n510), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n508), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U574 ( .A1(n510), .A2(n517), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n509), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U576 ( .A(G106GAT), .B(KEYINPUT109), .ZN(n514) );
  XOR2_X1 U577 ( .A(KEYINPUT44), .B(KEYINPUT110), .Z(n512) );
  NAND2_X1 U578 ( .A1(n510), .A2(n520), .ZN(n511) );
  XNOR2_X1 U579 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n514), .B(n513), .ZN(G1339GAT) );
  NOR2_X1 U581 ( .A1(n516), .A2(n515), .ZN(n534) );
  NAND2_X1 U582 ( .A1(n517), .A2(n534), .ZN(n518) );
  XOR2_X1 U583 ( .A(KEYINPUT115), .B(n518), .Z(n519) );
  NOR2_X1 U584 ( .A1(n520), .A2(n519), .ZN(n530) );
  NAND2_X1 U585 ( .A1(n530), .A2(n547), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n521), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U587 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n523) );
  NAND2_X1 U588 ( .A1(n530), .A2(n549), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U590 ( .A(G120GAT), .B(n524), .ZN(G1341GAT) );
  INV_X1 U591 ( .A(n530), .ZN(n525) );
  NOR2_X1 U592 ( .A1(n555), .A2(n525), .ZN(n527) );
  XNOR2_X1 U593 ( .A(KEYINPUT50), .B(KEYINPUT117), .ZN(n526) );
  XNOR2_X1 U594 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U595 ( .A(G127GAT), .B(n528), .ZN(G1342GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n532) );
  NAND2_X1 U597 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U598 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U599 ( .A(G134GAT), .B(n533), .ZN(G1343GAT) );
  NAND2_X1 U600 ( .A1(n534), .A2(n557), .ZN(n543) );
  NOR2_X1 U601 ( .A1(n559), .A2(n543), .ZN(n535) );
  XOR2_X1 U602 ( .A(G141GAT), .B(n535), .Z(G1344GAT) );
  INV_X1 U603 ( .A(n549), .ZN(n536) );
  NOR2_X1 U604 ( .A1(n543), .A2(n536), .ZN(n540) );
  XOR2_X1 U605 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n538) );
  XNOR2_X1 U606 ( .A(G148GAT), .B(KEYINPUT119), .ZN(n537) );
  XNOR2_X1 U607 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U608 ( .A(n540), .B(n539), .ZN(G1345GAT) );
  NOR2_X1 U609 ( .A1(n568), .A2(n543), .ZN(n541) );
  XOR2_X1 U610 ( .A(KEYINPUT120), .B(n541), .Z(n542) );
  XNOR2_X1 U611 ( .A(G155GAT), .B(n542), .ZN(G1346GAT) );
  NOR2_X1 U612 ( .A1(n544), .A2(n543), .ZN(n546) );
  XNOR2_X1 U613 ( .A(G162GAT), .B(KEYINPUT121), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n546), .B(n545), .ZN(G1347GAT) );
  NAND2_X1 U615 ( .A1(n550), .A2(n547), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n548), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U617 ( .A1(n550), .A2(n549), .ZN(n552) );
  XOR2_X1 U618 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U620 ( .A(G176GAT), .B(n553), .ZN(G1349GAT) );
  NOR2_X1 U621 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U622 ( .A(G183GAT), .B(n556), .Z(G1350GAT) );
  NAND2_X1 U623 ( .A1(n558), .A2(n557), .ZN(n571) );
  NOR2_X1 U624 ( .A1(n571), .A2(n559), .ZN(n563) );
  XOR2_X1 U625 ( .A(KEYINPUT59), .B(KEYINPUT123), .Z(n561) );
  XNOR2_X1 U626 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n563), .B(n562), .ZN(G1352GAT) );
  NOR2_X1 U629 ( .A1(n564), .A2(n571), .ZN(n566) );
  XNOR2_X1 U630 ( .A(KEYINPUT124), .B(KEYINPUT61), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U632 ( .A(G204GAT), .B(n567), .ZN(G1353GAT) );
  NOR2_X1 U633 ( .A1(n568), .A2(n571), .ZN(n570) );
  XNOR2_X1 U634 ( .A(G211GAT), .B(KEYINPUT125), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G1354GAT) );
  NOR2_X1 U636 ( .A1(n572), .A2(n571), .ZN(n574) );
  XNOR2_X1 U637 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n574), .B(n573), .ZN(n575) );
  XOR2_X1 U639 ( .A(G218GAT), .B(n575), .Z(G1355GAT) );
endmodule

