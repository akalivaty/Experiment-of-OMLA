

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580;

  AND2_X1 U321 ( .A1(G230GAT), .A2(G233GAT), .ZN(n289) );
  AND2_X1 U322 ( .A1(G232GAT), .A2(G233GAT), .ZN(n290) );
  XOR2_X1 U323 ( .A(G85GAT), .B(G92GAT), .Z(n395) );
  XNOR2_X1 U324 ( .A(n381), .B(n380), .ZN(n385) );
  AND2_X1 U325 ( .A1(n419), .A2(n418), .ZN(n420) );
  XNOR2_X1 U326 ( .A(n403), .B(n290), .ZN(n404) );
  XOR2_X1 U327 ( .A(n556), .B(KEYINPUT36), .Z(n577) );
  XNOR2_X1 U328 ( .A(n405), .B(n404), .ZN(n411) );
  NOR2_X1 U329 ( .A1(n497), .A2(n450), .ZN(n557) );
  XOR2_X1 U330 ( .A(KEYINPUT41), .B(n568), .Z(n546) );
  XNOR2_X1 U331 ( .A(G183GAT), .B(KEYINPUT122), .ZN(n451) );
  XNOR2_X1 U332 ( .A(n452), .B(n451), .ZN(G1350GAT) );
  XOR2_X1 U333 ( .A(KEYINPUT14), .B(KEYINPUT81), .Z(n292) );
  XNOR2_X1 U334 ( .A(KEYINPUT15), .B(KEYINPUT80), .ZN(n291) );
  XNOR2_X1 U335 ( .A(n292), .B(n291), .ZN(n297) );
  XNOR2_X1 U336 ( .A(G57GAT), .B(KEYINPUT71), .ZN(n293) );
  XNOR2_X1 U337 ( .A(n293), .B(KEYINPUT13), .ZN(n380) );
  XOR2_X1 U338 ( .A(n380), .B(G155GAT), .Z(n295) );
  XOR2_X1 U339 ( .A(G8GAT), .B(G1GAT), .Z(n374) );
  XNOR2_X1 U340 ( .A(n374), .B(G211GAT), .ZN(n294) );
  XNOR2_X1 U341 ( .A(n295), .B(n294), .ZN(n296) );
  XNOR2_X1 U342 ( .A(n297), .B(n296), .ZN(n310) );
  XOR2_X1 U343 ( .A(G78GAT), .B(G71GAT), .Z(n299) );
  XNOR2_X1 U344 ( .A(G15GAT), .B(G22GAT), .ZN(n298) );
  XNOR2_X1 U345 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U346 ( .A(KEYINPUT83), .B(G64GAT), .Z(n301) );
  XNOR2_X1 U347 ( .A(G183GAT), .B(G127GAT), .ZN(n300) );
  XNOR2_X1 U348 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U349 ( .A(n303), .B(n302), .Z(n308) );
  XOR2_X1 U350 ( .A(KEYINPUT84), .B(KEYINPUT82), .Z(n305) );
  NAND2_X1 U351 ( .A1(G231GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U352 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U353 ( .A(KEYINPUT12), .B(n306), .ZN(n307) );
  XNOR2_X1 U354 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U355 ( .A(n310), .B(n309), .Z(n572) );
  XOR2_X1 U356 ( .A(KEYINPUT20), .B(KEYINPUT87), .Z(n312) );
  XOR2_X1 U357 ( .A(G190GAT), .B(G134GAT), .Z(n396) );
  XOR2_X1 U358 ( .A(KEYINPUT0), .B(G127GAT), .Z(n428) );
  XNOR2_X1 U359 ( .A(n396), .B(n428), .ZN(n311) );
  XNOR2_X1 U360 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U361 ( .A(n313), .B(G176GAT), .Z(n319) );
  XNOR2_X1 U362 ( .A(G99GAT), .B(G71GAT), .ZN(n314) );
  XNOR2_X1 U363 ( .A(n314), .B(G120GAT), .ZN(n387) );
  XOR2_X1 U364 ( .A(n387), .B(KEYINPUT65), .Z(n316) );
  NAND2_X1 U365 ( .A1(G227GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U366 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U367 ( .A(G43GAT), .B(n317), .ZN(n318) );
  XNOR2_X1 U368 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U369 ( .A(KEYINPUT88), .B(KEYINPUT86), .Z(n321) );
  XNOR2_X1 U370 ( .A(KEYINPUT85), .B(KEYINPUT89), .ZN(n320) );
  XNOR2_X1 U371 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U372 ( .A(n323), .B(n322), .ZN(n328) );
  XNOR2_X1 U373 ( .A(G169GAT), .B(G15GAT), .ZN(n324) );
  XNOR2_X1 U374 ( .A(n324), .B(G113GAT), .ZN(n370) );
  XOR2_X1 U375 ( .A(G183GAT), .B(KEYINPUT17), .Z(n326) );
  XNOR2_X1 U376 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n325) );
  XNOR2_X1 U377 ( .A(n326), .B(n325), .ZN(n351) );
  XNOR2_X1 U378 ( .A(n370), .B(n351), .ZN(n327) );
  XNOR2_X1 U379 ( .A(n328), .B(n327), .ZN(n528) );
  INV_X1 U380 ( .A(n528), .ZN(n497) );
  XOR2_X1 U381 ( .A(KEYINPUT93), .B(G218GAT), .Z(n330) );
  XNOR2_X1 U382 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n329) );
  XNOR2_X1 U383 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U384 ( .A(G197GAT), .B(n331), .Z(n350) );
  XOR2_X1 U385 ( .A(G148GAT), .B(G106GAT), .Z(n333) );
  XNOR2_X1 U386 ( .A(KEYINPUT72), .B(G78GAT), .ZN(n332) );
  XNOR2_X1 U387 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U388 ( .A(KEYINPUT73), .B(n334), .ZN(n390) );
  XOR2_X1 U389 ( .A(n350), .B(n390), .Z(n349) );
  XOR2_X1 U390 ( .A(G204GAT), .B(KEYINPUT22), .Z(n336) );
  XNOR2_X1 U391 ( .A(KEYINPUT94), .B(KEYINPUT91), .ZN(n335) );
  XNOR2_X1 U392 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U393 ( .A(KEYINPUT23), .B(n337), .Z(n339) );
  NAND2_X1 U394 ( .A1(G228GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U395 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U396 ( .A(n340), .B(KEYINPUT92), .Z(n347) );
  XOR2_X1 U397 ( .A(G155GAT), .B(KEYINPUT3), .Z(n342) );
  XNOR2_X1 U398 ( .A(G162GAT), .B(KEYINPUT2), .ZN(n341) );
  XNOR2_X1 U399 ( .A(n342), .B(n341), .ZN(n432) );
  XOR2_X1 U400 ( .A(KEYINPUT24), .B(n432), .Z(n344) );
  XOR2_X1 U401 ( .A(G141GAT), .B(G22GAT), .Z(n375) );
  XNOR2_X1 U402 ( .A(G50GAT), .B(n375), .ZN(n343) );
  XNOR2_X1 U403 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U404 ( .A(n345), .B(KEYINPUT95), .ZN(n346) );
  XNOR2_X1 U405 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U406 ( .A(n349), .B(n348), .ZN(n465) );
  XOR2_X1 U407 ( .A(KEYINPUT102), .B(KEYINPUT101), .Z(n353) );
  XNOR2_X1 U408 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U409 ( .A(n353), .B(n352), .ZN(n359) );
  XOR2_X1 U410 ( .A(G64GAT), .B(KEYINPUT75), .Z(n355) );
  XNOR2_X1 U411 ( .A(G176GAT), .B(G204GAT), .ZN(n354) );
  XNOR2_X1 U412 ( .A(n355), .B(n354), .ZN(n386) );
  XOR2_X1 U413 ( .A(KEYINPUT78), .B(n386), .Z(n357) );
  NAND2_X1 U414 ( .A1(G226GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U415 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U416 ( .A(n359), .B(n358), .Z(n364) );
  XOR2_X1 U417 ( .A(G92GAT), .B(G8GAT), .Z(n361) );
  XNOR2_X1 U418 ( .A(G169GAT), .B(G36GAT), .ZN(n360) );
  XNOR2_X1 U419 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U420 ( .A(G190GAT), .B(n362), .ZN(n363) );
  XOR2_X1 U421 ( .A(n364), .B(n363), .Z(n519) );
  INV_X1 U422 ( .A(n519), .ZN(n493) );
  XOR2_X1 U423 ( .A(G43GAT), .B(G29GAT), .Z(n366) );
  XNOR2_X1 U424 ( .A(KEYINPUT7), .B(G50GAT), .ZN(n365) );
  XNOR2_X1 U425 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U426 ( .A(n367), .B(KEYINPUT8), .Z(n369) );
  XNOR2_X1 U427 ( .A(G36GAT), .B(KEYINPUT69), .ZN(n368) );
  XNOR2_X1 U428 ( .A(n369), .B(n368), .ZN(n409) );
  XNOR2_X1 U429 ( .A(n409), .B(n370), .ZN(n379) );
  XOR2_X1 U430 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n372) );
  NAND2_X1 U431 ( .A1(G229GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U432 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U433 ( .A(n373), .B(G197GAT), .Z(n377) );
  XNOR2_X1 U434 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U435 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U436 ( .A(n379), .B(n378), .Z(n504) );
  XOR2_X1 U437 ( .A(n504), .B(KEYINPUT70), .Z(n554) );
  XNOR2_X1 U438 ( .A(n395), .B(n289), .ZN(n381) );
  XOR2_X1 U439 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n383) );
  XNOR2_X1 U440 ( .A(KEYINPUT74), .B(KEYINPUT32), .ZN(n382) );
  XNOR2_X1 U441 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U442 ( .A(n385), .B(n384), .Z(n389) );
  XNOR2_X1 U443 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U444 ( .A(n389), .B(n388), .ZN(n392) );
  INV_X1 U445 ( .A(n390), .ZN(n391) );
  XOR2_X1 U446 ( .A(n392), .B(n391), .Z(n474) );
  XOR2_X1 U447 ( .A(KEYINPUT66), .B(KEYINPUT45), .Z(n413) );
  INV_X1 U448 ( .A(n572), .ZN(n484) );
  XOR2_X1 U449 ( .A(KEYINPUT64), .B(KEYINPUT77), .Z(n394) );
  XNOR2_X1 U450 ( .A(G99GAT), .B(G106GAT), .ZN(n393) );
  XNOR2_X1 U451 ( .A(n394), .B(n393), .ZN(n400) );
  XOR2_X1 U452 ( .A(n395), .B(G162GAT), .Z(n398) );
  XNOR2_X1 U453 ( .A(n396), .B(G218GAT), .ZN(n397) );
  XNOR2_X1 U454 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U455 ( .A(n400), .B(n399), .Z(n405) );
  XOR2_X1 U456 ( .A(KEYINPUT79), .B(KEYINPUT10), .Z(n402) );
  XNOR2_X1 U457 ( .A(KEYINPUT78), .B(KEYINPUT11), .ZN(n401) );
  XNOR2_X1 U458 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U459 ( .A(KEYINPUT76), .B(KEYINPUT67), .Z(n407) );
  XNOR2_X1 U460 ( .A(KEYINPUT9), .B(KEYINPUT68), .ZN(n406) );
  XNOR2_X1 U461 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U462 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U463 ( .A(n411), .B(n410), .ZN(n556) );
  NOR2_X1 U464 ( .A1(n484), .A2(n577), .ZN(n412) );
  XOR2_X1 U465 ( .A(n413), .B(n412), .Z(n414) );
  NAND2_X1 U466 ( .A1(n474), .A2(n414), .ZN(n415) );
  NOR2_X1 U467 ( .A1(n554), .A2(n415), .ZN(n416) );
  XNOR2_X1 U468 ( .A(n416), .B(KEYINPUT116), .ZN(n422) );
  INV_X1 U469 ( .A(n504), .ZN(n565) );
  INV_X1 U470 ( .A(n474), .ZN(n568) );
  NAND2_X1 U471 ( .A1(n565), .A2(n546), .ZN(n417) );
  XNOR2_X1 U472 ( .A(KEYINPUT46), .B(n417), .ZN(n419) );
  NOR2_X1 U473 ( .A1(n556), .A2(n572), .ZN(n418) );
  XOR2_X1 U474 ( .A(KEYINPUT47), .B(n420), .Z(n421) );
  NOR2_X1 U475 ( .A1(n422), .A2(n421), .ZN(n423) );
  XNOR2_X1 U476 ( .A(n423), .B(KEYINPUT48), .ZN(n542) );
  NOR2_X1 U477 ( .A1(n493), .A2(n542), .ZN(n424) );
  XNOR2_X1 U478 ( .A(n424), .B(KEYINPUT54), .ZN(n447) );
  XOR2_X1 U479 ( .A(G85GAT), .B(G148GAT), .Z(n426) );
  XNOR2_X1 U480 ( .A(G29GAT), .B(G134GAT), .ZN(n425) );
  XNOR2_X1 U481 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U482 ( .A(n428), .B(n427), .Z(n430) );
  NAND2_X1 U483 ( .A1(G225GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U484 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U485 ( .A(n431), .B(KEYINPUT99), .Z(n434) );
  XNOR2_X1 U486 ( .A(n432), .B(KEYINPUT97), .ZN(n433) );
  XNOR2_X1 U487 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U488 ( .A(G57GAT), .B(G120GAT), .Z(n436) );
  XNOR2_X1 U489 ( .A(G113GAT), .B(G141GAT), .ZN(n435) );
  XNOR2_X1 U490 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U491 ( .A(n438), .B(n437), .Z(n446) );
  XOR2_X1 U492 ( .A(KEYINPUT98), .B(KEYINPUT100), .Z(n440) );
  XNOR2_X1 U493 ( .A(KEYINPUT96), .B(KEYINPUT6), .ZN(n439) );
  XNOR2_X1 U494 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U495 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n442) );
  XNOR2_X1 U496 ( .A(G1GAT), .B(KEYINPUT1), .ZN(n441) );
  XNOR2_X1 U497 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U498 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U499 ( .A(n446), .B(n445), .Z(n540) );
  INV_X1 U500 ( .A(n540), .ZN(n489) );
  NAND2_X1 U501 ( .A1(n447), .A2(n489), .ZN(n564) );
  NOR2_X1 U502 ( .A1(n465), .A2(n564), .ZN(n449) );
  XNOR2_X1 U503 ( .A(KEYINPUT55), .B(KEYINPUT120), .ZN(n448) );
  XNOR2_X1 U504 ( .A(n449), .B(n448), .ZN(n450) );
  NAND2_X1 U505 ( .A1(n572), .A2(n557), .ZN(n452) );
  NAND2_X1 U506 ( .A1(n557), .A2(n546), .ZN(n456) );
  XOR2_X1 U507 ( .A(KEYINPUT121), .B(KEYINPUT57), .Z(n454) );
  XOR2_X1 U508 ( .A(G176GAT), .B(KEYINPUT56), .Z(n453) );
  XNOR2_X1 U509 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U510 ( .A(n456), .B(n455), .ZN(G1349GAT) );
  XNOR2_X1 U511 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n476) );
  XNOR2_X1 U512 ( .A(n528), .B(KEYINPUT90), .ZN(n459) );
  XOR2_X1 U513 ( .A(n519), .B(KEYINPUT27), .Z(n462) );
  XNOR2_X1 U514 ( .A(n465), .B(KEYINPUT28), .ZN(n523) );
  OR2_X1 U515 ( .A1(n462), .A2(n523), .ZN(n457) );
  NOR2_X1 U516 ( .A1(n489), .A2(n457), .ZN(n529) );
  XNOR2_X1 U517 ( .A(n529), .B(KEYINPUT103), .ZN(n458) );
  NOR2_X1 U518 ( .A1(n459), .A2(n458), .ZN(n470) );
  NAND2_X1 U519 ( .A1(n465), .A2(n497), .ZN(n460) );
  XNOR2_X1 U520 ( .A(n460), .B(KEYINPUT26), .ZN(n461) );
  XNOR2_X1 U521 ( .A(KEYINPUT104), .B(n461), .ZN(n563) );
  NOR2_X1 U522 ( .A1(n563), .A2(n462), .ZN(n541) );
  NOR2_X1 U523 ( .A1(n497), .A2(n493), .ZN(n463) );
  XOR2_X1 U524 ( .A(KEYINPUT105), .B(n463), .Z(n464) );
  NOR2_X1 U525 ( .A1(n465), .A2(n464), .ZN(n466) );
  XOR2_X1 U526 ( .A(KEYINPUT25), .B(n466), .Z(n467) );
  NOR2_X1 U527 ( .A1(n541), .A2(n467), .ZN(n468) );
  NOR2_X1 U528 ( .A1(n468), .A2(n540), .ZN(n469) );
  NOR2_X1 U529 ( .A1(n470), .A2(n469), .ZN(n483) );
  NOR2_X1 U530 ( .A1(n556), .A2(n484), .ZN(n471) );
  XOR2_X1 U531 ( .A(KEYINPUT16), .B(n471), .Z(n472) );
  NOR2_X1 U532 ( .A1(n483), .A2(n472), .ZN(n473) );
  XOR2_X1 U533 ( .A(KEYINPUT106), .B(n473), .Z(n505) );
  NAND2_X1 U534 ( .A1(n474), .A2(n554), .ZN(n487) );
  NOR2_X1 U535 ( .A1(n505), .A2(n487), .ZN(n480) );
  NAND2_X1 U536 ( .A1(n480), .A2(n540), .ZN(n475) );
  XNOR2_X1 U537 ( .A(n476), .B(n475), .ZN(G1324GAT) );
  NAND2_X1 U538 ( .A1(n480), .A2(n519), .ZN(n477) );
  XNOR2_X1 U539 ( .A(G8GAT), .B(n477), .ZN(G1325GAT) );
  XOR2_X1 U540 ( .A(G15GAT), .B(KEYINPUT35), .Z(n479) );
  NAND2_X1 U541 ( .A1(n480), .A2(n528), .ZN(n478) );
  XNOR2_X1 U542 ( .A(n479), .B(n478), .ZN(G1326GAT) );
  XOR2_X1 U543 ( .A(G22GAT), .B(KEYINPUT107), .Z(n482) );
  NAND2_X1 U544 ( .A1(n480), .A2(n523), .ZN(n481) );
  XNOR2_X1 U545 ( .A(n482), .B(n481), .ZN(G1327GAT) );
  XNOR2_X1 U546 ( .A(KEYINPUT108), .B(KEYINPUT39), .ZN(n491) );
  NOR2_X1 U547 ( .A1(n577), .A2(n483), .ZN(n485) );
  NAND2_X1 U548 ( .A1(n485), .A2(n484), .ZN(n486) );
  XOR2_X1 U549 ( .A(KEYINPUT37), .B(n486), .Z(n517) );
  NOR2_X1 U550 ( .A1(n517), .A2(n487), .ZN(n488) );
  XOR2_X1 U551 ( .A(KEYINPUT38), .B(n488), .Z(n501) );
  NOR2_X1 U552 ( .A1(n489), .A2(n501), .ZN(n490) );
  XNOR2_X1 U553 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U554 ( .A(G29GAT), .B(n492), .ZN(G1328GAT) );
  XNOR2_X1 U555 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n495) );
  NOR2_X1 U556 ( .A1(n493), .A2(n501), .ZN(n494) );
  XNOR2_X1 U557 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U558 ( .A(G36GAT), .B(n496), .ZN(G1329GAT) );
  INV_X1 U559 ( .A(KEYINPUT40), .ZN(n499) );
  NOR2_X1 U560 ( .A1(n497), .A2(n501), .ZN(n498) );
  XNOR2_X1 U561 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U562 ( .A(G43GAT), .B(n500), .ZN(G1330GAT) );
  INV_X1 U563 ( .A(n523), .ZN(n502) );
  NOR2_X1 U564 ( .A1(n502), .A2(n501), .ZN(n503) );
  XOR2_X1 U565 ( .A(G50GAT), .B(n503), .Z(G1331GAT) );
  XNOR2_X1 U566 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n507) );
  NAND2_X1 U567 ( .A1(n504), .A2(n546), .ZN(n516) );
  NOR2_X1 U568 ( .A1(n505), .A2(n516), .ZN(n512) );
  NAND2_X1 U569 ( .A1(n512), .A2(n540), .ZN(n506) );
  XNOR2_X1 U570 ( .A(n507), .B(n506), .ZN(G1332GAT) );
  XOR2_X1 U571 ( .A(G64GAT), .B(KEYINPUT111), .Z(n509) );
  NAND2_X1 U572 ( .A1(n512), .A2(n519), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n509), .B(n508), .ZN(G1333GAT) );
  NAND2_X1 U574 ( .A1(n528), .A2(n512), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n510), .B(KEYINPUT112), .ZN(n511) );
  XNOR2_X1 U576 ( .A(G71GAT), .B(n511), .ZN(G1334GAT) );
  XOR2_X1 U577 ( .A(KEYINPUT113), .B(KEYINPUT43), .Z(n514) );
  NAND2_X1 U578 ( .A1(n512), .A2(n523), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n514), .B(n513), .ZN(n515) );
  XOR2_X1 U580 ( .A(G78GAT), .B(n515), .Z(G1335GAT) );
  NOR2_X1 U581 ( .A1(n517), .A2(n516), .ZN(n524) );
  NAND2_X1 U582 ( .A1(n524), .A2(n540), .ZN(n518) );
  XNOR2_X1 U583 ( .A(G85GAT), .B(n518), .ZN(G1336GAT) );
  NAND2_X1 U584 ( .A1(n519), .A2(n524), .ZN(n520) );
  XNOR2_X1 U585 ( .A(n520), .B(KEYINPUT114), .ZN(n521) );
  XNOR2_X1 U586 ( .A(G92GAT), .B(n521), .ZN(G1337GAT) );
  NAND2_X1 U587 ( .A1(n528), .A2(n524), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n522), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT115), .B(KEYINPUT44), .Z(n526) );
  NAND2_X1 U590 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U592 ( .A(G106GAT), .B(n527), .ZN(G1339GAT) );
  XOR2_X1 U593 ( .A(G113GAT), .B(KEYINPUT117), .Z(n532) );
  NAND2_X1 U594 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U595 ( .A1(n542), .A2(n530), .ZN(n537) );
  NAND2_X1 U596 ( .A1(n537), .A2(n554), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n532), .B(n531), .ZN(G1340GAT) );
  XOR2_X1 U598 ( .A(G120GAT), .B(KEYINPUT49), .Z(n534) );
  NAND2_X1 U599 ( .A1(n537), .A2(n546), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n534), .B(n533), .ZN(G1341GAT) );
  NAND2_X1 U601 ( .A1(n572), .A2(n537), .ZN(n535) );
  XNOR2_X1 U602 ( .A(n535), .B(KEYINPUT50), .ZN(n536) );
  XNOR2_X1 U603 ( .A(G127GAT), .B(n536), .ZN(G1342GAT) );
  XOR2_X1 U604 ( .A(G134GAT), .B(KEYINPUT51), .Z(n539) );
  NAND2_X1 U605 ( .A1(n537), .A2(n556), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n539), .B(n538), .ZN(G1343GAT) );
  NAND2_X1 U607 ( .A1(n541), .A2(n540), .ZN(n543) );
  NOR2_X1 U608 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U609 ( .A(n544), .B(KEYINPUT118), .ZN(n552) );
  NAND2_X1 U610 ( .A1(n552), .A2(n565), .ZN(n545) );
  XNOR2_X1 U611 ( .A(n545), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n548) );
  NAND2_X1 U613 ( .A1(n552), .A2(n546), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(n549), .ZN(G1345GAT) );
  XOR2_X1 U616 ( .A(G155GAT), .B(KEYINPUT119), .Z(n551) );
  NAND2_X1 U617 ( .A1(n552), .A2(n572), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n551), .B(n550), .ZN(G1346GAT) );
  NAND2_X1 U619 ( .A1(n552), .A2(n556), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n553), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U621 ( .A1(n554), .A2(n557), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n555), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(KEYINPUT58), .ZN(n559) );
  XNOR2_X1 U625 ( .A(G190GAT), .B(n559), .ZN(G1351GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n561) );
  XNOR2_X1 U627 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(n562) );
  XOR2_X1 U629 ( .A(KEYINPUT60), .B(n562), .Z(n567) );
  NOR2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n575) );
  NAND2_X1 U631 ( .A1(n575), .A2(n565), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(G1352GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n570) );
  NAND2_X1 U634 ( .A1(n575), .A2(n568), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(n571) );
  XOR2_X1 U636 ( .A(G204GAT), .B(n571), .Z(G1353GAT) );
  NAND2_X1 U637 ( .A1(n572), .A2(n575), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n573), .B(KEYINPUT126), .ZN(n574) );
  XNOR2_X1 U639 ( .A(G211GAT), .B(n574), .ZN(G1354GAT) );
  INV_X1 U640 ( .A(n575), .ZN(n576) );
  NOR2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n579) );
  XNOR2_X1 U642 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U644 ( .A(G218GAT), .B(n580), .ZN(G1355GAT) );
endmodule

