

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U550 ( .A(n771), .B(KEYINPUT103), .ZN(n775) );
  OR2_X1 U551 ( .A1(n774), .A2(n773), .ZN(n516) );
  AND2_X1 U552 ( .A1(n518), .A2(n815), .ZN(n517) );
  AND2_X1 U553 ( .A1(n808), .A2(n796), .ZN(n518) );
  NOR2_X1 U554 ( .A1(n696), .A2(n695), .ZN(n700) );
  XOR2_X1 U555 ( .A(n719), .B(KEYINPUT93), .Z(n717) );
  AND2_X1 U556 ( .A1(n778), .A2(n776), .ZN(n719) );
  INV_X1 U557 ( .A(G2105), .ZN(n524) );
  NOR2_X1 U558 ( .A1(G164), .A2(G1384), .ZN(n778) );
  XOR2_X1 U559 ( .A(G543), .B(KEYINPUT0), .Z(n641) );
  NOR2_X1 U560 ( .A1(G651), .A2(n641), .ZN(n653) );
  NOR2_X1 U561 ( .A1(n539), .A2(n538), .ZN(G160) );
  NOR2_X1 U562 ( .A1(G2104), .A2(G2105), .ZN(n519) );
  XOR2_X1 U563 ( .A(KEYINPUT17), .B(n519), .Z(n529) );
  NAND2_X1 U564 ( .A1(G138), .A2(n529), .ZN(n523) );
  NAND2_X1 U565 ( .A1(n524), .A2(G2104), .ZN(n520) );
  XNOR2_X1 U566 ( .A(n520), .B(KEYINPUT65), .ZN(n534) );
  INV_X1 U567 ( .A(n534), .ZN(n521) );
  INV_X1 U568 ( .A(n521), .ZN(n872) );
  NAND2_X1 U569 ( .A1(G102), .A2(n872), .ZN(n522) );
  NAND2_X1 U570 ( .A1(n523), .A2(n522), .ZN(n528) );
  NOR2_X1 U571 ( .A1(G2104), .A2(n524), .ZN(n532) );
  BUF_X1 U572 ( .A(n532), .Z(n876) );
  NAND2_X1 U573 ( .A1(G126), .A2(n876), .ZN(n526) );
  AND2_X1 U574 ( .A1(G2104), .A2(G2105), .ZN(n877) );
  NAND2_X1 U575 ( .A1(G114), .A2(n877), .ZN(n525) );
  NAND2_X1 U576 ( .A1(n526), .A2(n525), .ZN(n527) );
  NOR2_X1 U577 ( .A1(n528), .A2(n527), .ZN(G164) );
  BUF_X1 U578 ( .A(n529), .Z(n870) );
  NAND2_X1 U579 ( .A1(G137), .A2(n870), .ZN(n531) );
  NAND2_X1 U580 ( .A1(G113), .A2(n877), .ZN(n530) );
  NAND2_X1 U581 ( .A1(n531), .A2(n530), .ZN(n539) );
  NAND2_X1 U582 ( .A1(G125), .A2(n532), .ZN(n533) );
  XNOR2_X1 U583 ( .A(n533), .B(KEYINPUT64), .ZN(n537) );
  NAND2_X1 U584 ( .A1(G101), .A2(n534), .ZN(n535) );
  XOR2_X1 U585 ( .A(KEYINPUT23), .B(n535), .Z(n536) );
  NAND2_X1 U586 ( .A1(n537), .A2(n536), .ZN(n538) );
  INV_X1 U587 ( .A(G651), .ZN(n543) );
  NOR2_X1 U588 ( .A1(G543), .A2(n543), .ZN(n540) );
  XOR2_X1 U589 ( .A(KEYINPUT1), .B(n540), .Z(n649) );
  NAND2_X1 U590 ( .A1(G64), .A2(n649), .ZN(n542) );
  NAND2_X1 U591 ( .A1(G52), .A2(n653), .ZN(n541) );
  NAND2_X1 U592 ( .A1(n542), .A2(n541), .ZN(n549) );
  NOR2_X1 U593 ( .A1(G651), .A2(G543), .ZN(n650) );
  NAND2_X1 U594 ( .A1(G90), .A2(n650), .ZN(n546) );
  OR2_X1 U595 ( .A1(n543), .A2(n641), .ZN(n544) );
  XOR2_X1 U596 ( .A(KEYINPUT66), .B(n544), .Z(n567) );
  NAND2_X1 U597 ( .A1(G77), .A2(n567), .ZN(n545) );
  NAND2_X1 U598 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U599 ( .A(KEYINPUT9), .B(n547), .Z(n548) );
  NOR2_X1 U600 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U601 ( .A(KEYINPUT69), .B(n550), .Z(G171) );
  INV_X1 U602 ( .A(G171), .ZN(G301) );
  AND2_X1 U603 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U604 ( .A(G120), .ZN(G236) );
  INV_X1 U605 ( .A(G132), .ZN(G219) );
  INV_X1 U606 ( .A(G82), .ZN(G220) );
  NAND2_X1 U607 ( .A1(n650), .A2(G89), .ZN(n551) );
  XNOR2_X1 U608 ( .A(n551), .B(KEYINPUT4), .ZN(n553) );
  BUF_X1 U609 ( .A(n567), .Z(n647) );
  NAND2_X1 U610 ( .A1(G76), .A2(n647), .ZN(n552) );
  NAND2_X1 U611 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U612 ( .A(n554), .B(KEYINPUT5), .ZN(n559) );
  NAND2_X1 U613 ( .A1(G63), .A2(n649), .ZN(n556) );
  NAND2_X1 U614 ( .A1(G51), .A2(n653), .ZN(n555) );
  NAND2_X1 U615 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U616 ( .A(KEYINPUT6), .B(n557), .Z(n558) );
  NAND2_X1 U617 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U618 ( .A(n560), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U619 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U620 ( .A(KEYINPUT71), .B(KEYINPUT10), .Z(n562) );
  NAND2_X1 U621 ( .A1(G7), .A2(G661), .ZN(n561) );
  XNOR2_X1 U622 ( .A(n562), .B(n561), .ZN(G223) );
  INV_X1 U623 ( .A(G223), .ZN(n824) );
  NAND2_X1 U624 ( .A1(n824), .A2(G567), .ZN(n563) );
  XOR2_X1 U625 ( .A(KEYINPUT11), .B(n563), .Z(G234) );
  NAND2_X1 U626 ( .A1(n649), .A2(G56), .ZN(n564) );
  XOR2_X1 U627 ( .A(KEYINPUT14), .B(n564), .Z(n573) );
  XOR2_X1 U628 ( .A(KEYINPUT72), .B(KEYINPUT12), .Z(n566) );
  NAND2_X1 U629 ( .A1(G81), .A2(n650), .ZN(n565) );
  XNOR2_X1 U630 ( .A(n566), .B(n565), .ZN(n570) );
  NAND2_X1 U631 ( .A1(G68), .A2(n567), .ZN(n568) );
  XNOR2_X1 U632 ( .A(KEYINPUT73), .B(n568), .ZN(n569) );
  NOR2_X1 U633 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U634 ( .A(n571), .B(KEYINPUT13), .ZN(n572) );
  NOR2_X1 U635 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U636 ( .A(n574), .B(KEYINPUT74), .ZN(n576) );
  NAND2_X1 U637 ( .A1(G43), .A2(n653), .ZN(n575) );
  NAND2_X1 U638 ( .A1(n576), .A2(n575), .ZN(n696) );
  INV_X1 U639 ( .A(G860), .ZN(n598) );
  OR2_X1 U640 ( .A1(n696), .A2(n598), .ZN(n577) );
  XOR2_X1 U641 ( .A(KEYINPUT75), .B(n577), .Z(G153) );
  NAND2_X1 U642 ( .A1(G868), .A2(G301), .ZN(n588) );
  NAND2_X1 U643 ( .A1(G66), .A2(n649), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n578), .B(KEYINPUT76), .ZN(n585) );
  NAND2_X1 U645 ( .A1(G54), .A2(n653), .ZN(n580) );
  NAND2_X1 U646 ( .A1(G92), .A2(n650), .ZN(n579) );
  NAND2_X1 U647 ( .A1(n580), .A2(n579), .ZN(n583) );
  NAND2_X1 U648 ( .A1(G79), .A2(n647), .ZN(n581) );
  XNOR2_X1 U649 ( .A(KEYINPUT77), .B(n581), .ZN(n582) );
  NOR2_X1 U650 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U651 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U652 ( .A(KEYINPUT15), .B(n586), .ZN(n944) );
  BUF_X1 U653 ( .A(n944), .Z(n897) );
  OR2_X1 U654 ( .A1(n897), .A2(G868), .ZN(n587) );
  NAND2_X1 U655 ( .A1(n588), .A2(n587), .ZN(G284) );
  NAND2_X1 U656 ( .A1(G65), .A2(n649), .ZN(n590) );
  NAND2_X1 U657 ( .A1(G53), .A2(n653), .ZN(n589) );
  NAND2_X1 U658 ( .A1(n590), .A2(n589), .ZN(n594) );
  NAND2_X1 U659 ( .A1(G91), .A2(n650), .ZN(n592) );
  NAND2_X1 U660 ( .A1(G78), .A2(n647), .ZN(n591) );
  NAND2_X1 U661 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U662 ( .A1(n594), .A2(n593), .ZN(n948) );
  XOR2_X1 U663 ( .A(n948), .B(KEYINPUT70), .Z(G299) );
  INV_X1 U664 ( .A(G868), .ZN(n670) );
  XNOR2_X1 U665 ( .A(KEYINPUT78), .B(n670), .ZN(n595) );
  NOR2_X1 U666 ( .A1(G286), .A2(n595), .ZN(n597) );
  NOR2_X1 U667 ( .A1(G868), .A2(G299), .ZN(n596) );
  NOR2_X1 U668 ( .A1(n597), .A2(n596), .ZN(G297) );
  NAND2_X1 U669 ( .A1(n598), .A2(G559), .ZN(n599) );
  NAND2_X1 U670 ( .A1(n599), .A2(n897), .ZN(n600) );
  XNOR2_X1 U671 ( .A(n600), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U672 ( .A1(G868), .A2(n696), .ZN(n601) );
  XOR2_X1 U673 ( .A(KEYINPUT79), .B(n601), .Z(n605) );
  NAND2_X1 U674 ( .A1(n897), .A2(G868), .ZN(n602) );
  XNOR2_X1 U675 ( .A(KEYINPUT80), .B(n602), .ZN(n603) );
  NOR2_X1 U676 ( .A1(G559), .A2(n603), .ZN(n604) );
  NOR2_X1 U677 ( .A1(n605), .A2(n604), .ZN(G282) );
  NAND2_X1 U678 ( .A1(G123), .A2(n876), .ZN(n606) );
  XOR2_X1 U679 ( .A(KEYINPUT81), .B(n606), .Z(n607) );
  XNOR2_X1 U680 ( .A(n607), .B(KEYINPUT18), .ZN(n609) );
  NAND2_X1 U681 ( .A1(G111), .A2(n877), .ZN(n608) );
  NAND2_X1 U682 ( .A1(n609), .A2(n608), .ZN(n613) );
  NAND2_X1 U683 ( .A1(G135), .A2(n870), .ZN(n611) );
  NAND2_X1 U684 ( .A1(G99), .A2(n872), .ZN(n610) );
  NAND2_X1 U685 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U686 ( .A1(n613), .A2(n612), .ZN(n921) );
  XNOR2_X1 U687 ( .A(n921), .B(G2096), .ZN(n614) );
  XNOR2_X1 U688 ( .A(n614), .B(KEYINPUT82), .ZN(n616) );
  INV_X1 U689 ( .A(G2100), .ZN(n615) );
  NAND2_X1 U690 ( .A1(n616), .A2(n615), .ZN(G156) );
  NAND2_X1 U691 ( .A1(G93), .A2(n650), .ZN(n618) );
  NAND2_X1 U692 ( .A1(G80), .A2(n647), .ZN(n617) );
  NAND2_X1 U693 ( .A1(n618), .A2(n617), .ZN(n621) );
  NAND2_X1 U694 ( .A1(G67), .A2(n649), .ZN(n619) );
  XNOR2_X1 U695 ( .A(KEYINPUT83), .B(n619), .ZN(n620) );
  NOR2_X1 U696 ( .A1(n621), .A2(n620), .ZN(n623) );
  NAND2_X1 U697 ( .A1(n653), .A2(G55), .ZN(n622) );
  NAND2_X1 U698 ( .A1(n623), .A2(n622), .ZN(n671) );
  NAND2_X1 U699 ( .A1(G559), .A2(n897), .ZN(n624) );
  XNOR2_X1 U700 ( .A(n624), .B(n696), .ZN(n667) );
  NOR2_X1 U701 ( .A1(G860), .A2(n667), .ZN(n625) );
  XOR2_X1 U702 ( .A(n671), .B(n625), .Z(G145) );
  NAND2_X1 U703 ( .A1(n649), .A2(G60), .ZN(n626) );
  XOR2_X1 U704 ( .A(KEYINPUT67), .B(n626), .Z(n628) );
  NAND2_X1 U705 ( .A1(n653), .A2(G47), .ZN(n627) );
  NAND2_X1 U706 ( .A1(n628), .A2(n627), .ZN(n629) );
  XOR2_X1 U707 ( .A(KEYINPUT68), .B(n629), .Z(n633) );
  NAND2_X1 U708 ( .A1(n647), .A2(G72), .ZN(n631) );
  NAND2_X1 U709 ( .A1(G85), .A2(n650), .ZN(n630) );
  AND2_X1 U710 ( .A1(n631), .A2(n630), .ZN(n632) );
  NAND2_X1 U711 ( .A1(n633), .A2(n632), .ZN(G290) );
  NAND2_X1 U712 ( .A1(G88), .A2(n650), .ZN(n635) );
  NAND2_X1 U713 ( .A1(G75), .A2(n647), .ZN(n634) );
  NAND2_X1 U714 ( .A1(n635), .A2(n634), .ZN(n639) );
  NAND2_X1 U715 ( .A1(G62), .A2(n649), .ZN(n637) );
  NAND2_X1 U716 ( .A1(G50), .A2(n653), .ZN(n636) );
  NAND2_X1 U717 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U718 ( .A1(n639), .A2(n638), .ZN(G166) );
  NAND2_X1 U719 ( .A1(G49), .A2(n653), .ZN(n640) );
  XNOR2_X1 U720 ( .A(n640), .B(KEYINPUT84), .ZN(n646) );
  NAND2_X1 U721 ( .A1(G87), .A2(n641), .ZN(n643) );
  NAND2_X1 U722 ( .A1(G74), .A2(G651), .ZN(n642) );
  NAND2_X1 U723 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U724 ( .A1(n649), .A2(n644), .ZN(n645) );
  NAND2_X1 U725 ( .A1(n646), .A2(n645), .ZN(G288) );
  NAND2_X1 U726 ( .A1(n647), .A2(G73), .ZN(n648) );
  XNOR2_X1 U727 ( .A(n648), .B(KEYINPUT2), .ZN(n658) );
  NAND2_X1 U728 ( .A1(G61), .A2(n649), .ZN(n652) );
  NAND2_X1 U729 ( .A1(G86), .A2(n650), .ZN(n651) );
  NAND2_X1 U730 ( .A1(n652), .A2(n651), .ZN(n656) );
  NAND2_X1 U731 ( .A1(G48), .A2(n653), .ZN(n654) );
  XNOR2_X1 U732 ( .A(KEYINPUT85), .B(n654), .ZN(n655) );
  NOR2_X1 U733 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U734 ( .A1(n658), .A2(n657), .ZN(G305) );
  XNOR2_X1 U735 ( .A(G299), .B(G290), .ZN(n666) );
  XOR2_X1 U736 ( .A(KEYINPUT19), .B(KEYINPUT88), .Z(n659) );
  XNOR2_X1 U737 ( .A(G288), .B(n659), .ZN(n660) );
  XNOR2_X1 U738 ( .A(KEYINPUT87), .B(n660), .ZN(n662) );
  XNOR2_X1 U739 ( .A(G305), .B(KEYINPUT86), .ZN(n661) );
  XNOR2_X1 U740 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U741 ( .A(G166), .B(n663), .ZN(n664) );
  XNOR2_X1 U742 ( .A(n664), .B(n671), .ZN(n665) );
  XNOR2_X1 U743 ( .A(n666), .B(n665), .ZN(n896) );
  XNOR2_X1 U744 ( .A(n896), .B(n667), .ZN(n668) );
  NAND2_X1 U745 ( .A1(n668), .A2(G868), .ZN(n669) );
  XOR2_X1 U746 ( .A(KEYINPUT89), .B(n669), .Z(n673) );
  NAND2_X1 U747 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U748 ( .A1(n673), .A2(n672), .ZN(G295) );
  NAND2_X1 U749 ( .A1(G2084), .A2(G2078), .ZN(n674) );
  XOR2_X1 U750 ( .A(KEYINPUT20), .B(n674), .Z(n675) );
  NAND2_X1 U751 ( .A1(n675), .A2(G2090), .ZN(n676) );
  XNOR2_X1 U752 ( .A(n676), .B(KEYINPUT90), .ZN(n677) );
  XNOR2_X1 U753 ( .A(KEYINPUT21), .B(n677), .ZN(n678) );
  NAND2_X1 U754 ( .A1(G2072), .A2(n678), .ZN(G158) );
  XNOR2_X1 U755 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U756 ( .A1(G220), .A2(G219), .ZN(n679) );
  XOR2_X1 U757 ( .A(KEYINPUT22), .B(n679), .Z(n680) );
  NOR2_X1 U758 ( .A1(G218), .A2(n680), .ZN(n681) );
  NAND2_X1 U759 ( .A1(G96), .A2(n681), .ZN(n829) );
  NAND2_X1 U760 ( .A1(n829), .A2(G2106), .ZN(n685) );
  NAND2_X1 U761 ( .A1(G69), .A2(G108), .ZN(n682) );
  NOR2_X1 U762 ( .A1(G236), .A2(n682), .ZN(n683) );
  NAND2_X1 U763 ( .A1(G57), .A2(n683), .ZN(n830) );
  NAND2_X1 U764 ( .A1(n830), .A2(G567), .ZN(n684) );
  NAND2_X1 U765 ( .A1(n685), .A2(n684), .ZN(n831) );
  NAND2_X1 U766 ( .A1(G483), .A2(G661), .ZN(n686) );
  NOR2_X1 U767 ( .A1(n831), .A2(n686), .ZN(n828) );
  NAND2_X1 U768 ( .A1(n828), .A2(G36), .ZN(G176) );
  INV_X1 U769 ( .A(G166), .ZN(G303) );
  NOR2_X1 U770 ( .A1(G2090), .A2(G303), .ZN(n687) );
  NAND2_X1 U771 ( .A1(G8), .A2(n687), .ZN(n752) );
  AND2_X1 U772 ( .A1(G160), .A2(G40), .ZN(n776) );
  NAND2_X1 U773 ( .A1(n778), .A2(n776), .ZN(n735) );
  NAND2_X1 U774 ( .A1(n735), .A2(G1348), .ZN(n691) );
  NAND2_X1 U775 ( .A1(G2067), .A2(n717), .ZN(n688) );
  XNOR2_X1 U776 ( .A(KEYINPUT95), .B(n688), .ZN(n689) );
  INV_X1 U777 ( .A(n689), .ZN(n690) );
  NAND2_X1 U778 ( .A1(n691), .A2(n690), .ZN(n698) );
  INV_X1 U779 ( .A(G1996), .ZN(n971) );
  NOR2_X1 U780 ( .A1(n735), .A2(n971), .ZN(n692) );
  XOR2_X1 U781 ( .A(n692), .B(KEYINPUT26), .Z(n694) );
  NAND2_X1 U782 ( .A1(n735), .A2(G1341), .ZN(n693) );
  NAND2_X1 U783 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U784 ( .A1(n700), .A2(n944), .ZN(n697) );
  NAND2_X1 U785 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U786 ( .A(n699), .B(KEYINPUT96), .ZN(n703) );
  NOR2_X1 U787 ( .A1(n944), .A2(n700), .ZN(n701) );
  XNOR2_X1 U788 ( .A(KEYINPUT97), .B(n701), .ZN(n702) );
  NAND2_X1 U789 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U790 ( .A(n704), .B(KEYINPUT98), .ZN(n709) );
  NAND2_X1 U791 ( .A1(n717), .A2(G2072), .ZN(n705) );
  XNOR2_X1 U792 ( .A(n705), .B(KEYINPUT27), .ZN(n707) );
  INV_X1 U793 ( .A(G1956), .ZN(n1008) );
  NOR2_X1 U794 ( .A1(n1008), .A2(n717), .ZN(n706) );
  NOR2_X1 U795 ( .A1(n707), .A2(n706), .ZN(n710) );
  NAND2_X1 U796 ( .A1(n710), .A2(n948), .ZN(n708) );
  NAND2_X1 U797 ( .A1(n709), .A2(n708), .ZN(n714) );
  NOR2_X1 U798 ( .A1(n710), .A2(n948), .ZN(n712) );
  XOR2_X1 U799 ( .A(KEYINPUT94), .B(KEYINPUT28), .Z(n711) );
  XNOR2_X1 U800 ( .A(n712), .B(n711), .ZN(n713) );
  NAND2_X1 U801 ( .A1(n714), .A2(n713), .ZN(n716) );
  XNOR2_X1 U802 ( .A(KEYINPUT99), .B(KEYINPUT29), .ZN(n715) );
  XNOR2_X1 U803 ( .A(n716), .B(n715), .ZN(n723) );
  XOR2_X1 U804 ( .A(G2078), .B(KEYINPUT25), .Z(n978) );
  INV_X1 U805 ( .A(n717), .ZN(n718) );
  NOR2_X1 U806 ( .A1(n978), .A2(n718), .ZN(n721) );
  NOR2_X1 U807 ( .A1(n719), .A2(G1961), .ZN(n720) );
  NOR2_X1 U808 ( .A1(n721), .A2(n720), .ZN(n724) );
  OR2_X1 U809 ( .A1(n724), .A2(G301), .ZN(n722) );
  NAND2_X1 U810 ( .A1(n723), .A2(n722), .ZN(n733) );
  NAND2_X1 U811 ( .A1(n724), .A2(G301), .ZN(n725) );
  XOR2_X1 U812 ( .A(KEYINPUT100), .B(n725), .Z(n730) );
  NAND2_X1 U813 ( .A1(G8), .A2(n735), .ZN(n774) );
  NOR2_X1 U814 ( .A1(G1966), .A2(n774), .ZN(n746) );
  NOR2_X1 U815 ( .A1(G2084), .A2(n735), .ZN(n747) );
  NOR2_X1 U816 ( .A1(n746), .A2(n747), .ZN(n726) );
  NAND2_X1 U817 ( .A1(G8), .A2(n726), .ZN(n727) );
  XNOR2_X1 U818 ( .A(KEYINPUT30), .B(n727), .ZN(n728) );
  NOR2_X1 U819 ( .A1(G168), .A2(n728), .ZN(n729) );
  NOR2_X1 U820 ( .A1(n730), .A2(n729), .ZN(n731) );
  XOR2_X1 U821 ( .A(KEYINPUT31), .B(n731), .Z(n732) );
  NAND2_X1 U822 ( .A1(n733), .A2(n732), .ZN(n744) );
  AND2_X1 U823 ( .A1(G286), .A2(G8), .ZN(n734) );
  NAND2_X1 U824 ( .A1(n744), .A2(n734), .ZN(n742) );
  INV_X1 U825 ( .A(G8), .ZN(n740) );
  NOR2_X1 U826 ( .A1(G1971), .A2(n774), .ZN(n737) );
  NOR2_X1 U827 ( .A1(G2090), .A2(n735), .ZN(n736) );
  NOR2_X1 U828 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U829 ( .A1(n738), .A2(G303), .ZN(n739) );
  OR2_X1 U830 ( .A1(n740), .A2(n739), .ZN(n741) );
  AND2_X1 U831 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U832 ( .A(n743), .B(KEYINPUT32), .ZN(n751) );
  XNOR2_X1 U833 ( .A(KEYINPUT101), .B(n744), .ZN(n745) );
  NOR2_X1 U834 ( .A1(n746), .A2(n745), .ZN(n749) );
  NAND2_X1 U835 ( .A1(G8), .A2(n747), .ZN(n748) );
  NAND2_X1 U836 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U837 ( .A1(n751), .A2(n750), .ZN(n757) );
  NAND2_X1 U838 ( .A1(n752), .A2(n757), .ZN(n753) );
  NAND2_X1 U839 ( .A1(n753), .A2(n774), .ZN(n770) );
  NOR2_X1 U840 ( .A1(G1976), .A2(G288), .ZN(n761) );
  NOR2_X1 U841 ( .A1(G1971), .A2(G303), .ZN(n754) );
  NOR2_X1 U842 ( .A1(n761), .A2(n754), .ZN(n952) );
  INV_X1 U843 ( .A(KEYINPUT33), .ZN(n755) );
  AND2_X1 U844 ( .A1(n952), .A2(n755), .ZN(n756) );
  NAND2_X1 U845 ( .A1(n757), .A2(n756), .ZN(n768) );
  INV_X1 U846 ( .A(n774), .ZN(n759) );
  NAND2_X1 U847 ( .A1(G288), .A2(G1976), .ZN(n758) );
  XNOR2_X1 U848 ( .A(n758), .B(KEYINPUT102), .ZN(n956) );
  AND2_X1 U849 ( .A1(n759), .A2(n956), .ZN(n760) );
  OR2_X1 U850 ( .A1(KEYINPUT33), .A2(n760), .ZN(n764) );
  NAND2_X1 U851 ( .A1(n761), .A2(KEYINPUT33), .ZN(n762) );
  OR2_X1 U852 ( .A1(n774), .A2(n762), .ZN(n763) );
  NAND2_X1 U853 ( .A1(n764), .A2(n763), .ZN(n766) );
  XOR2_X1 U854 ( .A(G1981), .B(G305), .Z(n961) );
  INV_X1 U855 ( .A(n961), .ZN(n765) );
  NOR2_X1 U856 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U857 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U858 ( .A1(n770), .A2(n769), .ZN(n771) );
  NOR2_X1 U859 ( .A1(G1981), .A2(G305), .ZN(n772) );
  XOR2_X1 U860 ( .A(n772), .B(KEYINPUT24), .Z(n773) );
  NAND2_X1 U861 ( .A1(n775), .A2(n516), .ZN(n806) );
  INV_X1 U862 ( .A(n776), .ZN(n777) );
  NOR2_X1 U863 ( .A1(n778), .A2(n777), .ZN(n820) );
  NAND2_X1 U864 ( .A1(G131), .A2(n870), .ZN(n780) );
  NAND2_X1 U865 ( .A1(G119), .A2(n876), .ZN(n779) );
  NAND2_X1 U866 ( .A1(n780), .A2(n779), .ZN(n784) );
  NAND2_X1 U867 ( .A1(G95), .A2(n872), .ZN(n782) );
  NAND2_X1 U868 ( .A1(G107), .A2(n877), .ZN(n781) );
  NAND2_X1 U869 ( .A1(n782), .A2(n781), .ZN(n783) );
  OR2_X1 U870 ( .A1(n784), .A2(n783), .ZN(n860) );
  NAND2_X1 U871 ( .A1(G1991), .A2(n860), .ZN(n794) );
  NAND2_X1 U872 ( .A1(G129), .A2(n876), .ZN(n786) );
  NAND2_X1 U873 ( .A1(G117), .A2(n877), .ZN(n785) );
  NAND2_X1 U874 ( .A1(n786), .A2(n785), .ZN(n789) );
  NAND2_X1 U875 ( .A1(n872), .A2(G105), .ZN(n787) );
  XOR2_X1 U876 ( .A(KEYINPUT38), .B(n787), .Z(n788) );
  NOR2_X1 U877 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U878 ( .A(n790), .B(KEYINPUT92), .ZN(n792) );
  NAND2_X1 U879 ( .A1(G141), .A2(n870), .ZN(n791) );
  NAND2_X1 U880 ( .A1(n792), .A2(n791), .ZN(n890) );
  NAND2_X1 U881 ( .A1(G1996), .A2(n890), .ZN(n793) );
  NAND2_X1 U882 ( .A1(n794), .A2(n793), .ZN(n939) );
  NAND2_X1 U883 ( .A1(n820), .A2(n939), .ZN(n808) );
  XOR2_X1 U884 ( .A(G1986), .B(KEYINPUT91), .Z(n795) );
  XNOR2_X1 U885 ( .A(G290), .B(n795), .ZN(n954) );
  NAND2_X1 U886 ( .A1(n820), .A2(n954), .ZN(n796) );
  NAND2_X1 U887 ( .A1(G140), .A2(n870), .ZN(n798) );
  NAND2_X1 U888 ( .A1(G104), .A2(n872), .ZN(n797) );
  NAND2_X1 U889 ( .A1(n798), .A2(n797), .ZN(n799) );
  XNOR2_X1 U890 ( .A(KEYINPUT34), .B(n799), .ZN(n804) );
  NAND2_X1 U891 ( .A1(G128), .A2(n876), .ZN(n801) );
  NAND2_X1 U892 ( .A1(G116), .A2(n877), .ZN(n800) );
  NAND2_X1 U893 ( .A1(n801), .A2(n800), .ZN(n802) );
  XOR2_X1 U894 ( .A(KEYINPUT35), .B(n802), .Z(n803) );
  NOR2_X1 U895 ( .A1(n804), .A2(n803), .ZN(n805) );
  XNOR2_X1 U896 ( .A(KEYINPUT36), .B(n805), .ZN(n893) );
  XNOR2_X1 U897 ( .A(G2067), .B(KEYINPUT37), .ZN(n817) );
  NOR2_X1 U898 ( .A1(n893), .A2(n817), .ZN(n926) );
  NAND2_X1 U899 ( .A1(n820), .A2(n926), .ZN(n815) );
  NAND2_X1 U900 ( .A1(n806), .A2(n517), .ZN(n807) );
  XNOR2_X1 U901 ( .A(n807), .B(KEYINPUT104), .ZN(n822) );
  XOR2_X1 U902 ( .A(KEYINPUT105), .B(KEYINPUT39), .Z(n814) );
  NOR2_X1 U903 ( .A1(G1996), .A2(n890), .ZN(n919) );
  INV_X1 U904 ( .A(n808), .ZN(n811) );
  NOR2_X1 U905 ( .A1(G1991), .A2(n860), .ZN(n922) );
  NOR2_X1 U906 ( .A1(G1986), .A2(G290), .ZN(n809) );
  NOR2_X1 U907 ( .A1(n922), .A2(n809), .ZN(n810) );
  NOR2_X1 U908 ( .A1(n811), .A2(n810), .ZN(n812) );
  NOR2_X1 U909 ( .A1(n919), .A2(n812), .ZN(n813) );
  XNOR2_X1 U910 ( .A(n814), .B(n813), .ZN(n816) );
  NAND2_X1 U911 ( .A1(n816), .A2(n815), .ZN(n818) );
  NAND2_X1 U912 ( .A1(n893), .A2(n817), .ZN(n927) );
  NAND2_X1 U913 ( .A1(n818), .A2(n927), .ZN(n819) );
  NAND2_X1 U914 ( .A1(n820), .A2(n819), .ZN(n821) );
  NAND2_X1 U915 ( .A1(n822), .A2(n821), .ZN(n823) );
  XNOR2_X1 U916 ( .A(n823), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U917 ( .A1(n824), .A2(G2106), .ZN(n825) );
  XOR2_X1 U918 ( .A(KEYINPUT107), .B(n825), .Z(G217) );
  AND2_X1 U919 ( .A1(G15), .A2(G2), .ZN(n826) );
  NAND2_X1 U920 ( .A1(G661), .A2(n826), .ZN(G259) );
  NAND2_X1 U921 ( .A1(G3), .A2(G1), .ZN(n827) );
  NAND2_X1 U922 ( .A1(n828), .A2(n827), .ZN(G188) );
  XOR2_X1 U923 ( .A(G69), .B(KEYINPUT108), .Z(G235) );
  XNOR2_X1 U924 ( .A(G108), .B(KEYINPUT117), .ZN(G238) );
  INV_X1 U926 ( .A(G96), .ZN(G221) );
  NOR2_X1 U927 ( .A1(n830), .A2(n829), .ZN(G325) );
  INV_X1 U928 ( .A(G325), .ZN(G261) );
  INV_X1 U929 ( .A(n831), .ZN(G319) );
  XOR2_X1 U930 ( .A(KEYINPUT109), .B(G2084), .Z(n833) );
  XNOR2_X1 U931 ( .A(G2067), .B(G2090), .ZN(n832) );
  XNOR2_X1 U932 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U933 ( .A(n834), .B(G2100), .Z(n836) );
  XNOR2_X1 U934 ( .A(G2072), .B(G2078), .ZN(n835) );
  XNOR2_X1 U935 ( .A(n836), .B(n835), .ZN(n840) );
  XOR2_X1 U936 ( .A(G2096), .B(G2678), .Z(n838) );
  XNOR2_X1 U937 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n837) );
  XNOR2_X1 U938 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U939 ( .A(n840), .B(n839), .Z(G227) );
  XNOR2_X1 U940 ( .A(G1966), .B(KEYINPUT110), .ZN(n850) );
  XOR2_X1 U941 ( .A(G1976), .B(G1971), .Z(n842) );
  XNOR2_X1 U942 ( .A(G1986), .B(G1961), .ZN(n841) );
  XNOR2_X1 U943 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U944 ( .A(G1956), .B(G1981), .Z(n844) );
  XNOR2_X1 U945 ( .A(G1996), .B(G1991), .ZN(n843) );
  XNOR2_X1 U946 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U947 ( .A(n846), .B(n845), .Z(n848) );
  XNOR2_X1 U948 ( .A(G2474), .B(KEYINPUT41), .ZN(n847) );
  XNOR2_X1 U949 ( .A(n848), .B(n847), .ZN(n849) );
  XNOR2_X1 U950 ( .A(n850), .B(n849), .ZN(G229) );
  NAND2_X1 U951 ( .A1(G112), .A2(n877), .ZN(n857) );
  NAND2_X1 U952 ( .A1(G136), .A2(n870), .ZN(n852) );
  NAND2_X1 U953 ( .A1(G100), .A2(n872), .ZN(n851) );
  NAND2_X1 U954 ( .A1(n852), .A2(n851), .ZN(n855) );
  NAND2_X1 U955 ( .A1(n876), .A2(G124), .ZN(n853) );
  XOR2_X1 U956 ( .A(KEYINPUT44), .B(n853), .Z(n854) );
  NOR2_X1 U957 ( .A1(n855), .A2(n854), .ZN(n856) );
  NAND2_X1 U958 ( .A1(n857), .A2(n856), .ZN(n858) );
  XNOR2_X1 U959 ( .A(n858), .B(KEYINPUT111), .ZN(G162) );
  XOR2_X1 U960 ( .A(G164), .B(n921), .Z(n859) );
  XNOR2_X1 U961 ( .A(n860), .B(n859), .ZN(n886) );
  NAND2_X1 U962 ( .A1(G130), .A2(n876), .ZN(n862) );
  NAND2_X1 U963 ( .A1(G118), .A2(n877), .ZN(n861) );
  NAND2_X1 U964 ( .A1(n862), .A2(n861), .ZN(n868) );
  NAND2_X1 U965 ( .A1(G142), .A2(n870), .ZN(n864) );
  NAND2_X1 U966 ( .A1(G106), .A2(n872), .ZN(n863) );
  NAND2_X1 U967 ( .A1(n864), .A2(n863), .ZN(n865) );
  XOR2_X1 U968 ( .A(KEYINPUT112), .B(n865), .Z(n866) );
  XNOR2_X1 U969 ( .A(KEYINPUT45), .B(n866), .ZN(n867) );
  NOR2_X1 U970 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U971 ( .A(n869), .B(G162), .Z(n884) );
  NAND2_X1 U972 ( .A1(G139), .A2(n870), .ZN(n871) );
  XNOR2_X1 U973 ( .A(n871), .B(KEYINPUT114), .ZN(n875) );
  NAND2_X1 U974 ( .A1(G103), .A2(n872), .ZN(n873) );
  XOR2_X1 U975 ( .A(KEYINPUT113), .B(n873), .Z(n874) );
  NAND2_X1 U976 ( .A1(n875), .A2(n874), .ZN(n882) );
  NAND2_X1 U977 ( .A1(G127), .A2(n876), .ZN(n879) );
  NAND2_X1 U978 ( .A1(G115), .A2(n877), .ZN(n878) );
  NAND2_X1 U979 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U980 ( .A(KEYINPUT47), .B(n880), .Z(n881) );
  NOR2_X1 U981 ( .A1(n882), .A2(n881), .ZN(n929) );
  XNOR2_X1 U982 ( .A(G160), .B(n929), .ZN(n883) );
  XNOR2_X1 U983 ( .A(n884), .B(n883), .ZN(n885) );
  XNOR2_X1 U984 ( .A(n886), .B(n885), .ZN(n892) );
  XOR2_X1 U985 ( .A(KEYINPUT116), .B(KEYINPUT46), .Z(n888) );
  XNOR2_X1 U986 ( .A(KEYINPUT115), .B(KEYINPUT48), .ZN(n887) );
  XNOR2_X1 U987 ( .A(n888), .B(n887), .ZN(n889) );
  XNOR2_X1 U988 ( .A(n890), .B(n889), .ZN(n891) );
  XNOR2_X1 U989 ( .A(n892), .B(n891), .ZN(n894) );
  XNOR2_X1 U990 ( .A(n894), .B(n893), .ZN(n895) );
  NOR2_X1 U991 ( .A1(G37), .A2(n895), .ZN(G395) );
  XOR2_X1 U992 ( .A(n896), .B(G286), .Z(n899) );
  XNOR2_X1 U993 ( .A(n897), .B(G171), .ZN(n898) );
  XNOR2_X1 U994 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U995 ( .A(n900), .B(n696), .ZN(n901) );
  NOR2_X1 U996 ( .A1(G37), .A2(n901), .ZN(G397) );
  XOR2_X1 U997 ( .A(G2443), .B(G2427), .Z(n903) );
  XNOR2_X1 U998 ( .A(G2438), .B(G2454), .ZN(n902) );
  XNOR2_X1 U999 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U1000 ( .A(n904), .B(G2435), .Z(n906) );
  XNOR2_X1 U1001 ( .A(G1341), .B(G1348), .ZN(n905) );
  XNOR2_X1 U1002 ( .A(n906), .B(n905), .ZN(n910) );
  XOR2_X1 U1003 ( .A(G2430), .B(G2446), .Z(n908) );
  XNOR2_X1 U1004 ( .A(KEYINPUT106), .B(G2451), .ZN(n907) );
  XNOR2_X1 U1005 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1006 ( .A(n910), .B(n909), .Z(n911) );
  NAND2_X1 U1007 ( .A1(G14), .A2(n911), .ZN(n917) );
  NAND2_X1 U1008 ( .A1(G319), .A2(n917), .ZN(n914) );
  NOR2_X1 U1009 ( .A1(G227), .A2(G229), .ZN(n912) );
  XNOR2_X1 U1010 ( .A(KEYINPUT49), .B(n912), .ZN(n913) );
  NOR2_X1 U1011 ( .A1(n914), .A2(n913), .ZN(n916) );
  NOR2_X1 U1012 ( .A1(G395), .A2(G397), .ZN(n915) );
  NAND2_X1 U1013 ( .A1(n916), .A2(n915), .ZN(G225) );
  INV_X1 U1014 ( .A(G225), .ZN(G308) );
  INV_X1 U1015 ( .A(G57), .ZN(G237) );
  INV_X1 U1016 ( .A(n917), .ZN(G401) );
  INV_X1 U1017 ( .A(KEYINPUT55), .ZN(n989) );
  XOR2_X1 U1018 ( .A(G2090), .B(G162), .Z(n918) );
  NOR2_X1 U1019 ( .A1(n919), .A2(n918), .ZN(n920) );
  XOR2_X1 U1020 ( .A(KEYINPUT51), .B(n920), .Z(n937) );
  XNOR2_X1 U1021 ( .A(G160), .B(G2084), .ZN(n924) );
  NOR2_X1 U1022 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n925) );
  NOR2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n928) );
  NAND2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n935) );
  XOR2_X1 U1026 ( .A(G2072), .B(n929), .Z(n931) );
  XOR2_X1 U1027 ( .A(G164), .B(G2078), .Z(n930) );
  NOR2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1029 ( .A(KEYINPUT118), .B(n932), .Z(n933) );
  XNOR2_X1 U1030 ( .A(KEYINPUT50), .B(n933), .ZN(n934) );
  NOR2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1032 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1033 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1034 ( .A(KEYINPUT52), .B(n940), .Z(n941) );
  XNOR2_X1 U1035 ( .A(KEYINPUT119), .B(n941), .ZN(n942) );
  NAND2_X1 U1036 ( .A1(n989), .A2(n942), .ZN(n943) );
  NAND2_X1 U1037 ( .A1(n943), .A2(G29), .ZN(n996) );
  XOR2_X1 U1038 ( .A(n944), .B(G1348), .Z(n946) );
  XNOR2_X1 U1039 ( .A(G301), .B(G1961), .ZN(n945) );
  NOR2_X1 U1040 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1041 ( .A(KEYINPUT122), .B(n947), .ZN(n960) );
  XNOR2_X1 U1042 ( .A(n1008), .B(n948), .ZN(n950) );
  AND2_X1 U1043 ( .A1(G1971), .A2(G303), .ZN(n949) );
  NOR2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1045 ( .A1(n952), .A2(n951), .ZN(n953) );
  NOR2_X1 U1046 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1047 ( .A1(n956), .A2(n955), .ZN(n958) );
  XNOR2_X1 U1048 ( .A(G1341), .B(n696), .ZN(n957) );
  NOR2_X1 U1049 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1050 ( .A1(n960), .A2(n959), .ZN(n965) );
  XNOR2_X1 U1051 ( .A(G1966), .B(G168), .ZN(n962) );
  NAND2_X1 U1052 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1053 ( .A(KEYINPUT57), .B(n963), .Z(n964) );
  NOR2_X1 U1054 ( .A1(n965), .A2(n964), .ZN(n967) );
  XOR2_X1 U1055 ( .A(G16), .B(KEYINPUT56), .Z(n966) );
  NOR2_X1 U1056 ( .A1(n967), .A2(n966), .ZN(n968) );
  XOR2_X1 U1057 ( .A(KEYINPUT123), .B(n968), .Z(n994) );
  XNOR2_X1 U1058 ( .A(G2090), .B(G35), .ZN(n984) );
  XNOR2_X1 U1059 ( .A(G1991), .B(G25), .ZN(n970) );
  XNOR2_X1 U1060 ( .A(G33), .B(G2072), .ZN(n969) );
  NOR2_X1 U1061 ( .A1(n970), .A2(n969), .ZN(n977) );
  XNOR2_X1 U1062 ( .A(G32), .B(n971), .ZN(n972) );
  NAND2_X1 U1063 ( .A1(n972), .A2(G28), .ZN(n975) );
  XNOR2_X1 U1064 ( .A(KEYINPUT120), .B(G2067), .ZN(n973) );
  XNOR2_X1 U1065 ( .A(G26), .B(n973), .ZN(n974) );
  NOR2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1067 ( .A1(n977), .A2(n976), .ZN(n981) );
  XOR2_X1 U1068 ( .A(G27), .B(n978), .Z(n979) );
  XNOR2_X1 U1069 ( .A(KEYINPUT121), .B(n979), .ZN(n980) );
  NOR2_X1 U1070 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1071 ( .A(KEYINPUT53), .B(n982), .ZN(n983) );
  NOR2_X1 U1072 ( .A1(n984), .A2(n983), .ZN(n987) );
  XOR2_X1 U1073 ( .A(G2084), .B(G34), .Z(n985) );
  XNOR2_X1 U1074 ( .A(KEYINPUT54), .B(n985), .ZN(n986) );
  NAND2_X1 U1075 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1076 ( .A(n989), .B(n988), .ZN(n991) );
  INV_X1 U1077 ( .A(G29), .ZN(n990) );
  NAND2_X1 U1078 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1079 ( .A1(G11), .A2(n992), .ZN(n993) );
  NOR2_X1 U1080 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1081 ( .A1(n996), .A2(n995), .ZN(n1023) );
  XOR2_X1 U1082 ( .A(G1986), .B(KEYINPUT126), .Z(n997) );
  XNOR2_X1 U1083 ( .A(G24), .B(n997), .ZN(n1001) );
  XNOR2_X1 U1084 ( .A(G1971), .B(G22), .ZN(n999) );
  XNOR2_X1 U1085 ( .A(G23), .B(G1976), .ZN(n998) );
  NOR2_X1 U1086 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1087 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1088 ( .A(n1002), .B(KEYINPUT58), .ZN(n1005) );
  XOR2_X1 U1089 ( .A(G1966), .B(G21), .Z(n1003) );
  XNOR2_X1 U1090 ( .A(KEYINPUT125), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1091 ( .A1(n1005), .A2(n1004), .ZN(n1017) );
  XOR2_X1 U1092 ( .A(G4), .B(KEYINPUT124), .Z(n1007) );
  XNOR2_X1 U1093 ( .A(G1348), .B(KEYINPUT59), .ZN(n1006) );
  XNOR2_X1 U1094 ( .A(n1007), .B(n1006), .ZN(n1014) );
  XNOR2_X1 U1095 ( .A(G20), .B(n1008), .ZN(n1012) );
  XNOR2_X1 U1096 ( .A(G1981), .B(G6), .ZN(n1010) );
  XNOR2_X1 U1097 ( .A(G19), .B(G1341), .ZN(n1009) );
  NOR2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NOR2_X1 U1100 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1101 ( .A(n1015), .B(KEYINPUT60), .ZN(n1016) );
  NAND2_X1 U1102 ( .A1(n1017), .A2(n1016), .ZN(n1019) );
  XNOR2_X1 U1103 ( .A(G5), .B(G1961), .ZN(n1018) );
  NOR2_X1 U1104 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XOR2_X1 U1105 ( .A(KEYINPUT61), .B(n1020), .Z(n1021) );
  NOR2_X1 U1106 ( .A1(G16), .A2(n1021), .ZN(n1022) );
  NOR2_X1 U1107 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1108 ( .A(KEYINPUT127), .B(n1024), .Z(n1025) );
  XNOR2_X1 U1109 ( .A(KEYINPUT62), .B(n1025), .ZN(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

