

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584;

  XOR2_X1 U322 ( .A(KEYINPUT97), .B(n529), .Z(n290) );
  AND2_X1 U323 ( .A1(G226GAT), .A2(G233GAT), .ZN(n291) );
  INV_X1 U324 ( .A(KEYINPUT15), .ZN(n401) );
  XNOR2_X1 U325 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U326 ( .A(n377), .B(n291), .ZN(n357) );
  XNOR2_X1 U327 ( .A(n404), .B(n403), .ZN(n407) );
  XNOR2_X1 U328 ( .A(n357), .B(n405), .ZN(n361) );
  XNOR2_X1 U329 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U330 ( .A(n412), .B(n411), .ZN(n413) );
  NOR2_X1 U331 ( .A1(n476), .A2(n475), .ZN(n560) );
  INV_X1 U332 ( .A(G43GAT), .ZN(n453) );
  XOR2_X1 U333 ( .A(n368), .B(n367), .Z(n522) );
  XNOR2_X1 U334 ( .A(n477), .B(G190GAT), .ZN(n478) );
  XNOR2_X1 U335 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U336 ( .A(n479), .B(n478), .ZN(G1351GAT) );
  XNOR2_X1 U337 ( .A(n456), .B(n455), .ZN(G1330GAT) );
  XOR2_X1 U338 ( .A(KEYINPUT83), .B(G183GAT), .Z(n293) );
  XNOR2_X1 U339 ( .A(G43GAT), .B(G134GAT), .ZN(n292) );
  XNOR2_X1 U340 ( .A(n293), .B(n292), .ZN(n297) );
  XOR2_X1 U341 ( .A(KEYINPUT88), .B(KEYINPUT85), .Z(n295) );
  XNOR2_X1 U342 ( .A(KEYINPUT84), .B(KEYINPUT20), .ZN(n294) );
  XNOR2_X1 U343 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U344 ( .A(n297), .B(n296), .Z(n302) );
  XOR2_X1 U345 ( .A(G71GAT), .B(G176GAT), .Z(n299) );
  NAND2_X1 U346 ( .A1(G227GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U347 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U348 ( .A(G113GAT), .B(n300), .ZN(n301) );
  XNOR2_X1 U349 ( .A(n302), .B(n301), .ZN(n312) );
  XOR2_X1 U350 ( .A(G15GAT), .B(G127GAT), .Z(n408) );
  XNOR2_X1 U351 ( .A(G120GAT), .B(KEYINPUT82), .ZN(n303) );
  XNOR2_X1 U352 ( .A(n303), .B(KEYINPUT0), .ZN(n347) );
  XOR2_X1 U353 ( .A(n408), .B(n347), .Z(n305) );
  XNOR2_X1 U354 ( .A(G190GAT), .B(G99GAT), .ZN(n304) );
  XNOR2_X1 U355 ( .A(n305), .B(n304), .ZN(n310) );
  XOR2_X1 U356 ( .A(KEYINPUT87), .B(KEYINPUT18), .Z(n307) );
  XNOR2_X1 U357 ( .A(G169GAT), .B(KEYINPUT86), .ZN(n306) );
  XNOR2_X1 U358 ( .A(n307), .B(n306), .ZN(n309) );
  XOR2_X1 U359 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n308) );
  XNOR2_X1 U360 ( .A(n309), .B(n308), .ZN(n367) );
  XOR2_X1 U361 ( .A(n310), .B(n367), .Z(n311) );
  XOR2_X1 U362 ( .A(n312), .B(n311), .Z(n530) );
  INV_X1 U363 ( .A(n530), .ZN(n476) );
  XNOR2_X1 U364 ( .A(KEYINPUT36), .B(KEYINPUT106), .ZN(n333) );
  XOR2_X1 U365 ( .A(KEYINPUT64), .B(KEYINPUT66), .Z(n314) );
  XNOR2_X1 U366 ( .A(KEYINPUT9), .B(KEYINPUT76), .ZN(n313) );
  XNOR2_X1 U367 ( .A(n314), .B(n313), .ZN(n332) );
  XOR2_X1 U368 ( .A(KEYINPUT11), .B(KEYINPUT65), .Z(n316) );
  XNOR2_X1 U369 ( .A(G92GAT), .B(KEYINPUT78), .ZN(n315) );
  XNOR2_X1 U370 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U371 ( .A(n317), .B(KEYINPUT10), .Z(n319) );
  XOR2_X1 U372 ( .A(G134GAT), .B(KEYINPUT77), .Z(n336) );
  XNOR2_X1 U373 ( .A(G106GAT), .B(n336), .ZN(n318) );
  XNOR2_X1 U374 ( .A(n319), .B(n318), .ZN(n325) );
  XOR2_X1 U375 ( .A(G99GAT), .B(G85GAT), .Z(n441) );
  XNOR2_X1 U376 ( .A(G29GAT), .B(G43GAT), .ZN(n321) );
  XNOR2_X1 U377 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n320) );
  XOR2_X1 U378 ( .A(n321), .B(n320), .Z(n429) );
  XNOR2_X1 U379 ( .A(n441), .B(n429), .ZN(n323) );
  AND2_X1 U380 ( .A1(G232GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U381 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U382 ( .A(n325), .B(n324), .Z(n330) );
  XOR2_X1 U383 ( .A(G162GAT), .B(KEYINPUT75), .Z(n327) );
  XNOR2_X1 U384 ( .A(G50GAT), .B(G218GAT), .ZN(n326) );
  XNOR2_X1 U385 ( .A(n327), .B(n326), .ZN(n370) );
  XNOR2_X1 U386 ( .A(G36GAT), .B(G190GAT), .ZN(n328) );
  XNOR2_X1 U387 ( .A(n328), .B(KEYINPUT79), .ZN(n364) );
  XNOR2_X1 U388 ( .A(n370), .B(n364), .ZN(n329) );
  XNOR2_X1 U389 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U390 ( .A(n332), .B(n331), .ZN(n555) );
  XNOR2_X1 U391 ( .A(n333), .B(n555), .ZN(n581) );
  XOR2_X1 U392 ( .A(KEYINPUT90), .B(KEYINPUT6), .Z(n335) );
  XNOR2_X1 U393 ( .A(KEYINPUT5), .B(KEYINPUT91), .ZN(n334) );
  XNOR2_X1 U394 ( .A(n335), .B(n334), .ZN(n355) );
  XOR2_X1 U395 ( .A(G85GAT), .B(n336), .Z(n338) );
  XOR2_X1 U396 ( .A(G113GAT), .B(G1GAT), .Z(n428) );
  XNOR2_X1 U397 ( .A(n428), .B(G162GAT), .ZN(n337) );
  XNOR2_X1 U398 ( .A(n338), .B(n337), .ZN(n351) );
  XOR2_X1 U399 ( .A(G148GAT), .B(G155GAT), .Z(n340) );
  XNOR2_X1 U400 ( .A(G29GAT), .B(G127GAT), .ZN(n339) );
  XNOR2_X1 U401 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U402 ( .A(KEYINPUT92), .B(KEYINPUT4), .Z(n342) );
  XNOR2_X1 U403 ( .A(G57GAT), .B(KEYINPUT1), .ZN(n341) );
  XNOR2_X1 U404 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U405 ( .A(n344), .B(n343), .Z(n349) );
  XOR2_X1 U406 ( .A(KEYINPUT2), .B(KEYINPUT89), .Z(n346) );
  XNOR2_X1 U407 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n345) );
  XNOR2_X1 U408 ( .A(n346), .B(n345), .ZN(n382) );
  XNOR2_X1 U409 ( .A(n347), .B(n382), .ZN(n348) );
  XNOR2_X1 U410 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U411 ( .A(n351), .B(n350), .Z(n353) );
  NAND2_X1 U412 ( .A1(G225GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U413 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U414 ( .A(n355), .B(n354), .ZN(n520) );
  INV_X1 U415 ( .A(n520), .ZN(n496) );
  XOR2_X1 U416 ( .A(G197GAT), .B(KEYINPUT21), .Z(n377) );
  XNOR2_X1 U417 ( .A(G8GAT), .B(G183GAT), .ZN(n356) );
  XNOR2_X1 U418 ( .A(n356), .B(G211GAT), .ZN(n405) );
  XOR2_X1 U419 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n359) );
  XNOR2_X1 U420 ( .A(G218GAT), .B(KEYINPUT95), .ZN(n358) );
  XNOR2_X1 U421 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U422 ( .A(n361), .B(n360), .Z(n366) );
  XOR2_X1 U423 ( .A(G64GAT), .B(G92GAT), .Z(n363) );
  XNOR2_X1 U424 ( .A(G176GAT), .B(G204GAT), .ZN(n362) );
  XNOR2_X1 U425 ( .A(n363), .B(n362), .ZN(n446) );
  XNOR2_X1 U426 ( .A(n364), .B(n446), .ZN(n365) );
  XNOR2_X1 U427 ( .A(n366), .B(n365), .ZN(n368) );
  XOR2_X1 U428 ( .A(n522), .B(KEYINPUT96), .Z(n369) );
  XNOR2_X1 U429 ( .A(n369), .B(KEYINPUT27), .ZN(n390) );
  NOR2_X1 U430 ( .A1(n496), .A2(n390), .ZN(n544) );
  XOR2_X1 U431 ( .A(KEYINPUT22), .B(n370), .Z(n372) );
  NAND2_X1 U432 ( .A1(G228GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U433 ( .A(n372), .B(n371), .ZN(n376) );
  XOR2_X1 U434 ( .A(G204GAT), .B(G211GAT), .Z(n374) );
  XNOR2_X1 U435 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n373) );
  XNOR2_X1 U436 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U437 ( .A(n376), .B(n375), .Z(n379) );
  XOR2_X1 U438 ( .A(G22GAT), .B(G155GAT), .Z(n400) );
  XNOR2_X1 U439 ( .A(n377), .B(n400), .ZN(n378) );
  XNOR2_X1 U440 ( .A(n379), .B(n378), .ZN(n384) );
  XOR2_X1 U441 ( .A(G78GAT), .B(G148GAT), .Z(n381) );
  XNOR2_X1 U442 ( .A(G106GAT), .B(KEYINPUT73), .ZN(n380) );
  XNOR2_X1 U443 ( .A(n381), .B(n380), .ZN(n447) );
  XOR2_X1 U444 ( .A(n382), .B(n447), .Z(n383) );
  XNOR2_X1 U445 ( .A(n384), .B(n383), .ZN(n473) );
  XNOR2_X1 U446 ( .A(KEYINPUT28), .B(n473), .ZN(n525) );
  INV_X1 U447 ( .A(n525), .ZN(n503) );
  NAND2_X1 U448 ( .A1(n544), .A2(n503), .ZN(n529) );
  NOR2_X1 U449 ( .A1(n530), .A2(n290), .ZN(n395) );
  INV_X1 U450 ( .A(n522), .ZN(n499) );
  NOR2_X1 U451 ( .A1(n476), .A2(n499), .ZN(n385) );
  NOR2_X1 U452 ( .A1(n473), .A2(n385), .ZN(n386) );
  XNOR2_X1 U453 ( .A(n386), .B(KEYINPUT99), .ZN(n387) );
  XNOR2_X1 U454 ( .A(n387), .B(KEYINPUT25), .ZN(n392) );
  NAND2_X1 U455 ( .A1(n473), .A2(n476), .ZN(n388) );
  XNOR2_X1 U456 ( .A(n388), .B(KEYINPUT26), .ZN(n389) );
  XNOR2_X1 U457 ( .A(KEYINPUT98), .B(n389), .ZN(n570) );
  NOR2_X1 U458 ( .A1(n390), .A2(n570), .ZN(n391) );
  NOR2_X1 U459 ( .A1(n392), .A2(n391), .ZN(n393) );
  NOR2_X1 U460 ( .A1(n520), .A2(n393), .ZN(n394) );
  NOR2_X1 U461 ( .A1(n395), .A2(n394), .ZN(n396) );
  XNOR2_X1 U462 ( .A(n396), .B(KEYINPUT100), .ZN(n484) );
  XOR2_X1 U463 ( .A(KEYINPUT14), .B(KEYINPUT80), .Z(n398) );
  XNOR2_X1 U464 ( .A(G1GAT), .B(KEYINPUT12), .ZN(n397) );
  XNOR2_X1 U465 ( .A(n398), .B(n397), .ZN(n414) );
  XNOR2_X1 U466 ( .A(G71GAT), .B(G57GAT), .ZN(n399) );
  XNOR2_X1 U467 ( .A(n399), .B(KEYINPUT13), .ZN(n444) );
  XNOR2_X1 U468 ( .A(n444), .B(n400), .ZN(n404) );
  AND2_X1 U469 ( .A1(G231GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U470 ( .A(n405), .B(KEYINPUT81), .ZN(n406) );
  XNOR2_X1 U471 ( .A(n407), .B(n406), .ZN(n412) );
  XNOR2_X1 U472 ( .A(n408), .B(G78GAT), .ZN(n410) );
  INV_X1 U473 ( .A(G64GAT), .ZN(n409) );
  XNOR2_X1 U474 ( .A(n414), .B(n413), .ZN(n579) );
  NOR2_X1 U475 ( .A1(n484), .A2(n579), .ZN(n415) );
  XNOR2_X1 U476 ( .A(n415), .B(KEYINPUT107), .ZN(n416) );
  NOR2_X1 U477 ( .A1(n581), .A2(n416), .ZN(n417) );
  XNOR2_X1 U478 ( .A(n417), .B(KEYINPUT37), .ZN(n519) );
  XOR2_X1 U479 ( .A(KEYINPUT70), .B(KEYINPUT69), .Z(n419) );
  XNOR2_X1 U480 ( .A(KEYINPUT29), .B(KEYINPUT68), .ZN(n418) );
  XNOR2_X1 U481 ( .A(n419), .B(n418), .ZN(n437) );
  XOR2_X1 U482 ( .A(G197GAT), .B(G141GAT), .Z(n421) );
  XNOR2_X1 U483 ( .A(G50GAT), .B(G36GAT), .ZN(n420) );
  XNOR2_X1 U484 ( .A(n421), .B(n420), .ZN(n425) );
  XOR2_X1 U485 ( .A(G8GAT), .B(G15GAT), .Z(n423) );
  XNOR2_X1 U486 ( .A(G169GAT), .B(G22GAT), .ZN(n422) );
  XNOR2_X1 U487 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U488 ( .A(n425), .B(n424), .Z(n435) );
  XOR2_X1 U489 ( .A(KEYINPUT30), .B(KEYINPUT71), .Z(n427) );
  XNOR2_X1 U490 ( .A(KEYINPUT72), .B(KEYINPUT67), .ZN(n426) );
  XNOR2_X1 U491 ( .A(n427), .B(n426), .ZN(n433) );
  XOR2_X1 U492 ( .A(n429), .B(n428), .Z(n431) );
  NAND2_X1 U493 ( .A1(G229GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U494 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U495 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U496 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U497 ( .A(n437), .B(n436), .Z(n545) );
  INV_X1 U498 ( .A(n545), .ZN(n572) );
  XOR2_X1 U499 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n439) );
  XNOR2_X1 U500 ( .A(G120GAT), .B(KEYINPUT32), .ZN(n438) );
  XNOR2_X1 U501 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U502 ( .A(n441), .B(n440), .Z(n443) );
  NAND2_X1 U503 ( .A1(G230GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U504 ( .A(n443), .B(n442), .ZN(n445) );
  XOR2_X1 U505 ( .A(n445), .B(n444), .Z(n449) );
  XNOR2_X1 U506 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U507 ( .A(n449), .B(n448), .ZN(n575) );
  NAND2_X1 U508 ( .A1(n572), .A2(n575), .ZN(n450) );
  XNOR2_X1 U509 ( .A(n450), .B(KEYINPUT74), .ZN(n485) );
  NOR2_X1 U510 ( .A1(n519), .A2(n485), .ZN(n452) );
  XOR2_X1 U511 ( .A(KEYINPUT38), .B(KEYINPUT108), .Z(n451) );
  XNOR2_X1 U512 ( .A(n452), .B(n451), .ZN(n502) );
  NOR2_X1 U513 ( .A1(n476), .A2(n502), .ZN(n456) );
  XNOR2_X1 U514 ( .A(KEYINPUT40), .B(KEYINPUT110), .ZN(n454) );
  XNOR2_X1 U515 ( .A(n575), .B(KEYINPUT41), .ZN(n559) );
  NAND2_X1 U516 ( .A1(n559), .A2(n572), .ZN(n459) );
  XOR2_X1 U517 ( .A(KEYINPUT118), .B(KEYINPUT46), .Z(n457) );
  XNOR2_X1 U518 ( .A(KEYINPUT117), .B(n457), .ZN(n458) );
  XNOR2_X1 U519 ( .A(n459), .B(n458), .ZN(n460) );
  XOR2_X1 U520 ( .A(n579), .B(KEYINPUT116), .Z(n565) );
  NAND2_X1 U521 ( .A1(n460), .A2(n565), .ZN(n461) );
  XNOR2_X1 U522 ( .A(n461), .B(KEYINPUT119), .ZN(n462) );
  NAND2_X1 U523 ( .A1(n462), .A2(n555), .ZN(n463) );
  XNOR2_X1 U524 ( .A(n463), .B(KEYINPUT47), .ZN(n469) );
  INV_X1 U525 ( .A(n579), .ZN(n552) );
  NOR2_X1 U526 ( .A1(n552), .A2(n581), .ZN(n464) );
  XNOR2_X1 U527 ( .A(KEYINPUT45), .B(n464), .ZN(n465) );
  NAND2_X1 U528 ( .A1(n465), .A2(n575), .ZN(n466) );
  XNOR2_X1 U529 ( .A(KEYINPUT120), .B(n466), .ZN(n467) );
  NOR2_X1 U530 ( .A1(n572), .A2(n467), .ZN(n468) );
  NOR2_X1 U531 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U532 ( .A(n470), .B(KEYINPUT48), .ZN(n542) );
  NOR2_X1 U533 ( .A1(n499), .A2(n542), .ZN(n471) );
  XNOR2_X1 U534 ( .A(n471), .B(KEYINPUT54), .ZN(n472) );
  NAND2_X1 U535 ( .A1(n472), .A2(n496), .ZN(n569) );
  NOR2_X1 U536 ( .A1(n473), .A2(n569), .ZN(n474) );
  XNOR2_X1 U537 ( .A(n474), .B(KEYINPUT55), .ZN(n475) );
  INV_X1 U538 ( .A(n560), .ZN(n564) );
  NOR2_X1 U539 ( .A1(n555), .A2(n564), .ZN(n479) );
  XNOR2_X1 U540 ( .A(KEYINPUT125), .B(KEYINPUT58), .ZN(n477) );
  XNOR2_X1 U541 ( .A(G1GAT), .B(KEYINPUT102), .ZN(n480) );
  XNOR2_X1 U542 ( .A(n480), .B(KEYINPUT34), .ZN(n481) );
  XOR2_X1 U543 ( .A(KEYINPUT101), .B(n481), .Z(n487) );
  NAND2_X1 U544 ( .A1(n555), .A2(n579), .ZN(n482) );
  XNOR2_X1 U545 ( .A(KEYINPUT16), .B(n482), .ZN(n483) );
  OR2_X1 U546 ( .A1(n484), .A2(n483), .ZN(n506) );
  NOR2_X1 U547 ( .A1(n485), .A2(n506), .ZN(n493) );
  NAND2_X1 U548 ( .A1(n493), .A2(n520), .ZN(n486) );
  XNOR2_X1 U549 ( .A(n487), .B(n486), .ZN(G1324GAT) );
  NAND2_X1 U550 ( .A1(n522), .A2(n493), .ZN(n488) );
  XNOR2_X1 U551 ( .A(n488), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U552 ( .A(KEYINPUT35), .B(KEYINPUT104), .Z(n490) );
  NAND2_X1 U553 ( .A1(n493), .A2(n530), .ZN(n489) );
  XNOR2_X1 U554 ( .A(n490), .B(n489), .ZN(n492) );
  XOR2_X1 U555 ( .A(G15GAT), .B(KEYINPUT103), .Z(n491) );
  XNOR2_X1 U556 ( .A(n492), .B(n491), .ZN(G1326GAT) );
  XOR2_X1 U557 ( .A(G22GAT), .B(KEYINPUT105), .Z(n495) );
  NAND2_X1 U558 ( .A1(n493), .A2(n525), .ZN(n494) );
  XNOR2_X1 U559 ( .A(n495), .B(n494), .ZN(G1327GAT) );
  NOR2_X1 U560 ( .A1(n496), .A2(n502), .ZN(n498) );
  XNOR2_X1 U561 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n497) );
  XNOR2_X1 U562 ( .A(n498), .B(n497), .ZN(G1328GAT) );
  NOR2_X1 U563 ( .A1(n499), .A2(n502), .ZN(n501) );
  XNOR2_X1 U564 ( .A(G36GAT), .B(KEYINPUT109), .ZN(n500) );
  XNOR2_X1 U565 ( .A(n501), .B(n500), .ZN(G1329GAT) );
  NOR2_X1 U566 ( .A1(n503), .A2(n502), .ZN(n504) );
  XOR2_X1 U567 ( .A(G50GAT), .B(n504), .Z(G1331GAT) );
  XOR2_X1 U568 ( .A(KEYINPUT42), .B(KEYINPUT113), .Z(n509) );
  NAND2_X1 U569 ( .A1(n559), .A2(n545), .ZN(n505) );
  XOR2_X1 U570 ( .A(KEYINPUT111), .B(n505), .Z(n518) );
  NOR2_X1 U571 ( .A1(n518), .A2(n506), .ZN(n507) );
  XNOR2_X1 U572 ( .A(KEYINPUT112), .B(n507), .ZN(n515) );
  NAND2_X1 U573 ( .A1(n515), .A2(n520), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U575 ( .A(G57GAT), .B(n510), .ZN(G1332GAT) );
  NAND2_X1 U576 ( .A1(n515), .A2(n522), .ZN(n511) );
  XNOR2_X1 U577 ( .A(n511), .B(KEYINPUT114), .ZN(n512) );
  XNOR2_X1 U578 ( .A(G64GAT), .B(n512), .ZN(G1333GAT) );
  XOR2_X1 U579 ( .A(G71GAT), .B(KEYINPUT115), .Z(n514) );
  NAND2_X1 U580 ( .A1(n515), .A2(n530), .ZN(n513) );
  XNOR2_X1 U581 ( .A(n514), .B(n513), .ZN(G1334GAT) );
  XOR2_X1 U582 ( .A(G78GAT), .B(KEYINPUT43), .Z(n517) );
  NAND2_X1 U583 ( .A1(n525), .A2(n515), .ZN(n516) );
  XNOR2_X1 U584 ( .A(n517), .B(n516), .ZN(G1335GAT) );
  NOR2_X1 U585 ( .A1(n519), .A2(n518), .ZN(n526) );
  NAND2_X1 U586 ( .A1(n520), .A2(n526), .ZN(n521) );
  XNOR2_X1 U587 ( .A(n521), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U588 ( .A1(n526), .A2(n522), .ZN(n523) );
  XNOR2_X1 U589 ( .A(G92GAT), .B(n523), .ZN(G1337GAT) );
  NAND2_X1 U590 ( .A1(n530), .A2(n526), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n524), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U592 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n527), .B(KEYINPUT44), .ZN(n528) );
  XNOR2_X1 U594 ( .A(G106GAT), .B(n528), .ZN(G1339GAT) );
  NOR2_X1 U595 ( .A1(n542), .A2(n529), .ZN(n531) );
  NAND2_X1 U596 ( .A1(n531), .A2(n530), .ZN(n538) );
  NOR2_X1 U597 ( .A1(n545), .A2(n538), .ZN(n532) );
  XOR2_X1 U598 ( .A(G113GAT), .B(n532), .Z(G1340GAT) );
  INV_X1 U599 ( .A(n559), .ZN(n547) );
  NOR2_X1 U600 ( .A1(n547), .A2(n538), .ZN(n534) );
  XNOR2_X1 U601 ( .A(KEYINPUT121), .B(KEYINPUT49), .ZN(n533) );
  XNOR2_X1 U602 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U603 ( .A(G120GAT), .B(n535), .Z(G1341GAT) );
  NOR2_X1 U604 ( .A1(n565), .A2(n538), .ZN(n536) );
  XOR2_X1 U605 ( .A(KEYINPUT50), .B(n536), .Z(n537) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(n537), .ZN(G1342GAT) );
  NOR2_X1 U607 ( .A1(n555), .A2(n538), .ZN(n540) );
  XNOR2_X1 U608 ( .A(KEYINPUT51), .B(KEYINPUT122), .ZN(n539) );
  XNOR2_X1 U609 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U610 ( .A(G134GAT), .B(n541), .ZN(G1343GAT) );
  NOR2_X1 U611 ( .A1(n542), .A2(n570), .ZN(n543) );
  NAND2_X1 U612 ( .A1(n544), .A2(n543), .ZN(n554) );
  NOR2_X1 U613 ( .A1(n545), .A2(n554), .ZN(n546) );
  XOR2_X1 U614 ( .A(G141GAT), .B(n546), .Z(G1344GAT) );
  NOR2_X1 U615 ( .A1(n554), .A2(n547), .ZN(n551) );
  XOR2_X1 U616 ( .A(KEYINPUT123), .B(KEYINPUT52), .Z(n549) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n548) );
  XNOR2_X1 U618 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U619 ( .A(n551), .B(n550), .ZN(G1345GAT) );
  NOR2_X1 U620 ( .A1(n552), .A2(n554), .ZN(n553) );
  XOR2_X1 U621 ( .A(G155GAT), .B(n553), .Z(G1346GAT) );
  NOR2_X1 U622 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U623 ( .A(G162GAT), .B(n556), .Z(G1347GAT) );
  NAND2_X1 U624 ( .A1(n572), .A2(n560), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n557), .B(KEYINPUT124), .ZN(n558) );
  XNOR2_X1 U626 ( .A(G169GAT), .B(n558), .ZN(G1348GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n562) );
  NAND2_X1 U628 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U630 ( .A(G176GAT), .B(n563), .ZN(G1349GAT) );
  NOR2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U632 ( .A(G183GAT), .B(n566), .Z(G1350GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT127), .B(KEYINPUT59), .Z(n568) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(n574) );
  NOR2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U637 ( .A(n571), .B(KEYINPUT126), .Z(n582) );
  INV_X1 U638 ( .A(n582), .ZN(n578) );
  NAND2_X1 U639 ( .A1(n578), .A2(n572), .ZN(n573) );
  XOR2_X1 U640 ( .A(n574), .B(n573), .Z(G1352GAT) );
  XOR2_X1 U641 ( .A(G204GAT), .B(KEYINPUT61), .Z(n577) );
  OR2_X1 U642 ( .A1(n582), .A2(n575), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  NAND2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(G211GAT), .B(n580), .ZN(G1354GAT) );
  NOR2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U647 ( .A(KEYINPUT62), .B(n583), .Z(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

