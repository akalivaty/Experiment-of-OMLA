//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 1 0 0 1 1 0 0 0 1 0 1 1 1 1 0 0 1 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 1 0 0 0 0 0 0 1 1 0 1 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n811, new_n812, new_n813,
    new_n815, new_n816, new_n817, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947;
  INV_X1    g000(.A(G71gat), .ZN(new_n202));
  INV_X1    g001(.A(G78gat), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n202), .A2(new_n203), .A3(KEYINPUT9), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(new_n202), .B2(new_n203), .ZN(new_n205));
  INV_X1    g004(.A(G57gat), .ZN(new_n206));
  INV_X1    g005(.A(G64gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(G57gat), .A2(G64gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n205), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  AND2_X1   g009(.A1(G57gat), .A2(G64gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(G57gat), .A2(G64gat), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT95), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT95), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n208), .A2(new_n214), .A3(new_n209), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n213), .A2(new_n215), .A3(KEYINPUT9), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT96), .ZN(new_n217));
  XOR2_X1   g016(.A(G71gat), .B(G78gat), .Z(new_n218));
  AND3_X1   g017(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n217), .B1(new_n216), .B2(new_n218), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n210), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT21), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(G231gat), .A2(G233gat), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n223), .B(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G127gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n225), .B(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT91), .ZN(new_n228));
  INV_X1    g027(.A(G15gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n229), .A2(G22gat), .ZN(new_n230));
  INV_X1    g029(.A(G22gat), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n231), .A2(G15gat), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n228), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(G15gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n229), .A2(G22gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n234), .A2(new_n235), .A3(KEYINPUT91), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(G1gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(KEYINPUT16), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n239), .B(KEYINPUT92), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n233), .A2(new_n238), .A3(new_n236), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(G8gat), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n244), .B1(new_n242), .B2(KEYINPUT93), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  OAI211_X1 g045(.A(new_n241), .B(new_n242), .C1(KEYINPUT93), .C2(new_n244), .ZN(new_n247));
  AND2_X1   g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n248), .B1(new_n222), .B2(new_n221), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n227), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n251), .B(KEYINPUT97), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n252), .B(G155gat), .ZN(new_n253));
  XOR2_X1   g052(.A(G183gat), .B(G211gat), .Z(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  OR2_X1    g054(.A1(new_n250), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n250), .A2(new_n255), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(G29gat), .A2(G36gat), .ZN(new_n260));
  INV_X1    g059(.A(G43gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(G50gat), .ZN(new_n262));
  INV_X1    g061(.A(G50gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(G43gat), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n262), .A2(new_n264), .A3(KEYINPUT15), .ZN(new_n265));
  OAI21_X1  g064(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n266));
  NOR3_X1   g065(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n266), .B1(new_n267), .B2(KEYINPUT90), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT14), .ZN(new_n269));
  INV_X1    g068(.A(G29gat), .ZN(new_n270));
  INV_X1    g069(.A(G36gat), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT90), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n260), .B(new_n265), .C1(new_n268), .C2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT88), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n276), .B1(new_n261), .B2(G50gat), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n263), .A2(KEYINPUT88), .A3(G43gat), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n277), .A2(new_n262), .A3(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT89), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT15), .ZN(new_n281));
  AND3_X1   g080(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n280), .B1(new_n279), .B2(new_n281), .ZN(new_n283));
  OR3_X1    g082(.A1(new_n275), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  AOI22_X1  g083(.A1(new_n272), .A2(new_n266), .B1(G29gat), .B2(G36gat), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n285), .A2(new_n265), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n284), .A2(KEYINPUT17), .A3(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT17), .ZN(new_n289));
  NOR3_X1   g088(.A1(new_n275), .A2(new_n282), .A3(new_n283), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n289), .B1(new_n290), .B2(new_n286), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n248), .A2(new_n288), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(G229gat), .A2(G233gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n284), .A2(new_n287), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n246), .A2(new_n247), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n292), .A2(new_n293), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT18), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n292), .A2(KEYINPUT18), .A3(new_n293), .A4(new_n296), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n294), .B(new_n295), .ZN(new_n301));
  XOR2_X1   g100(.A(new_n293), .B(KEYINPUT13), .Z(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n299), .A2(new_n300), .A3(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G113gat), .B(G141gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n305), .B(G197gat), .ZN(new_n306));
  XOR2_X1   g105(.A(KEYINPUT11), .B(G169gat), .Z(new_n307));
  XNOR2_X1  g106(.A(new_n306), .B(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n308), .B(KEYINPUT12), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n304), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT94), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n299), .A2(new_n309), .A3(new_n303), .A4(new_n300), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n304), .A2(KEYINPUT94), .A3(new_n310), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G99gat), .B(G106gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(G85gat), .A2(G92gat), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT7), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n318), .A2(KEYINPUT98), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(G85gat), .ZN(new_n321));
  INV_X1    g120(.A(G92gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(G99gat), .A2(G106gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT8), .ZN(new_n325));
  AND3_X1   g124(.A1(new_n320), .A2(new_n323), .A3(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT98), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT7), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n319), .A2(KEYINPUT98), .ZN(new_n329));
  AND2_X1   g128(.A1(G85gat), .A2(G92gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n317), .B1(new_n326), .B2(new_n331), .ZN(new_n332));
  AOI22_X1  g131(.A1(KEYINPUT8), .A2(new_n324), .B1(new_n321), .B2(new_n322), .ZN(new_n333));
  AND4_X1   g132(.A1(new_n317), .A2(new_n331), .A3(new_n320), .A4(new_n333), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n221), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT10), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n335), .B(new_n210), .C1(new_n220), .C2(new_n219), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n216), .A2(new_n218), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT96), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n344), .A2(KEYINPUT10), .A3(new_n210), .A4(new_n335), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n340), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G230gat), .A2(G233gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AND2_X1   g147(.A1(new_n337), .A2(new_n339), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n348), .B1(new_n349), .B2(new_n347), .ZN(new_n350));
  XOR2_X1   g149(.A(G120gat), .B(G148gat), .Z(new_n351));
  XNOR2_X1  g150(.A(new_n351), .B(KEYINPUT100), .ZN(new_n352));
  XNOR2_X1  g151(.A(G176gat), .B(G204gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n352), .B(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  OR2_X1    g154(.A1(new_n350), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n350), .A2(new_n355), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT99), .ZN(new_n359));
  AND2_X1   g158(.A1(G232gat), .A2(G233gat), .ZN(new_n360));
  AOI22_X1  g159(.A1(new_n294), .A2(new_n335), .B1(KEYINPUT41), .B2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n288), .A2(new_n291), .A3(new_n336), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n359), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n361), .A2(new_n362), .A3(new_n359), .ZN(new_n365));
  XNOR2_X1  g164(.A(G134gat), .B(G162gat), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  AND3_X1   g166(.A1(new_n364), .A2(new_n365), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n367), .B1(new_n364), .B2(new_n365), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n360), .A2(KEYINPUT41), .ZN(new_n370));
  XNOR2_X1  g169(.A(G190gat), .B(G218gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n370), .B(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  OR3_X1    g172(.A1(new_n368), .A2(new_n369), .A3(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n373), .B1(new_n368), .B2(new_n369), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NOR4_X1   g175(.A1(new_n259), .A2(new_n316), .A3(new_n358), .A4(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(G155gat), .ZN(new_n378));
  INV_X1    g177(.A(G162gat), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g179(.A1(G155gat), .A2(G162gat), .ZN(new_n381));
  XOR2_X1   g180(.A(G141gat), .B(G148gat), .Z(new_n382));
  XNOR2_X1  g181(.A(KEYINPUT75), .B(KEYINPUT2), .ZN(new_n383));
  AOI211_X1 g182(.A(new_n380), .B(new_n381), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(G148gat), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n385), .A2(G141gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(KEYINPUT76), .B(G148gat), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n386), .B1(new_n387), .B2(G141gat), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT2), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n380), .B1(new_n389), .B2(new_n381), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n384), .A2(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(G197gat), .B(G204gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(G211gat), .A2(G218gat), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT22), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n394), .A2(KEYINPUT73), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT73), .B1(new_n394), .B2(new_n395), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(G211gat), .B(G218gat), .ZN(new_n400));
  OR2_X1    g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n399), .A2(new_n400), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT82), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT29), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n405), .B(new_n406), .C1(KEYINPUT82), .C2(new_n401), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT3), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n392), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  AND2_X1   g208(.A1(G228gat), .A2(G233gat), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n392), .A2(new_n408), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n403), .B1(new_n411), .B2(new_n406), .ZN(new_n412));
  OR3_X1    g211(.A1(new_n409), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n412), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT3), .B1(new_n403), .B2(new_n406), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n414), .B1(new_n392), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(new_n410), .ZN(new_n417));
  XNOR2_X1  g216(.A(KEYINPUT31), .B(G50gat), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n413), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(G78gat), .B(G106gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n421), .B(G22gat), .ZN(new_n422));
  NOR3_X1   g221(.A1(new_n409), .A2(new_n410), .A3(new_n412), .ZN(new_n423));
  INV_X1    g222(.A(new_n417), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n418), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AND3_X1   g224(.A1(new_n420), .A2(new_n422), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n422), .B1(new_n420), .B2(new_n425), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(G113gat), .B(G120gat), .ZN(new_n429));
  OR2_X1    g228(.A1(new_n429), .A2(KEYINPUT1), .ZN(new_n430));
  XNOR2_X1  g229(.A(G127gat), .B(G134gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n430), .B(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n392), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n432), .A2(new_n392), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(G225gat), .A2(G233gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n439), .B(KEYINPUT77), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(KEYINPUT5), .B1(new_n438), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n434), .A2(KEYINPUT3), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n444), .A2(new_n433), .A3(new_n411), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT4), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n436), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n432), .A2(new_n392), .A3(KEYINPUT4), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n445), .A2(new_n441), .A3(new_n447), .A4(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT78), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n443), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n442), .A2(KEYINPUT78), .A3(new_n449), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XOR2_X1   g252(.A(G1gat), .B(G29gat), .Z(new_n454));
  XNOR2_X1  g253(.A(new_n454), .B(KEYINPUT80), .ZN(new_n455));
  XOR2_X1   g254(.A(G57gat), .B(G85gat), .Z(new_n456));
  XNOR2_X1  g255(.A(new_n455), .B(new_n456), .ZN(new_n457));
  XNOR2_X1  g256(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n457), .B(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT6), .B1(new_n453), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n459), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT83), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT83), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n459), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n451), .A2(new_n465), .A3(new_n452), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n460), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n451), .A2(new_n452), .A3(KEYINPUT6), .A4(new_n461), .ZN(new_n468));
  XNOR2_X1  g267(.A(KEYINPUT27), .B(G183gat), .ZN(new_n469));
  INV_X1    g268(.A(G190gat), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n469), .A2(KEYINPUT28), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT27), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT27), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n474), .A2(KEYINPUT65), .A3(G183gat), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n473), .A2(new_n475), .A3(new_n470), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT66), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n473), .A2(new_n475), .A3(KEYINPUT66), .A4(new_n470), .ZN(new_n479));
  XNOR2_X1  g278(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n471), .B1(new_n478), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT26), .ZN(new_n483));
  INV_X1    g282(.A(G169gat), .ZN(new_n484));
  INV_X1    g283(.A(G176gat), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n487));
  NAND2_X1  g286(.A1(G169gat), .A2(G176gat), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(G183gat), .A2(G190gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n482), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n484), .A2(new_n485), .A3(KEYINPUT23), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT23), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n495), .B1(G169gat), .B2(G176gat), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT24), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n497), .A2(G183gat), .A3(G190gat), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n494), .A2(new_n496), .A3(new_n498), .A4(new_n488), .ZN(new_n499));
  AND2_X1   g298(.A1(G183gat), .A2(G190gat), .ZN(new_n500));
  NOR2_X1   g299(.A1(G183gat), .A2(G190gat), .ZN(new_n501));
  NOR3_X1   g300(.A1(new_n500), .A2(new_n501), .A3(new_n497), .ZN(new_n502));
  OAI21_X1  g301(.A(KEYINPUT64), .B1(new_n499), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT25), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT25), .ZN(new_n505));
  OAI211_X1 g304(.A(KEYINPUT64), .B(new_n505), .C1(new_n499), .C2(new_n502), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n493), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n508), .A2(G226gat), .A3(G233gat), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  AOI22_X1  g309(.A1(new_n508), .A2(new_n406), .B1(G226gat), .B2(G233gat), .ZN(new_n511));
  NOR3_X1   g310(.A1(new_n510), .A2(new_n511), .A3(new_n404), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n404), .B1(new_n510), .B2(new_n511), .ZN(new_n514));
  XNOR2_X1  g313(.A(G8gat), .B(G36gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(G64gat), .B(G92gat), .ZN(new_n516));
  XOR2_X1   g315(.A(new_n515), .B(new_n516), .Z(new_n517));
  NAND3_X1  g316(.A1(new_n513), .A2(new_n514), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n467), .A2(new_n468), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n513), .A2(KEYINPUT74), .A3(new_n514), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT74), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n508), .A2(new_n406), .ZN(new_n522));
  INV_X1    g321(.A(G226gat), .ZN(new_n523));
  INV_X1    g322(.A(G233gat), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n403), .B1(new_n525), .B2(new_n509), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n521), .B1(new_n526), .B2(new_n512), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n520), .A2(KEYINPUT37), .A3(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n517), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT87), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(KEYINPUT85), .B(KEYINPUT38), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT37), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n513), .A2(new_n535), .A3(new_n514), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(KEYINPUT86), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n528), .A2(KEYINPUT87), .A3(new_n529), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n532), .A2(new_n534), .A3(new_n537), .A4(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n513), .A2(new_n514), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n517), .B1(new_n540), .B2(KEYINPUT37), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(new_n533), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n519), .B1(new_n539), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n445), .A2(new_n447), .A3(new_n448), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT39), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n545), .A2(new_n546), .A3(new_n440), .ZN(new_n547));
  AND3_X1   g346(.A1(new_n462), .A2(new_n464), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n545), .A2(new_n440), .ZN(new_n549));
  OAI211_X1 g348(.A(new_n549), .B(KEYINPUT39), .C1(new_n440), .C2(new_n437), .ZN(new_n550));
  AND2_X1   g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  OR2_X1    g350(.A1(new_n551), .A2(KEYINPUT40), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n548), .A2(KEYINPUT40), .A3(new_n550), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT84), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n548), .A2(KEYINPUT84), .A3(KEYINPUT40), .A4(new_n550), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT30), .ZN(new_n558));
  OR2_X1    g357(.A1(new_n518), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n520), .A2(new_n529), .A3(new_n527), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n518), .A2(new_n558), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  AND4_X1   g361(.A1(new_n466), .A2(new_n552), .A3(new_n557), .A4(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n428), .B1(new_n544), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n428), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT81), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n566), .B1(new_n453), .B2(new_n459), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n451), .A2(new_n452), .A3(KEYINPUT81), .A4(new_n461), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n567), .A2(new_n460), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n562), .B1(new_n569), .B2(new_n468), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n565), .A2(new_n570), .ZN(new_n571));
  AOI22_X1  g370(.A1(new_n500), .A2(new_n497), .B1(G169gat), .B2(G176gat), .ZN(new_n572));
  OR2_X1    g371(.A1(G183gat), .A2(G190gat), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n573), .A2(KEYINPUT24), .A3(new_n490), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n572), .A2(new_n574), .A3(new_n496), .A4(new_n494), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n505), .B1(new_n575), .B2(KEYINPUT64), .ZN(new_n576));
  INV_X1    g375(.A(new_n506), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n476), .A2(new_n477), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n579), .A2(new_n480), .A3(new_n479), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n491), .B1(new_n580), .B2(new_n471), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n433), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n493), .A2(new_n507), .A3(new_n432), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(G227gat), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n585), .A2(new_n524), .ZN(new_n586));
  AOI21_X1  g385(.A(KEYINPUT68), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT68), .ZN(new_n588));
  INV_X1    g387(.A(new_n586), .ZN(new_n589));
  AOI211_X1 g388(.A(new_n588), .B(new_n589), .C1(new_n582), .C2(new_n583), .ZN(new_n590));
  OAI21_X1  g389(.A(KEYINPUT32), .B1(new_n587), .B2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G15gat), .B(G43gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(G71gat), .B(G99gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n591), .B1(KEYINPUT33), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  AND3_X1   g396(.A1(new_n493), .A2(new_n432), .A3(new_n507), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n432), .B1(new_n493), .B2(new_n507), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n586), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(new_n588), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n584), .A2(KEYINPUT68), .A3(new_n586), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n594), .B1(new_n603), .B2(KEYINPUT32), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT33), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n605), .B1(new_n587), .B2(new_n590), .ZN(new_n606));
  AOI21_X1  g405(.A(KEYINPUT69), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  AND4_X1   g406(.A1(KEYINPUT69), .A2(new_n591), .A3(new_n606), .A4(new_n595), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n597), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n582), .A2(new_n589), .A3(new_n583), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT34), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n591), .A2(new_n606), .A3(new_n595), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT69), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n604), .A2(KEYINPUT69), .A3(new_n606), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n611), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n617), .A2(new_n618), .A3(new_n597), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n612), .A2(KEYINPUT36), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(KEYINPUT70), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT70), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n612), .A2(new_n622), .A3(KEYINPUT36), .A4(new_n619), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT72), .ZN(new_n625));
  AOI211_X1 g424(.A(new_n625), .B(new_n618), .C1(new_n617), .C2(new_n597), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n612), .A2(new_n625), .A3(new_n619), .ZN(new_n628));
  XNOR2_X1  g427(.A(KEYINPUT71), .B(KEYINPUT36), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  AOI22_X1  g429(.A1(new_n564), .A2(new_n571), .B1(new_n624), .B2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT35), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n467), .A2(new_n468), .ZN(new_n633));
  INV_X1    g432(.A(new_n562), .ZN(new_n634));
  AND4_X1   g433(.A1(new_n632), .A2(new_n428), .A3(new_n633), .A4(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n627), .A2(new_n628), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n618), .B1(new_n617), .B2(new_n597), .ZN(new_n637));
  AOI211_X1 g436(.A(new_n611), .B(new_n596), .C1(new_n615), .C2(new_n616), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n639), .A2(new_n428), .A3(new_n570), .ZN(new_n640));
  AOI22_X1  g439(.A1(new_n635), .A2(new_n636), .B1(new_n640), .B2(KEYINPUT35), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n377), .B1(new_n631), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n569), .A2(new_n468), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(KEYINPUT101), .B(G1gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(G1324gat));
  INV_X1    g445(.A(new_n642), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n244), .B1(new_n647), .B2(new_n562), .ZN(new_n648));
  XNOR2_X1  g447(.A(KEYINPUT16), .B(G8gat), .ZN(new_n649));
  NOR3_X1   g448(.A1(new_n642), .A2(new_n634), .A3(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(KEYINPUT42), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n651), .B1(KEYINPUT42), .B2(new_n650), .ZN(G1325gat));
  NAND3_X1  g451(.A1(new_n647), .A2(new_n229), .A3(new_n636), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n624), .A2(new_n630), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT102), .ZN(new_n655));
  OAI21_X1  g454(.A(G15gat), .B1(new_n655), .B2(new_n642), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n653), .A2(new_n656), .ZN(G1326gat));
  NOR2_X1   g456(.A1(new_n642), .A2(new_n428), .ZN(new_n658));
  XOR2_X1   g457(.A(KEYINPUT43), .B(G22gat), .Z(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(G1327gat));
  OAI21_X1  g459(.A(new_n376), .B1(new_n631), .B2(new_n641), .ZN(new_n661));
  NOR3_X1   g460(.A1(new_n258), .A2(new_n316), .A3(new_n358), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n643), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n664), .A2(new_n270), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(KEYINPUT45), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT44), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n661), .A2(new_n668), .ZN(new_n669));
  OAI211_X1 g468(.A(KEYINPUT44), .B(new_n376), .C1(new_n631), .C2(new_n641), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g470(.A(new_n662), .B(KEYINPUT103), .Z(new_n672));
  AND3_X1   g471(.A1(new_n671), .A2(new_n665), .A3(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n667), .B1(new_n270), .B2(new_n673), .ZN(G1328gat));
  NAND3_X1  g473(.A1(new_n664), .A2(new_n271), .A3(new_n562), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(KEYINPUT46), .ZN(new_n676));
  OR2_X1    g475(.A1(new_n675), .A2(KEYINPUT46), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n671), .A2(new_n562), .A3(new_n672), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(KEYINPUT104), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(G36gat), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n678), .A2(KEYINPUT104), .ZN(new_n681));
  OAI211_X1 g480(.A(new_n676), .B(new_n677), .C1(new_n680), .C2(new_n681), .ZN(G1329gat));
  AOI21_X1  g481(.A(new_n626), .B1(new_n639), .B2(new_n625), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n683), .A2(G43gat), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n664), .A2(new_n684), .ZN(new_n685));
  AOI22_X1  g484(.A1(new_n683), .A2(new_n629), .B1(new_n621), .B2(new_n623), .ZN(new_n686));
  AND3_X1   g485(.A1(new_n671), .A2(new_n686), .A3(new_n672), .ZN(new_n687));
  OAI211_X1 g486(.A(KEYINPUT47), .B(new_n685), .C1(new_n687), .C2(new_n261), .ZN(new_n688));
  INV_X1    g487(.A(new_n655), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n671), .A2(new_n689), .A3(new_n672), .ZN(new_n690));
  AOI22_X1  g489(.A1(new_n690), .A2(G43gat), .B1(new_n664), .B2(new_n684), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n688), .B1(new_n691), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g491(.A(KEYINPUT48), .ZN(new_n693));
  NOR4_X1   g492(.A1(new_n661), .A2(G50gat), .A3(new_n428), .A4(new_n663), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT106), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n693), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n669), .A2(new_n565), .A3(new_n670), .A4(new_n672), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(G50gat), .ZN(new_n698));
  OAI211_X1 g497(.A(new_n696), .B(new_n698), .C1(new_n695), .C2(new_n694), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT105), .ZN(new_n700));
  AND3_X1   g499(.A1(new_n697), .A2(new_n700), .A3(G50gat), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n700), .B1(new_n697), .B2(G50gat), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n701), .A2(new_n702), .A3(new_n694), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n699), .B1(new_n703), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g503(.A1(new_n631), .A2(new_n641), .ZN(new_n705));
  INV_X1    g504(.A(new_n376), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n258), .A2(new_n316), .A3(new_n358), .A4(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(new_n665), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g509(.A1(new_n708), .A2(KEYINPUT107), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT107), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n712), .B1(new_n705), .B2(new_n707), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n634), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n711), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(KEYINPUT108), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT108), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n711), .A2(new_n717), .A3(new_n713), .A4(new_n714), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n719), .B(new_n720), .ZN(G1333gat));
  AND3_X1   g520(.A1(new_n708), .A2(KEYINPUT109), .A3(new_n636), .ZN(new_n722));
  AOI21_X1  g521(.A(KEYINPUT109), .B1(new_n708), .B2(new_n636), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n202), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n711), .A2(new_n689), .A3(new_n713), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(G71gat), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT50), .ZN(new_n727));
  AND3_X1   g526(.A1(new_n724), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n727), .B1(new_n724), .B2(new_n726), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n728), .A2(new_n729), .ZN(G1334gat));
  NAND3_X1  g529(.A1(new_n711), .A2(new_n565), .A3(new_n713), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(G78gat), .ZN(G1335gat));
  INV_X1    g531(.A(new_n316), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n258), .A2(new_n733), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n376), .B(new_n734), .C1(new_n631), .C2(new_n641), .ZN(new_n735));
  NAND2_X1  g534(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XOR2_X1   g536(.A(KEYINPUT110), .B(KEYINPUT51), .Z(new_n738));
  OAI21_X1  g537(.A(new_n737), .B1(new_n735), .B2(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n665), .A2(new_n321), .A3(new_n358), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT111), .ZN(new_n741));
  INV_X1    g540(.A(new_n734), .ZN(new_n742));
  INV_X1    g541(.A(new_n358), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n669), .A2(new_n665), .A3(new_n670), .A4(new_n744), .ZN(new_n745));
  AOI22_X1  g544(.A1(new_n739), .A2(new_n741), .B1(new_n745), .B2(G85gat), .ZN(new_n746));
  XOR2_X1   g545(.A(new_n746), .B(KEYINPUT112), .Z(G1336gat));
  NAND4_X1  g546(.A1(new_n669), .A2(new_n562), .A3(new_n670), .A4(new_n744), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(G92gat), .ZN(new_n749));
  AOI21_X1  g548(.A(KEYINPUT52), .B1(new_n749), .B2(KEYINPUT114), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n562), .A2(new_n322), .A3(new_n358), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT113), .ZN(new_n752));
  AOI22_X1  g551(.A1(new_n739), .A2(new_n752), .B1(new_n748), .B2(G92gat), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n750), .B(new_n753), .ZN(G1337gat));
  NAND3_X1  g553(.A1(new_n671), .A2(new_n689), .A3(new_n744), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(G99gat), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n683), .A2(G99gat), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n739), .A2(new_n358), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(G1338gat));
  NOR2_X1   g558(.A1(new_n428), .A2(G106gat), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n739), .A2(new_n358), .A3(new_n760), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n669), .A2(new_n565), .A3(new_n670), .A4(new_n744), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(G106gat), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g564(.A(KEYINPUT54), .ZN(new_n766));
  INV_X1    g565(.A(new_n347), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n345), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n766), .B1(new_n768), .B2(new_n340), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n348), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n767), .B1(new_n340), .B2(new_n345), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n354), .B1(new_n771), .B2(new_n766), .ZN(new_n772));
  AOI211_X1 g571(.A(KEYINPUT116), .B(KEYINPUT55), .C1(new_n770), .C2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT116), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n346), .A2(new_n766), .A3(new_n347), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n345), .A2(new_n767), .ZN(new_n777));
  OAI21_X1  g576(.A(KEYINPUT54), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n775), .B(new_n355), .C1(new_n778), .C2(new_n771), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT55), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n774), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OR2_X1    g580(.A1(new_n773), .A2(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(KEYINPUT55), .B1(new_n778), .B2(new_n771), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n775), .A2(new_n355), .ZN(new_n784));
  OAI21_X1  g583(.A(KEYINPUT115), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT115), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n770), .A2(new_n772), .A3(new_n786), .A4(KEYINPUT55), .ZN(new_n787));
  AND3_X1   g586(.A1(new_n356), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n782), .A2(new_n788), .A3(new_n315), .A4(new_n314), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n301), .A2(new_n302), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n293), .B1(new_n292), .B2(new_n296), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n308), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n313), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n358), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n376), .B1(new_n789), .B2(new_n794), .ZN(new_n795));
  AND4_X1   g594(.A1(new_n376), .A2(new_n782), .A3(new_n793), .A4(new_n788), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n259), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n258), .A2(new_n316), .A3(new_n743), .A4(new_n706), .ZN(new_n798));
  AOI211_X1 g597(.A(new_n683), .B(new_n565), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n643), .A2(new_n562), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  XOR2_X1   g600(.A(new_n801), .B(KEYINPUT117), .Z(new_n802));
  NAND3_X1  g601(.A1(new_n802), .A2(G113gat), .A3(new_n733), .ZN(new_n803));
  INV_X1    g602(.A(G113gat), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n797), .A2(new_n798), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n639), .A2(new_n428), .ZN(new_n806));
  AND3_X1   g605(.A1(new_n805), .A2(new_n665), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n634), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n804), .B1(new_n808), .B2(new_n316), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n803), .A2(new_n809), .ZN(G1340gat));
  NAND3_X1  g609(.A1(new_n802), .A2(G120gat), .A3(new_n358), .ZN(new_n811));
  INV_X1    g610(.A(G120gat), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n812), .B1(new_n808), .B2(new_n743), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n811), .A2(new_n813), .ZN(G1341gat));
  INV_X1    g613(.A(new_n802), .ZN(new_n815));
  OAI21_X1  g614(.A(G127gat), .B1(new_n815), .B2(new_n259), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n258), .A2(new_n226), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n816), .B1(new_n808), .B2(new_n817), .ZN(G1342gat));
  OAI21_X1  g617(.A(G134gat), .B1(new_n815), .B2(new_n706), .ZN(new_n819));
  INV_X1    g618(.A(G134gat), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n706), .A2(new_n562), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n807), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  XOR2_X1   g621(.A(new_n822), .B(KEYINPUT56), .Z(new_n823));
  NAND2_X1  g622(.A1(new_n819), .A2(new_n823), .ZN(G1343gat));
  INV_X1    g623(.A(new_n800), .ZN(new_n825));
  OAI21_X1  g624(.A(KEYINPUT118), .B1(new_n686), .B2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT118), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n654), .A2(new_n827), .A3(new_n800), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n779), .A2(new_n780), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n788), .A2(new_n315), .A3(new_n314), .A4(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n376), .B1(new_n832), .B2(new_n794), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n259), .B1(new_n833), .B2(new_n796), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n798), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT57), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n428), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n428), .B1(new_n797), .B2(new_n798), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n838), .B1(new_n839), .B2(KEYINPUT57), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n830), .A2(new_n733), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT58), .B1(new_n841), .B2(G141gat), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n643), .B1(new_n797), .B2(new_n798), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n655), .A2(new_n565), .A3(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT121), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n844), .B(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n634), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n316), .A2(G141gat), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n842), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(new_n837), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n851), .B1(new_n834), .B2(new_n798), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n773), .A2(new_n781), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n356), .A2(new_n785), .A3(new_n787), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n316), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n794), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n706), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n853), .A2(new_n854), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(new_n376), .A3(new_n793), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n258), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n798), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n565), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n852), .B1(new_n862), .B2(new_n836), .ZN(new_n863));
  OAI21_X1  g662(.A(KEYINPUT119), .B1(new_n829), .B2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT119), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n840), .A2(new_n865), .A3(new_n826), .A4(new_n828), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n864), .A2(new_n733), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(G141gat), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n848), .A2(new_n634), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n844), .A2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(KEYINPUT120), .B1(new_n872), .B2(KEYINPUT58), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n870), .B1(new_n867), .B2(G141gat), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT120), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT58), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n850), .B1(new_n873), .B2(new_n877), .ZN(G1344gat));
  NAND2_X1  g677(.A1(new_n830), .A2(new_n358), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n858), .A2(new_n376), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT122), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n858), .A2(KEYINPUT122), .A3(new_n376), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n882), .A2(new_n793), .A3(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(new_n833), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n258), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n565), .B1(new_n886), .B2(new_n861), .ZN(new_n887));
  AOI22_X1  g686(.A1(new_n887), .A2(new_n836), .B1(new_n805), .B2(new_n837), .ZN(new_n888));
  OAI211_X1 g687(.A(KEYINPUT59), .B(G148gat), .C1(new_n879), .C2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n358), .A2(new_n387), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n864), .A2(new_n866), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n891), .A2(new_n743), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n892), .A2(new_n387), .ZN(new_n893));
  OAI221_X1 g692(.A(new_n889), .B1(new_n847), .B2(new_n890), .C1(new_n893), .C2(KEYINPUT59), .ZN(G1345gat));
  OAI21_X1  g693(.A(G155gat), .B1(new_n891), .B2(new_n259), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n258), .A2(new_n378), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n895), .B1(new_n847), .B2(new_n896), .ZN(G1346gat));
  NAND3_X1  g696(.A1(new_n846), .A2(new_n379), .A3(new_n821), .ZN(new_n898));
  OAI21_X1  g697(.A(G162gat), .B1(new_n891), .B2(new_n706), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(G1347gat));
  NOR2_X1   g699(.A1(new_n665), .A2(new_n634), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n799), .A2(new_n901), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n902), .A2(new_n484), .A3(new_n316), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n806), .A2(new_n562), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n904), .B(KEYINPUT123), .ZN(new_n905));
  AND3_X1   g704(.A1(new_n905), .A2(new_n643), .A3(new_n805), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(new_n733), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n903), .B1(new_n907), .B2(new_n484), .ZN(new_n908));
  XOR2_X1   g707(.A(new_n908), .B(KEYINPUT124), .Z(G1348gat));
  AOI21_X1  g708(.A(G176gat), .B1(new_n906), .B2(new_n358), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n910), .B(KEYINPUT125), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n902), .A2(new_n485), .A3(new_n743), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n911), .A2(new_n912), .ZN(G1349gat));
  NAND3_X1  g712(.A1(new_n906), .A2(new_n469), .A3(new_n258), .ZN(new_n914));
  OAI21_X1  g713(.A(G183gat), .B1(new_n902), .B2(new_n259), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g715(.A(KEYINPUT126), .B(KEYINPUT60), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n916), .B(new_n917), .ZN(G1350gat));
  OAI21_X1  g717(.A(G190gat), .B1(new_n902), .B2(new_n706), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT61), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n906), .A2(new_n470), .A3(new_n376), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1351gat));
  NAND2_X1  g721(.A1(new_n655), .A2(new_n901), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(new_n839), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(G197gat), .B1(new_n926), .B2(new_n733), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n923), .A2(new_n888), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n733), .A2(G197gat), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(G1352gat));
  NOR3_X1   g729(.A1(new_n925), .A2(G204gat), .A3(new_n743), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT62), .ZN(new_n932));
  OR2_X1    g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(new_n928), .ZN(new_n934));
  OAI21_X1  g733(.A(G204gat), .B1(new_n934), .B2(new_n743), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n931), .A2(new_n932), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n933), .A2(new_n935), .A3(new_n936), .ZN(G1353gat));
  OR3_X1    g736(.A1(new_n925), .A2(G211gat), .A3(new_n259), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n928), .A2(new_n258), .ZN(new_n939));
  AND3_X1   g738(.A1(new_n939), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n940));
  AOI21_X1  g739(.A(KEYINPUT63), .B1(new_n939), .B2(G211gat), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n938), .B1(new_n940), .B2(new_n941), .ZN(G1354gat));
  OAI21_X1  g741(.A(new_n376), .B1(new_n934), .B2(KEYINPUT127), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT127), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n928), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g744(.A(G218gat), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  OR2_X1    g745(.A1(new_n706), .A2(G218gat), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n946), .B1(new_n925), .B2(new_n947), .ZN(G1355gat));
endmodule


