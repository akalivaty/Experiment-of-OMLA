

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U546 ( .A1(G29), .A2(n1014), .ZN(n512) );
  INV_X1 U547 ( .A(KEYINPUT100), .ZN(n708) );
  INV_X1 U548 ( .A(KEYINPUT28), .ZN(n710) );
  NOR2_X1 U549 ( .A1(G651), .A2(n618), .ZN(n638) );
  NOR2_X2 U550 ( .A1(G2104), .A2(n515), .ZN(n891) );
  INV_X1 U551 ( .A(G2105), .ZN(n515) );
  NAND2_X1 U552 ( .A1(n515), .A2(G2104), .ZN(n513) );
  XNOR2_X1 U553 ( .A(n513), .B(KEYINPUT65), .ZN(n537) );
  NAND2_X1 U554 ( .A1(G101), .A2(n537), .ZN(n514) );
  XOR2_X1 U555 ( .A(KEYINPUT23), .B(n514), .Z(n517) );
  NAND2_X1 U556 ( .A1(n891), .A2(G125), .ZN(n516) );
  AND2_X1 U557 ( .A1(n517), .A2(n516), .ZN(n523) );
  AND2_X1 U558 ( .A1(G2105), .A2(G2104), .ZN(n890) );
  NAND2_X1 U559 ( .A1(G113), .A2(n890), .ZN(n521) );
  NOR2_X1 U560 ( .A1(G2105), .A2(G2104), .ZN(n518) );
  XOR2_X1 U561 ( .A(KEYINPUT17), .B(n518), .Z(n519) );
  XNOR2_X1 U562 ( .A(n519), .B(KEYINPUT66), .ZN(n543) );
  NAND2_X1 U563 ( .A1(G137), .A2(n543), .ZN(n520) );
  AND2_X1 U564 ( .A1(n521), .A2(n520), .ZN(n522) );
  AND2_X1 U565 ( .A1(n523), .A2(n522), .ZN(G160) );
  INV_X1 U566 ( .A(G651), .ZN(n527) );
  NOR2_X1 U567 ( .A1(G543), .A2(n527), .ZN(n524) );
  XOR2_X1 U568 ( .A(KEYINPUT1), .B(n524), .Z(n637) );
  NAND2_X1 U569 ( .A1(G64), .A2(n637), .ZN(n526) );
  XOR2_X1 U570 ( .A(KEYINPUT0), .B(G543), .Z(n618) );
  NAND2_X1 U571 ( .A1(G52), .A2(n638), .ZN(n525) );
  NAND2_X1 U572 ( .A1(n526), .A2(n525), .ZN(n533) );
  NOR2_X1 U573 ( .A1(n618), .A2(n527), .ZN(n646) );
  NAND2_X1 U574 ( .A1(n646), .A2(G77), .ZN(n528) );
  XOR2_X1 U575 ( .A(KEYINPUT69), .B(n528), .Z(n530) );
  NOR2_X1 U576 ( .A1(G651), .A2(G543), .ZN(n642) );
  NAND2_X1 U577 ( .A1(n642), .A2(G90), .ZN(n529) );
  NAND2_X1 U578 ( .A1(n530), .A2(n529), .ZN(n531) );
  XOR2_X1 U579 ( .A(KEYINPUT9), .B(n531), .Z(n532) );
  NOR2_X1 U580 ( .A1(n533), .A2(n532), .ZN(G171) );
  INV_X1 U581 ( .A(G57), .ZN(G237) );
  NAND2_X1 U582 ( .A1(G126), .A2(n891), .ZN(n535) );
  NAND2_X1 U583 ( .A1(G114), .A2(n890), .ZN(n534) );
  NAND2_X1 U584 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U585 ( .A(n536), .B(KEYINPUT92), .ZN(n541) );
  BUF_X1 U586 ( .A(n537), .Z(n885) );
  NAND2_X1 U587 ( .A1(n885), .A2(G102), .ZN(n539) );
  NAND2_X1 U588 ( .A1(G138), .A2(n543), .ZN(n538) );
  NAND2_X1 U589 ( .A1(n539), .A2(n538), .ZN(n540) );
  NOR2_X1 U590 ( .A1(n541), .A2(n540), .ZN(n542) );
  XOR2_X1 U591 ( .A(n542), .B(KEYINPUT93), .Z(G164) );
  AND2_X1 U592 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U593 ( .A1(G111), .A2(n890), .ZN(n546) );
  INV_X1 U594 ( .A(n543), .ZN(n544) );
  INV_X1 U595 ( .A(n544), .ZN(n887) );
  NAND2_X1 U596 ( .A1(G135), .A2(n887), .ZN(n545) );
  NAND2_X1 U597 ( .A1(n546), .A2(n545), .ZN(n549) );
  NAND2_X1 U598 ( .A1(n891), .A2(G123), .ZN(n547) );
  XOR2_X1 U599 ( .A(KEYINPUT18), .B(n547), .Z(n548) );
  NOR2_X1 U600 ( .A1(n549), .A2(n548), .ZN(n551) );
  NAND2_X1 U601 ( .A1(n885), .A2(G99), .ZN(n550) );
  NAND2_X1 U602 ( .A1(n551), .A2(n550), .ZN(n990) );
  XNOR2_X1 U603 ( .A(G2096), .B(n990), .ZN(n552) );
  OR2_X1 U604 ( .A1(G2100), .A2(n552), .ZN(G156) );
  INV_X1 U605 ( .A(G108), .ZN(G238) );
  INV_X1 U606 ( .A(G120), .ZN(G236) );
  INV_X1 U607 ( .A(G132), .ZN(G219) );
  NAND2_X1 U608 ( .A1(G7), .A2(G661), .ZN(n553) );
  XNOR2_X1 U609 ( .A(n553), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U610 ( .A(KEYINPUT11), .B(KEYINPUT74), .Z(n555) );
  XNOR2_X1 U611 ( .A(G223), .B(KEYINPUT73), .ZN(n827) );
  NAND2_X1 U612 ( .A1(G567), .A2(n827), .ZN(n554) );
  XNOR2_X1 U613 ( .A(n555), .B(n554), .ZN(G234) );
  XNOR2_X1 U614 ( .A(KEYINPUT13), .B(KEYINPUT75), .ZN(n560) );
  NAND2_X1 U615 ( .A1(n642), .A2(G81), .ZN(n556) );
  XNOR2_X1 U616 ( .A(n556), .B(KEYINPUT12), .ZN(n558) );
  NAND2_X1 U617 ( .A1(G68), .A2(n646), .ZN(n557) );
  NAND2_X1 U618 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U619 ( .A(n560), .B(n559), .ZN(n563) );
  NAND2_X1 U620 ( .A1(n637), .A2(G56), .ZN(n561) );
  XOR2_X1 U621 ( .A(KEYINPUT14), .B(n561), .Z(n562) );
  NOR2_X1 U622 ( .A1(n563), .A2(n562), .ZN(n565) );
  NAND2_X1 U623 ( .A1(n638), .A2(G43), .ZN(n564) );
  NAND2_X1 U624 ( .A1(n565), .A2(n564), .ZN(n910) );
  INV_X1 U625 ( .A(G860), .ZN(n597) );
  OR2_X1 U626 ( .A1(n910), .A2(n597), .ZN(G153) );
  XOR2_X1 U627 ( .A(KEYINPUT76), .B(G171), .Z(G301) );
  NAND2_X1 U628 ( .A1(G868), .A2(G301), .ZN(n575) );
  NAND2_X1 U629 ( .A1(G66), .A2(n637), .ZN(n567) );
  NAND2_X1 U630 ( .A1(G92), .A2(n642), .ZN(n566) );
  NAND2_X1 U631 ( .A1(n567), .A2(n566), .ZN(n572) );
  NAND2_X1 U632 ( .A1(G54), .A2(n638), .ZN(n569) );
  NAND2_X1 U633 ( .A1(G79), .A2(n646), .ZN(n568) );
  NAND2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U635 ( .A(KEYINPUT77), .B(n570), .Z(n571) );
  NOR2_X1 U636 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U637 ( .A(KEYINPUT15), .B(n573), .ZN(n911) );
  INV_X1 U638 ( .A(G868), .ZN(n659) );
  NAND2_X1 U639 ( .A1(n911), .A2(n659), .ZN(n574) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(G284) );
  NAND2_X1 U641 ( .A1(G63), .A2(n637), .ZN(n577) );
  NAND2_X1 U642 ( .A1(G51), .A2(n638), .ZN(n576) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(KEYINPUT6), .B(n578), .ZN(n585) );
  NAND2_X1 U645 ( .A1(n642), .A2(G89), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n579), .B(KEYINPUT4), .ZN(n581) );
  NAND2_X1 U647 ( .A1(G76), .A2(n646), .ZN(n580) );
  NAND2_X1 U648 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U649 ( .A(KEYINPUT78), .B(n582), .Z(n583) );
  XNOR2_X1 U650 ( .A(KEYINPUT5), .B(n583), .ZN(n584) );
  NOR2_X1 U651 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U652 ( .A(KEYINPUT7), .B(n586), .Z(G168) );
  XOR2_X1 U653 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U654 ( .A1(n646), .A2(G78), .ZN(n587) );
  XNOR2_X1 U655 ( .A(n587), .B(KEYINPUT70), .ZN(n589) );
  NAND2_X1 U656 ( .A1(G91), .A2(n642), .ZN(n588) );
  NAND2_X1 U657 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U658 ( .A(KEYINPUT71), .B(n590), .ZN(n594) );
  NAND2_X1 U659 ( .A1(G65), .A2(n637), .ZN(n592) );
  NAND2_X1 U660 ( .A1(G53), .A2(n638), .ZN(n591) );
  AND2_X1 U661 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U662 ( .A1(n594), .A2(n593), .ZN(G299) );
  NOR2_X1 U663 ( .A1(G286), .A2(n659), .ZN(n596) );
  NOR2_X1 U664 ( .A1(G868), .A2(G299), .ZN(n595) );
  NOR2_X1 U665 ( .A1(n596), .A2(n595), .ZN(G297) );
  NAND2_X1 U666 ( .A1(n597), .A2(G559), .ZN(n598) );
  INV_X1 U667 ( .A(n911), .ZN(n611) );
  NAND2_X1 U668 ( .A1(n598), .A2(n611), .ZN(n599) );
  XNOR2_X1 U669 ( .A(n599), .B(KEYINPUT16), .ZN(n600) );
  XOR2_X1 U670 ( .A(KEYINPUT79), .B(n600), .Z(G148) );
  NOR2_X1 U671 ( .A1(n911), .A2(n659), .ZN(n601) );
  XOR2_X1 U672 ( .A(KEYINPUT80), .B(n601), .Z(n602) );
  NOR2_X1 U673 ( .A1(G559), .A2(n602), .ZN(n604) );
  NOR2_X1 U674 ( .A1(G868), .A2(n910), .ZN(n603) );
  NOR2_X1 U675 ( .A1(n604), .A2(n603), .ZN(G282) );
  NAND2_X1 U676 ( .A1(G67), .A2(n637), .ZN(n606) );
  NAND2_X1 U677 ( .A1(G55), .A2(n638), .ZN(n605) );
  NAND2_X1 U678 ( .A1(n606), .A2(n605), .ZN(n610) );
  NAND2_X1 U679 ( .A1(G93), .A2(n642), .ZN(n608) );
  NAND2_X1 U680 ( .A1(G80), .A2(n646), .ZN(n607) );
  NAND2_X1 U681 ( .A1(n608), .A2(n607), .ZN(n609) );
  NOR2_X1 U682 ( .A1(n610), .A2(n609), .ZN(n660) );
  NAND2_X1 U683 ( .A1(n611), .A2(G559), .ZN(n657) );
  XNOR2_X1 U684 ( .A(n910), .B(n657), .ZN(n612) );
  NOR2_X1 U685 ( .A1(G860), .A2(n612), .ZN(n613) );
  XOR2_X1 U686 ( .A(KEYINPUT81), .B(n613), .Z(n614) );
  XNOR2_X1 U687 ( .A(n660), .B(n614), .ZN(G145) );
  NAND2_X1 U688 ( .A1(G49), .A2(n638), .ZN(n616) );
  NAND2_X1 U689 ( .A1(G74), .A2(G651), .ZN(n615) );
  NAND2_X1 U690 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U691 ( .A1(n637), .A2(n617), .ZN(n620) );
  NAND2_X1 U692 ( .A1(n618), .A2(G87), .ZN(n619) );
  NAND2_X1 U693 ( .A1(n620), .A2(n619), .ZN(G288) );
  NAND2_X1 U694 ( .A1(G88), .A2(n642), .ZN(n622) );
  NAND2_X1 U695 ( .A1(G75), .A2(n646), .ZN(n621) );
  NAND2_X1 U696 ( .A1(n622), .A2(n621), .ZN(n626) );
  NAND2_X1 U697 ( .A1(G62), .A2(n637), .ZN(n624) );
  NAND2_X1 U698 ( .A1(G50), .A2(n638), .ZN(n623) );
  NAND2_X1 U699 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U700 ( .A1(n626), .A2(n625), .ZN(G166) );
  NAND2_X1 U701 ( .A1(G61), .A2(n637), .ZN(n628) );
  NAND2_X1 U702 ( .A1(G86), .A2(n642), .ZN(n627) );
  NAND2_X1 U703 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U704 ( .A(KEYINPUT82), .B(n629), .ZN(n635) );
  NAND2_X1 U705 ( .A1(G73), .A2(n646), .ZN(n630) );
  XOR2_X1 U706 ( .A(KEYINPUT2), .B(n630), .Z(n631) );
  XNOR2_X1 U707 ( .A(n631), .B(KEYINPUT83), .ZN(n633) );
  NAND2_X1 U708 ( .A1(G48), .A2(n638), .ZN(n632) );
  NAND2_X1 U709 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U710 ( .A1(n635), .A2(n634), .ZN(n636) );
  XOR2_X1 U711 ( .A(KEYINPUT84), .B(n636), .Z(G305) );
  NAND2_X1 U712 ( .A1(G60), .A2(n637), .ZN(n640) );
  NAND2_X1 U713 ( .A1(G47), .A2(n638), .ZN(n639) );
  NAND2_X1 U714 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U715 ( .A(KEYINPUT68), .B(n641), .ZN(n645) );
  NAND2_X1 U716 ( .A1(G85), .A2(n642), .ZN(n643) );
  XNOR2_X1 U717 ( .A(KEYINPUT67), .B(n643), .ZN(n644) );
  NOR2_X1 U718 ( .A1(n645), .A2(n644), .ZN(n648) );
  NAND2_X1 U719 ( .A1(n646), .A2(G72), .ZN(n647) );
  NAND2_X1 U720 ( .A1(n648), .A2(n647), .ZN(G290) );
  INV_X1 U721 ( .A(G299), .ZN(n916) );
  XNOR2_X1 U722 ( .A(KEYINPUT19), .B(KEYINPUT85), .ZN(n650) );
  XNOR2_X1 U723 ( .A(G288), .B(KEYINPUT86), .ZN(n649) );
  XNOR2_X1 U724 ( .A(n650), .B(n649), .ZN(n651) );
  XOR2_X1 U725 ( .A(n651), .B(n660), .Z(n653) );
  XNOR2_X1 U726 ( .A(G166), .B(G305), .ZN(n652) );
  XNOR2_X1 U727 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U728 ( .A(n654), .B(G290), .ZN(n655) );
  XNOR2_X1 U729 ( .A(n655), .B(n910), .ZN(n656) );
  XNOR2_X1 U730 ( .A(n916), .B(n656), .ZN(n836) );
  XOR2_X1 U731 ( .A(n836), .B(n657), .Z(n658) );
  NOR2_X1 U732 ( .A1(n659), .A2(n658), .ZN(n662) );
  NOR2_X1 U733 ( .A1(G868), .A2(n660), .ZN(n661) );
  NOR2_X1 U734 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U735 ( .A(KEYINPUT87), .B(n663), .ZN(G295) );
  XOR2_X1 U736 ( .A(KEYINPUT20), .B(KEYINPUT88), .Z(n665) );
  NAND2_X1 U737 ( .A1(G2084), .A2(G2078), .ZN(n664) );
  XNOR2_X1 U738 ( .A(n665), .B(n664), .ZN(n666) );
  NAND2_X1 U739 ( .A1(n666), .A2(G2090), .ZN(n667) );
  XOR2_X1 U740 ( .A(KEYINPUT89), .B(n667), .Z(n668) );
  XNOR2_X1 U741 ( .A(KEYINPUT21), .B(n668), .ZN(n669) );
  NAND2_X1 U742 ( .A1(n669), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U743 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U744 ( .A(KEYINPUT72), .B(G82), .Z(G220) );
  NOR2_X1 U745 ( .A1(G220), .A2(G219), .ZN(n670) );
  XNOR2_X1 U746 ( .A(KEYINPUT22), .B(n670), .ZN(n671) );
  NAND2_X1 U747 ( .A1(n671), .A2(G96), .ZN(n672) );
  NOR2_X1 U748 ( .A1(G218), .A2(n672), .ZN(n673) );
  XOR2_X1 U749 ( .A(KEYINPUT90), .B(n673), .Z(n834) );
  NAND2_X1 U750 ( .A1(n834), .A2(G2106), .ZN(n674) );
  XNOR2_X1 U751 ( .A(n674), .B(KEYINPUT91), .ZN(n678) );
  NOR2_X1 U752 ( .A1(G236), .A2(G238), .ZN(n675) );
  NAND2_X1 U753 ( .A1(G69), .A2(n675), .ZN(n676) );
  OR2_X1 U754 ( .A1(G237), .A2(n676), .ZN(n833) );
  AND2_X1 U755 ( .A1(G567), .A2(n833), .ZN(n677) );
  NOR2_X1 U756 ( .A1(n678), .A2(n677), .ZN(G319) );
  INV_X1 U757 ( .A(G319), .ZN(n907) );
  NAND2_X1 U758 ( .A1(G483), .A2(G661), .ZN(n679) );
  NOR2_X1 U759 ( .A1(n907), .A2(n679), .ZN(n830) );
  NAND2_X1 U760 ( .A1(n830), .A2(G36), .ZN(G176) );
  XOR2_X1 U761 ( .A(KEYINPUT94), .B(G166), .Z(G303) );
  NAND2_X1 U762 ( .A1(G105), .A2(n885), .ZN(n680) );
  XNOR2_X1 U763 ( .A(n680), .B(KEYINPUT38), .ZN(n687) );
  NAND2_X1 U764 ( .A1(G117), .A2(n890), .ZN(n682) );
  NAND2_X1 U765 ( .A1(G129), .A2(n891), .ZN(n681) );
  NAND2_X1 U766 ( .A1(n682), .A2(n681), .ZN(n685) );
  NAND2_X1 U767 ( .A1(n887), .A2(G141), .ZN(n683) );
  XOR2_X1 U768 ( .A(KEYINPUT96), .B(n683), .Z(n684) );
  NOR2_X1 U769 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U770 ( .A1(n687), .A2(n686), .ZN(n875) );
  NAND2_X1 U771 ( .A1(G1996), .A2(n875), .ZN(n688) );
  XNOR2_X1 U772 ( .A(n688), .B(KEYINPUT97), .ZN(n696) );
  XOR2_X1 U773 ( .A(KEYINPUT95), .B(G1991), .Z(n963) );
  NAND2_X1 U774 ( .A1(n885), .A2(G95), .ZN(n690) );
  NAND2_X1 U775 ( .A1(G131), .A2(n887), .ZN(n689) );
  NAND2_X1 U776 ( .A1(n690), .A2(n689), .ZN(n694) );
  NAND2_X1 U777 ( .A1(G107), .A2(n890), .ZN(n692) );
  NAND2_X1 U778 ( .A1(G119), .A2(n891), .ZN(n691) );
  NAND2_X1 U779 ( .A1(n692), .A2(n691), .ZN(n693) );
  OR2_X1 U780 ( .A1(n694), .A2(n693), .ZN(n870) );
  AND2_X1 U781 ( .A1(n963), .A2(n870), .ZN(n695) );
  NOR2_X1 U782 ( .A1(n696), .A2(n695), .ZN(n1000) );
  XOR2_X1 U783 ( .A(G1986), .B(G290), .Z(n917) );
  NAND2_X1 U784 ( .A1(n1000), .A2(n917), .ZN(n698) );
  NOR2_X1 U785 ( .A1(G164), .A2(G1384), .ZN(n701) );
  NAND2_X1 U786 ( .A1(G160), .A2(G40), .ZN(n699) );
  NOR2_X1 U787 ( .A1(n701), .A2(n699), .ZN(n813) );
  NAND2_X1 U788 ( .A1(n698), .A2(n813), .ZN(n803) );
  XOR2_X1 U789 ( .A(KEYINPUT98), .B(n699), .Z(n700) );
  AND2_X1 U790 ( .A1(n701), .A2(n700), .ZN(n733) );
  INV_X1 U791 ( .A(n733), .ZN(n740) );
  NAND2_X1 U792 ( .A1(G8), .A2(n740), .ZN(n785) );
  NOR2_X1 U793 ( .A1(G1971), .A2(n785), .ZN(n703) );
  NOR2_X1 U794 ( .A1(G2090), .A2(n740), .ZN(n702) );
  NOR2_X1 U795 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U796 ( .A1(n704), .A2(G303), .ZN(n750) );
  NAND2_X1 U797 ( .A1(n733), .A2(G2072), .ZN(n705) );
  XOR2_X1 U798 ( .A(KEYINPUT27), .B(n705), .Z(n707) );
  NAND2_X1 U799 ( .A1(G1956), .A2(n740), .ZN(n706) );
  NAND2_X1 U800 ( .A1(n707), .A2(n706), .ZN(n709) );
  XNOR2_X1 U801 ( .A(n709), .B(n708), .ZN(n712) );
  NOR2_X1 U802 ( .A1(n916), .A2(n712), .ZN(n711) );
  XNOR2_X1 U803 ( .A(n711), .B(n710), .ZN(n731) );
  NAND2_X1 U804 ( .A1(n916), .A2(n712), .ZN(n729) );
  XNOR2_X1 U805 ( .A(KEYINPUT64), .B(KEYINPUT26), .ZN(n719) );
  NOR2_X1 U806 ( .A1(G1996), .A2(n719), .ZN(n713) );
  NOR2_X1 U807 ( .A1(n910), .A2(n713), .ZN(n717) );
  NAND2_X1 U808 ( .A1(G1348), .A2(n740), .ZN(n715) );
  NAND2_X1 U809 ( .A1(G2067), .A2(n733), .ZN(n714) );
  NAND2_X1 U810 ( .A1(n715), .A2(n714), .ZN(n725) );
  NAND2_X1 U811 ( .A1(n911), .A2(n725), .ZN(n716) );
  NAND2_X1 U812 ( .A1(n717), .A2(n716), .ZN(n724) );
  INV_X1 U813 ( .A(G1341), .ZN(n938) );
  NAND2_X1 U814 ( .A1(n938), .A2(n719), .ZN(n718) );
  NAND2_X1 U815 ( .A1(n718), .A2(n740), .ZN(n722) );
  INV_X1 U816 ( .A(G1996), .ZN(n971) );
  NOR2_X1 U817 ( .A1(n971), .A2(n740), .ZN(n720) );
  NAND2_X1 U818 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U819 ( .A1(n722), .A2(n721), .ZN(n723) );
  NOR2_X1 U820 ( .A1(n724), .A2(n723), .ZN(n727) );
  NOR2_X1 U821 ( .A1(n725), .A2(n911), .ZN(n726) );
  NOR2_X1 U822 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U823 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U824 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U825 ( .A(n732), .B(KEYINPUT29), .ZN(n737) );
  XNOR2_X1 U826 ( .A(KEYINPUT25), .B(G2078), .ZN(n970) );
  NOR2_X1 U827 ( .A1(n740), .A2(n970), .ZN(n735) );
  INV_X1 U828 ( .A(G1961), .ZN(n937) );
  NOR2_X1 U829 ( .A1(n733), .A2(n937), .ZN(n734) );
  NOR2_X1 U830 ( .A1(n735), .A2(n734), .ZN(n739) );
  AND2_X1 U831 ( .A1(G171), .A2(n739), .ZN(n736) );
  NOR2_X1 U832 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U833 ( .A(n738), .B(KEYINPUT101), .ZN(n754) );
  NOR2_X1 U834 ( .A1(G171), .A2(n739), .ZN(n745) );
  NOR2_X1 U835 ( .A1(G1966), .A2(n785), .ZN(n756) );
  NOR2_X1 U836 ( .A1(G2084), .A2(n740), .ZN(n755) );
  NOR2_X1 U837 ( .A1(n756), .A2(n755), .ZN(n741) );
  NAND2_X1 U838 ( .A1(G8), .A2(n741), .ZN(n742) );
  XNOR2_X1 U839 ( .A(KEYINPUT30), .B(n742), .ZN(n743) );
  NOR2_X1 U840 ( .A1(G168), .A2(n743), .ZN(n744) );
  NOR2_X1 U841 ( .A1(n745), .A2(n744), .ZN(n746) );
  XOR2_X1 U842 ( .A(KEYINPUT31), .B(n746), .Z(n753) );
  NAND2_X1 U843 ( .A1(n754), .A2(n753), .ZN(n747) );
  NAND2_X1 U844 ( .A1(n747), .A2(G286), .ZN(n748) );
  XOR2_X1 U845 ( .A(KEYINPUT103), .B(n748), .Z(n749) );
  NAND2_X1 U846 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U847 ( .A1(n751), .A2(G8), .ZN(n752) );
  XNOR2_X1 U848 ( .A(n752), .B(KEYINPUT32), .ZN(n776) );
  AND2_X1 U849 ( .A1(n754), .A2(n753), .ZN(n759) );
  AND2_X1 U850 ( .A1(G8), .A2(n755), .ZN(n757) );
  OR2_X1 U851 ( .A1(n757), .A2(n756), .ZN(n758) );
  OR2_X1 U852 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U853 ( .A(KEYINPUT102), .B(n760), .ZN(n775) );
  NAND2_X1 U854 ( .A1(G1976), .A2(G288), .ZN(n915) );
  AND2_X1 U855 ( .A1(n775), .A2(n915), .ZN(n761) );
  NAND2_X1 U856 ( .A1(n776), .A2(n761), .ZN(n768) );
  INV_X1 U857 ( .A(n915), .ZN(n763) );
  NOR2_X1 U858 ( .A1(G1976), .A2(G288), .ZN(n769) );
  NOR2_X1 U859 ( .A1(G303), .A2(G1971), .ZN(n762) );
  NOR2_X1 U860 ( .A1(n769), .A2(n762), .ZN(n921) );
  OR2_X1 U861 ( .A1(n763), .A2(n921), .ZN(n764) );
  OR2_X1 U862 ( .A1(n785), .A2(n764), .ZN(n766) );
  INV_X1 U863 ( .A(KEYINPUT33), .ZN(n765) );
  AND2_X1 U864 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U865 ( .A1(n768), .A2(n767), .ZN(n774) );
  NAND2_X1 U866 ( .A1(n769), .A2(KEYINPUT33), .ZN(n770) );
  NOR2_X1 U867 ( .A1(n770), .A2(n785), .ZN(n772) );
  XOR2_X1 U868 ( .A(G1981), .B(G305), .Z(n928) );
  INV_X1 U869 ( .A(n928), .ZN(n771) );
  NOR2_X1 U870 ( .A1(n772), .A2(n771), .ZN(n773) );
  AND2_X1 U871 ( .A1(n774), .A2(n773), .ZN(n790) );
  NAND2_X1 U872 ( .A1(n776), .A2(n775), .ZN(n784) );
  NOR2_X1 U873 ( .A1(G2090), .A2(G303), .ZN(n777) );
  NAND2_X1 U874 ( .A1(G8), .A2(n777), .ZN(n782) );
  NOR2_X1 U875 ( .A1(G1981), .A2(G305), .ZN(n778) );
  XNOR2_X1 U876 ( .A(n778), .B(KEYINPUT99), .ZN(n779) );
  XNOR2_X1 U877 ( .A(n779), .B(KEYINPUT24), .ZN(n780) );
  NOR2_X1 U878 ( .A1(n785), .A2(n780), .ZN(n786) );
  INV_X1 U879 ( .A(n786), .ZN(n781) );
  AND2_X1 U880 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U881 ( .A1(n784), .A2(n783), .ZN(n788) );
  OR2_X1 U882 ( .A1(n786), .A2(n785), .ZN(n787) );
  AND2_X1 U883 ( .A1(n788), .A2(n787), .ZN(n789) );
  NOR2_X1 U884 ( .A1(n790), .A2(n789), .ZN(n801) );
  XNOR2_X1 U885 ( .A(G2067), .B(KEYINPUT37), .ZN(n811) );
  NAND2_X1 U886 ( .A1(n885), .A2(G104), .ZN(n792) );
  NAND2_X1 U887 ( .A1(G140), .A2(n887), .ZN(n791) );
  NAND2_X1 U888 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U889 ( .A(KEYINPUT34), .B(n793), .ZN(n798) );
  NAND2_X1 U890 ( .A1(G116), .A2(n890), .ZN(n795) );
  NAND2_X1 U891 ( .A1(G128), .A2(n891), .ZN(n794) );
  NAND2_X1 U892 ( .A1(n795), .A2(n794), .ZN(n796) );
  XOR2_X1 U893 ( .A(KEYINPUT35), .B(n796), .Z(n797) );
  NOR2_X1 U894 ( .A1(n798), .A2(n797), .ZN(n799) );
  XNOR2_X1 U895 ( .A(KEYINPUT36), .B(n799), .ZN(n900) );
  NOR2_X1 U896 ( .A1(n811), .A2(n900), .ZN(n1002) );
  NAND2_X1 U897 ( .A1(n813), .A2(n1002), .ZN(n809) );
  INV_X1 U898 ( .A(n809), .ZN(n800) );
  NOR2_X1 U899 ( .A1(n801), .A2(n800), .ZN(n802) );
  NAND2_X1 U900 ( .A1(n803), .A2(n802), .ZN(n816) );
  NOR2_X1 U901 ( .A1(G1996), .A2(n875), .ZN(n993) );
  INV_X1 U902 ( .A(n1000), .ZN(n806) );
  NOR2_X1 U903 ( .A1(G1986), .A2(G290), .ZN(n804) );
  NOR2_X1 U904 ( .A1(n963), .A2(n870), .ZN(n989) );
  NOR2_X1 U905 ( .A1(n804), .A2(n989), .ZN(n805) );
  NOR2_X1 U906 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U907 ( .A1(n993), .A2(n807), .ZN(n808) );
  XNOR2_X1 U908 ( .A(n808), .B(KEYINPUT39), .ZN(n810) );
  NAND2_X1 U909 ( .A1(n810), .A2(n809), .ZN(n812) );
  NAND2_X1 U910 ( .A1(n811), .A2(n900), .ZN(n1010) );
  NAND2_X1 U911 ( .A1(n812), .A2(n1010), .ZN(n814) );
  NAND2_X1 U912 ( .A1(n814), .A2(n813), .ZN(n815) );
  NAND2_X1 U913 ( .A1(n816), .A2(n815), .ZN(n817) );
  XNOR2_X1 U914 ( .A(n817), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U915 ( .A(G1348), .B(G2454), .ZN(n818) );
  XNOR2_X1 U916 ( .A(n818), .B(G2430), .ZN(n819) );
  XNOR2_X1 U917 ( .A(n819), .B(G1341), .ZN(n825) );
  XOR2_X1 U918 ( .A(G2443), .B(G2427), .Z(n821) );
  XNOR2_X1 U919 ( .A(G2438), .B(G2446), .ZN(n820) );
  XNOR2_X1 U920 ( .A(n821), .B(n820), .ZN(n823) );
  XOR2_X1 U921 ( .A(G2451), .B(G2435), .Z(n822) );
  XNOR2_X1 U922 ( .A(n823), .B(n822), .ZN(n824) );
  XNOR2_X1 U923 ( .A(n825), .B(n824), .ZN(n826) );
  NAND2_X1 U924 ( .A1(n826), .A2(G14), .ZN(n905) );
  XOR2_X1 U925 ( .A(KEYINPUT104), .B(n905), .Z(G401) );
  NAND2_X1 U926 ( .A1(n827), .A2(G2106), .ZN(n828) );
  XOR2_X1 U927 ( .A(KEYINPUT105), .B(n828), .Z(G217) );
  AND2_X1 U928 ( .A1(G15), .A2(G2), .ZN(n829) );
  NAND2_X1 U929 ( .A1(G661), .A2(n829), .ZN(G259) );
  NAND2_X1 U930 ( .A1(G1), .A2(G3), .ZN(n831) );
  NAND2_X1 U931 ( .A1(n831), .A2(n830), .ZN(n832) );
  XNOR2_X1 U932 ( .A(n832), .B(KEYINPUT106), .ZN(G188) );
  XNOR2_X1 U933 ( .A(G96), .B(KEYINPUT107), .ZN(G221) );
  NOR2_X1 U935 ( .A1(n834), .A2(n833), .ZN(n835) );
  XNOR2_X1 U936 ( .A(KEYINPUT108), .B(n835), .ZN(G325) );
  INV_X1 U937 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U938 ( .A(G286), .B(n911), .ZN(n837) );
  XNOR2_X1 U939 ( .A(n837), .B(n836), .ZN(n838) );
  XNOR2_X1 U940 ( .A(n838), .B(G171), .ZN(n839) );
  NOR2_X1 U941 ( .A1(G37), .A2(n839), .ZN(G397) );
  XOR2_X1 U942 ( .A(G1956), .B(G1961), .Z(n841) );
  XNOR2_X1 U943 ( .A(G1986), .B(G1966), .ZN(n840) );
  XNOR2_X1 U944 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U945 ( .A(n842), .B(G2474), .Z(n844) );
  XNOR2_X1 U946 ( .A(G1971), .B(G1976), .ZN(n843) );
  XNOR2_X1 U947 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U948 ( .A(KEYINPUT41), .B(G1981), .Z(n846) );
  XNOR2_X1 U949 ( .A(G1996), .B(G1991), .ZN(n845) );
  XNOR2_X1 U950 ( .A(n846), .B(n845), .ZN(n847) );
  XNOR2_X1 U951 ( .A(n848), .B(n847), .ZN(G229) );
  XOR2_X1 U952 ( .A(KEYINPUT109), .B(G2084), .Z(n850) );
  XNOR2_X1 U953 ( .A(G2067), .B(G2072), .ZN(n849) );
  XNOR2_X1 U954 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U955 ( .A(n851), .B(G2100), .Z(n853) );
  XNOR2_X1 U956 ( .A(G2078), .B(G2090), .ZN(n852) );
  XNOR2_X1 U957 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U958 ( .A(G2096), .B(G2678), .Z(n855) );
  XNOR2_X1 U959 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n854) );
  XNOR2_X1 U960 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U961 ( .A(n857), .B(n856), .Z(G227) );
  NAND2_X1 U962 ( .A1(n891), .A2(G124), .ZN(n858) );
  XNOR2_X1 U963 ( .A(n858), .B(KEYINPUT44), .ZN(n860) );
  NAND2_X1 U964 ( .A1(G136), .A2(n887), .ZN(n859) );
  NAND2_X1 U965 ( .A1(n860), .A2(n859), .ZN(n861) );
  XNOR2_X1 U966 ( .A(KEYINPUT110), .B(n861), .ZN(n865) );
  NAND2_X1 U967 ( .A1(G112), .A2(n890), .ZN(n863) );
  NAND2_X1 U968 ( .A1(G100), .A2(n885), .ZN(n862) );
  NAND2_X1 U969 ( .A1(n863), .A2(n862), .ZN(n864) );
  NOR2_X1 U970 ( .A1(n865), .A2(n864), .ZN(n866) );
  XOR2_X1 U971 ( .A(KEYINPUT111), .B(n866), .Z(G162) );
  XOR2_X1 U972 ( .A(KEYINPUT114), .B(KEYINPUT46), .Z(n868) );
  XNOR2_X1 U973 ( .A(KEYINPUT48), .B(KEYINPUT115), .ZN(n867) );
  XNOR2_X1 U974 ( .A(n868), .B(n867), .ZN(n869) );
  XNOR2_X1 U975 ( .A(n990), .B(n869), .ZN(n872) );
  XOR2_X1 U976 ( .A(G160), .B(n870), .Z(n871) );
  XNOR2_X1 U977 ( .A(n872), .B(n871), .ZN(n873) );
  XOR2_X1 U978 ( .A(G164), .B(n873), .Z(n874) );
  XNOR2_X1 U979 ( .A(n875), .B(n874), .ZN(n884) );
  NAND2_X1 U980 ( .A1(G118), .A2(n890), .ZN(n877) );
  NAND2_X1 U981 ( .A1(G130), .A2(n891), .ZN(n876) );
  NAND2_X1 U982 ( .A1(n877), .A2(n876), .ZN(n882) );
  NAND2_X1 U983 ( .A1(n885), .A2(G106), .ZN(n879) );
  NAND2_X1 U984 ( .A1(G142), .A2(n887), .ZN(n878) );
  NAND2_X1 U985 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U986 ( .A(KEYINPUT45), .B(n880), .Z(n881) );
  NOR2_X1 U987 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U988 ( .A(n884), .B(n883), .Z(n899) );
  NAND2_X1 U989 ( .A1(n885), .A2(G103), .ZN(n886) );
  XNOR2_X1 U990 ( .A(n886), .B(KEYINPUT112), .ZN(n889) );
  NAND2_X1 U991 ( .A1(G139), .A2(n887), .ZN(n888) );
  NAND2_X1 U992 ( .A1(n889), .A2(n888), .ZN(n896) );
  NAND2_X1 U993 ( .A1(G115), .A2(n890), .ZN(n893) );
  NAND2_X1 U994 ( .A1(G127), .A2(n891), .ZN(n892) );
  NAND2_X1 U995 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U996 ( .A(KEYINPUT47), .B(n894), .Z(n895) );
  NOR2_X1 U997 ( .A1(n896), .A2(n895), .ZN(n897) );
  XOR2_X1 U998 ( .A(KEYINPUT113), .B(n897), .Z(n1004) );
  XNOR2_X1 U999 ( .A(n1004), .B(G162), .ZN(n898) );
  XNOR2_X1 U1000 ( .A(n899), .B(n898), .ZN(n901) );
  XNOR2_X1 U1001 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n902), .ZN(G395) );
  NOR2_X1 U1003 ( .A1(G229), .A2(G227), .ZN(n903) );
  XOR2_X1 U1004 ( .A(KEYINPUT49), .B(n903), .Z(n904) );
  NAND2_X1 U1005 ( .A1(n905), .A2(n904), .ZN(n906) );
  NOR2_X1 U1006 ( .A1(G397), .A2(n906), .ZN(n909) );
  NOR2_X1 U1007 ( .A1(G395), .A2(n907), .ZN(n908) );
  NAND2_X1 U1008 ( .A1(n909), .A2(n908), .ZN(G225) );
  INV_X1 U1009 ( .A(G225), .ZN(G308) );
  INV_X1 U1010 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U1011 ( .A(G171), .B(G1961), .ZN(n927) );
  XNOR2_X1 U1012 ( .A(n938), .B(n910), .ZN(n913) );
  XOR2_X1 U1013 ( .A(G1348), .B(n911), .Z(n912) );
  NAND2_X1 U1014 ( .A1(n913), .A2(n912), .ZN(n925) );
  NAND2_X1 U1015 ( .A1(G303), .A2(G1971), .ZN(n914) );
  NAND2_X1 U1016 ( .A1(n915), .A2(n914), .ZN(n920) );
  XNOR2_X1 U1017 ( .A(n916), .B(G1956), .ZN(n918) );
  NAND2_X1 U1018 ( .A1(n918), .A2(n917), .ZN(n919) );
  NOR2_X1 U1019 ( .A1(n920), .A2(n919), .ZN(n922) );
  NAND2_X1 U1020 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1021 ( .A(KEYINPUT126), .B(n923), .ZN(n924) );
  NOR2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1023 ( .A1(n927), .A2(n926), .ZN(n933) );
  XNOR2_X1 U1024 ( .A(G1966), .B(G168), .ZN(n929) );
  NAND2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1026 ( .A(n930), .B(KEYINPUT125), .ZN(n931) );
  XNOR2_X1 U1027 ( .A(n931), .B(KEYINPUT57), .ZN(n932) );
  NOR2_X1 U1028 ( .A1(n933), .A2(n932), .ZN(n935) );
  XOR2_X1 U1029 ( .A(G16), .B(KEYINPUT56), .Z(n934) );
  NOR2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1031 ( .A(KEYINPUT127), .B(n936), .ZN(n1019) );
  XNOR2_X1 U1032 ( .A(G5), .B(n937), .ZN(n950) );
  XNOR2_X1 U1033 ( .A(G19), .B(n938), .ZN(n942) );
  XNOR2_X1 U1034 ( .A(G1956), .B(G20), .ZN(n940) );
  XNOR2_X1 U1035 ( .A(G1981), .B(G6), .ZN(n939) );
  NOR2_X1 U1036 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1037 ( .A1(n942), .A2(n941), .ZN(n945) );
  XOR2_X1 U1038 ( .A(KEYINPUT59), .B(G1348), .Z(n943) );
  XNOR2_X1 U1039 ( .A(G4), .B(n943), .ZN(n944) );
  NOR2_X1 U1040 ( .A1(n945), .A2(n944), .ZN(n946) );
  XOR2_X1 U1041 ( .A(KEYINPUT60), .B(n946), .Z(n948) );
  XNOR2_X1 U1042 ( .A(G1966), .B(G21), .ZN(n947) );
  NOR2_X1 U1043 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n957) );
  XNOR2_X1 U1045 ( .A(G1971), .B(G22), .ZN(n952) );
  XNOR2_X1 U1046 ( .A(G23), .B(G1976), .ZN(n951) );
  NOR2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n954) );
  XOR2_X1 U1048 ( .A(G1986), .B(G24), .Z(n953) );
  NAND2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1050 ( .A(KEYINPUT58), .B(n955), .ZN(n956) );
  NOR2_X1 U1051 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1052 ( .A(KEYINPUT61), .B(n958), .ZN(n960) );
  INV_X1 U1053 ( .A(G16), .ZN(n959) );
  NAND2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1055 ( .A1(n961), .A2(G11), .ZN(n1017) );
  XOR2_X1 U1056 ( .A(KEYINPUT55), .B(KEYINPUT120), .Z(n987) );
  XOR2_X1 U1057 ( .A(G2090), .B(G35), .Z(n962) );
  XNOR2_X1 U1058 ( .A(KEYINPUT121), .B(n962), .ZN(n979) );
  XOR2_X1 U1059 ( .A(G25), .B(n963), .Z(n969) );
  XOR2_X1 U1060 ( .A(G2067), .B(G26), .Z(n964) );
  NAND2_X1 U1061 ( .A1(n964), .A2(G28), .ZN(n967) );
  XNOR2_X1 U1062 ( .A(G33), .B(G2072), .ZN(n965) );
  XNOR2_X1 U1063 ( .A(KEYINPUT122), .B(n965), .ZN(n966) );
  NOR2_X1 U1064 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1065 ( .A1(n969), .A2(n968), .ZN(n976) );
  XOR2_X1 U1066 ( .A(n970), .B(G27), .Z(n973) );
  XOR2_X1 U1067 ( .A(n971), .B(G32), .Z(n972) );
  NOR2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1069 ( .A(n974), .B(KEYINPUT123), .ZN(n975) );
  NOR2_X1 U1070 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1071 ( .A(n977), .B(KEYINPUT53), .ZN(n978) );
  NOR2_X1 U1072 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1073 ( .A(n980), .B(KEYINPUT124), .ZN(n983) );
  XOR2_X1 U1074 ( .A(G2084), .B(G34), .Z(n981) );
  XNOR2_X1 U1075 ( .A(KEYINPUT54), .B(n981), .ZN(n982) );
  NAND2_X1 U1076 ( .A1(n983), .A2(n982), .ZN(n985) );
  INV_X1 U1077 ( .A(G29), .ZN(n984) );
  NAND2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1079 ( .A(n987), .B(n986), .ZN(n1015) );
  XOR2_X1 U1080 ( .A(KEYINPUT52), .B(KEYINPUT119), .Z(n1013) );
  XOR2_X1 U1081 ( .A(G160), .B(G2084), .Z(n988) );
  NOR2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n991) );
  NAND2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n998) );
  XNOR2_X1 U1084 ( .A(KEYINPUT51), .B(KEYINPUT117), .ZN(n996) );
  XOR2_X1 U1085 ( .A(G2090), .B(G162), .Z(n992) );
  XNOR2_X1 U1086 ( .A(KEYINPUT116), .B(n992), .ZN(n994) );
  NOR2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n995) );
  XOR2_X1 U1088 ( .A(n996), .B(n995), .Z(n997) );
  NOR2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NOR2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XOR2_X1 U1092 ( .A(KEYINPUT118), .B(n1003), .Z(n1009) );
  XOR2_X1 U1093 ( .A(G2072), .B(n1004), .Z(n1006) );
  XOR2_X1 U1094 ( .A(G164), .B(G2078), .Z(n1005) );
  NOR2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XOR2_X1 U1096 ( .A(KEYINPUT50), .B(n1007), .Z(n1008) );
  NOR2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1011) );
  NAND2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1099 ( .A(n1013), .B(n1012), .ZN(n1014) );
  NAND2_X1 U1100 ( .A1(n1015), .A2(n512), .ZN(n1016) );
  NOR2_X1 U1101 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1102 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XOR2_X1 U1103 ( .A(KEYINPUT62), .B(n1020), .Z(G311) );
  INV_X1 U1104 ( .A(G311), .ZN(G150) );
endmodule

