//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 0 1 1 1 0 1 1 0 1 1 1 1 1 1 1 0 0 1 0 0 1 1 0 0 1 0 1 0 1 0 1 1 1 1 0 0 1 0 1 1 0 0 0 1 1 0 1 1 1 0 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:38 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n449, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n564, new_n565, new_n566, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n609, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  INV_X1    g022(.A(G567), .ZN(new_n448));
  NOR2_X1   g023(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT66), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n448), .ZN(new_n457));
  INV_X1    g032(.A(new_n453), .ZN(new_n458));
  AOI21_X1  g033(.A(new_n457), .B1(new_n458), .B2(G2106), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT67), .Z(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n462), .A2(new_n464), .A3(G125), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT68), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n467));
  NAND4_X1  g042(.A1(new_n462), .A2(new_n464), .A3(new_n467), .A4(G125), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n466), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(KEYINPUT69), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n470), .A2(new_n473), .A3(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT72), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT71), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n477), .B1(new_n461), .B2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(G2105), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n479), .A2(KEYINPUT71), .A3(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n476), .B1(new_n481), .B2(G101), .ZN(new_n482));
  INV_X1    g057(.A(G101), .ZN(new_n483));
  AOI211_X1 g058(.A(KEYINPUT72), .B(new_n483), .C1(new_n478), .C2(new_n480), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n463), .B1(new_n461), .B2(KEYINPUT70), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT70), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n487), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n488));
  AOI21_X1  g063(.A(G2105), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n485), .B1(G137), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n475), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G160));
  AOI21_X1  g067(.A(new_n479), .B1(new_n486), .B2(new_n488), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G124), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n479), .A2(G112), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  XNOR2_X1  g072(.A(new_n489), .B(KEYINPUT73), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n497), .B1(new_n498), .B2(G136), .ZN(new_n499));
  XOR2_X1   g074(.A(new_n499), .B(KEYINPUT74), .Z(G162));
  OAI211_X1 g075(.A(new_n479), .B(G138), .C1(KEYINPUT75), .C2(KEYINPUT4), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n501), .B1(KEYINPUT75), .B2(KEYINPUT4), .ZN(new_n502));
  AND2_X1   g077(.A1(new_n462), .A2(new_n464), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G138), .ZN(new_n505));
  AOI211_X1 g080(.A(new_n505), .B(G2105), .C1(new_n486), .C2(new_n488), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT4), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n504), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n479), .A2(G114), .ZN(new_n509));
  OAI21_X1  g084(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n511), .B1(new_n493), .B2(G126), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(G164));
  XNOR2_X1  g089(.A(KEYINPUT5), .B(G543), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(KEYINPUT76), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT76), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n515), .A2(new_n516), .A3(new_n519), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G88), .ZN(new_n522));
  NAND2_X1  g097(.A1(G75), .A2(G543), .ZN(new_n523));
  INV_X1    g098(.A(new_n515), .ZN(new_n524));
  INV_X1    g099(.A(G62), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G543), .ZN(new_n527));
  OR2_X1    g102(.A1(KEYINPUT6), .A2(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(KEYINPUT6), .A2(G651), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n526), .A2(G651), .B1(G50), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n522), .A2(new_n531), .ZN(G303));
  INV_X1    g107(.A(G303), .ZN(G166));
  NAND2_X1  g108(.A1(new_n521), .A2(G89), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n516), .A2(KEYINPUT77), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT77), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n528), .A2(new_n536), .A3(new_n529), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n535), .A2(G543), .A3(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G51), .ZN(new_n540));
  NAND3_X1  g115(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n541), .A2(KEYINPUT7), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(KEYINPUT7), .ZN(new_n543));
  AND2_X1   g118(.A1(G63), .A2(G651), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n542), .A2(new_n543), .B1(new_n515), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n534), .A2(new_n540), .A3(new_n545), .ZN(G286));
  INV_X1    g121(.A(G286), .ZN(G168));
  NAND2_X1  g122(.A1(new_n521), .A2(G90), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n539), .A2(G52), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n550));
  INV_X1    g125(.A(G651), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n548), .A2(new_n549), .A3(new_n552), .ZN(G301));
  INV_X1    g128(.A(G301), .ZN(G171));
  NAND2_X1  g129(.A1(new_n521), .A2(G81), .ZN(new_n555));
  XNOR2_X1  g130(.A(KEYINPUT78), .B(G43), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n539), .A2(new_n556), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n558));
  OR2_X1    g133(.A1(new_n558), .A2(new_n551), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n555), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(G153));
  NAND4_X1  g137(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT79), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND4_X1  g141(.A1(G319), .A2(G483), .A3(G661), .A4(new_n566), .ZN(G188));
  NAND2_X1  g142(.A1(KEYINPUT80), .A2(G53), .ZN(new_n568));
  OR3_X1    g143(.A1(new_n538), .A2(KEYINPUT9), .A3(new_n568), .ZN(new_n569));
  OAI21_X1  g144(.A(KEYINPUT9), .B1(new_n538), .B2(new_n568), .ZN(new_n570));
  NAND2_X1  g145(.A1(G78), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(G65), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n524), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n569), .A2(new_n570), .B1(G651), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n518), .A2(G91), .A3(new_n520), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT81), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n576), .ZN(G299));
  NAND2_X1  g152(.A1(new_n539), .A2(G49), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n579));
  INV_X1    g154(.A(G87), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n518), .A2(new_n520), .ZN(new_n581));
  OAI211_X1 g156(.A(new_n578), .B(new_n579), .C1(new_n580), .C2(new_n581), .ZN(G288));
  NAND2_X1  g157(.A1(new_n515), .A2(G61), .ZN(new_n583));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n585), .A2(G651), .B1(G48), .B2(new_n530), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n518), .A2(G86), .A3(new_n520), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(G305));
  NAND2_X1  g163(.A1(new_n539), .A2(G47), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G85), .ZN(new_n591));
  OAI221_X1 g166(.A(new_n589), .B1(new_n551), .B2(new_n590), .C1(new_n591), .C2(new_n581), .ZN(G290));
  NAND2_X1  g167(.A1(G301), .A2(G868), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n521), .A2(G92), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n594), .B(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(G79), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G66), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n524), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n539), .A2(G54), .B1(G651), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n593), .B1(new_n602), .B2(G868), .ZN(G284));
  OAI21_X1  g178(.A(new_n593), .B1(new_n602), .B2(G868), .ZN(G321));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(G299), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(new_n605), .B2(G168), .ZN(G297));
  OAI21_X1  g182(.A(new_n606), .B1(new_n605), .B2(G168), .ZN(G280));
  XOR2_X1   g183(.A(KEYINPUT82), .B(G559), .Z(new_n609));
  OAI21_X1  g184(.A(new_n602), .B1(G860), .B2(new_n609), .ZN(G148));
  NAND2_X1  g185(.A1(new_n602), .A2(new_n609), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(G868), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(G868), .B2(new_n561), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g189(.A1(new_n503), .A2(new_n481), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT12), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT13), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(G2100), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n493), .A2(G123), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n479), .A2(G111), .ZN(new_n620));
  OAI21_X1  g195(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT73), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n489), .B(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(G135), .ZN(new_n624));
  OAI221_X1 g199(.A(new_n619), .B1(new_n620), .B2(new_n621), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(KEYINPUT83), .B(G2096), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n618), .A2(new_n627), .ZN(G156));
  XOR2_X1   g203(.A(KEYINPUT84), .B(KEYINPUT14), .Z(new_n629));
  XOR2_X1   g204(.A(KEYINPUT15), .B(G2435), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2438), .ZN(new_n631));
  XOR2_X1   g206(.A(G2427), .B(G2430), .Z(new_n632));
  AOI21_X1  g207(.A(new_n629), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(new_n631), .B2(new_n632), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2451), .B(G2454), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT16), .ZN(new_n636));
  XNOR2_X1  g211(.A(G1341), .B(G1348), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n634), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n641), .A2(new_n642), .A3(G14), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT85), .ZN(G401));
  XOR2_X1   g219(.A(G2072), .B(G2078), .Z(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT88), .B(KEYINPUT17), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2067), .B(G2678), .ZN(new_n648));
  INV_X1    g223(.A(KEYINPUT87), .ZN(new_n649));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  INV_X1    g225(.A(new_n648), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n650), .B1(new_n651), .B2(new_n645), .ZN(new_n652));
  AOI22_X1  g227(.A1(new_n647), .A2(new_n648), .B1(new_n649), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n653), .B1(new_n649), .B2(new_n652), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT89), .Z(new_n655));
  INV_X1    g230(.A(new_n650), .ZN(new_n656));
  NOR3_X1   g231(.A1(new_n656), .A2(new_n651), .A3(new_n645), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT86), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT18), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n651), .A2(new_n650), .ZN(new_n660));
  OAI211_X1 g235(.A(new_n655), .B(new_n659), .C1(new_n647), .C2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2096), .B(G2100), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(G227));
  XNOR2_X1  g238(.A(G1971), .B(G1976), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT19), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1956), .B(G2474), .ZN(new_n666));
  INV_X1    g241(.A(KEYINPUT90), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G1961), .B(G1966), .Z(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(KEYINPUT91), .B(KEYINPUT20), .Z(new_n671));
  OR2_X1    g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n668), .A2(new_n669), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n665), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n673), .A2(new_n670), .A3(new_n665), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n671), .B1(new_n670), .B2(new_n665), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT92), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n679), .B(new_n680), .Z(new_n681));
  XOR2_X1   g256(.A(G1991), .B(G1996), .Z(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n679), .B(new_n680), .ZN(new_n684));
  INV_X1    g259(.A(new_n682), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1981), .B(G1986), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n683), .A2(new_n686), .A3(new_n688), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(G229));
  XOR2_X1   g268(.A(KEYINPUT94), .B(G16), .Z(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n695), .A2(G22), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(G166), .B2(new_n695), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(G1971), .Z(new_n698));
  MUX2_X1   g273(.A(G23), .B(G288), .S(G16), .Z(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT33), .B(G1976), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NOR2_X1   g276(.A1(G6), .A2(G16), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n586), .A2(new_n587), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n702), .B1(new_n703), .B2(G16), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT32), .B(G1981), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n698), .A2(new_n701), .A3(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT34), .Z(new_n708));
  MUX2_X1   g283(.A(G24), .B(G290), .S(new_n695), .Z(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT95), .B(G1986), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n493), .A2(G119), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n479), .A2(G107), .ZN(new_n713));
  OAI21_X1  g288(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n712), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(new_n498), .B2(G131), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT93), .Z(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G29), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G25), .B2(G29), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT35), .B(G1991), .Z(new_n720));
  OAI21_X1  g295(.A(new_n711), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(new_n719), .B2(new_n720), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n708), .A2(new_n722), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT36), .Z(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT30), .B(G28), .ZN(new_n725));
  INV_X1    g300(.A(G29), .ZN(new_n726));
  OR2_X1    g301(.A1(KEYINPUT31), .A2(G11), .ZN(new_n727));
  NAND2_X1  g302(.A1(KEYINPUT31), .A2(G11), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n725), .A2(new_n726), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(new_n625), .B2(new_n726), .ZN(new_n730));
  MUX2_X1   g305(.A(G21), .B(G286), .S(G16), .Z(new_n731));
  AOI21_X1  g306(.A(new_n730), .B1(new_n731), .B2(G1966), .ZN(new_n732));
  INV_X1    g307(.A(G1961), .ZN(new_n733));
  INV_X1    g308(.A(G5), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n734), .A2(G16), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G301), .B2(G16), .ZN(new_n736));
  OAI221_X1 g311(.A(new_n732), .B1(new_n733), .B2(new_n736), .C1(G1966), .C2(new_n731), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT100), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n561), .A2(new_n695), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G19), .B2(new_n695), .ZN(new_n740));
  INV_X1    g315(.A(G1341), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n479), .A2(G103), .A3(G2104), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT25), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n503), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n746));
  INV_X1    g321(.A(G139), .ZN(new_n747));
  OAI221_X1 g322(.A(new_n745), .B1(new_n479), .B2(new_n746), .C1(new_n623), .C2(new_n747), .ZN(new_n748));
  MUX2_X1   g323(.A(G33), .B(new_n748), .S(G29), .Z(new_n749));
  OR2_X1    g324(.A1(new_n749), .A2(G2072), .ZN(new_n750));
  NOR2_X1   g325(.A1(G164), .A2(new_n726), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G27), .B2(new_n726), .ZN(new_n752));
  INV_X1    g327(.A(G2078), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n749), .A2(G2072), .ZN(new_n755));
  NAND4_X1  g330(.A1(new_n742), .A2(new_n750), .A3(new_n754), .A4(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n736), .A2(new_n733), .ZN(new_n757));
  OAI221_X1 g332(.A(new_n757), .B1(new_n752), .B2(new_n753), .C1(new_n740), .C2(new_n741), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(G29), .A2(G32), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n493), .A2(G129), .ZN(new_n761));
  NAND3_X1  g336(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT26), .Z(new_n763));
  NAND2_X1  g338(.A1(new_n481), .A2(G105), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n761), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(new_n765), .ZN(new_n766));
  AND3_X1   g341(.A1(new_n498), .A2(KEYINPUT97), .A3(G141), .ZN(new_n767));
  AOI21_X1  g342(.A(KEYINPUT97), .B1(new_n498), .B2(G141), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT98), .Z(new_n770));
  AOI21_X1  g345(.A(new_n760), .B1(new_n770), .B2(G29), .ZN(new_n771));
  XOR2_X1   g346(.A(KEYINPUT27), .B(G1996), .Z(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n726), .B1(KEYINPUT24), .B2(G34), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(KEYINPUT24), .B2(G34), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n491), .B2(G29), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G2084), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n759), .A2(new_n773), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n726), .A2(G35), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G162), .B2(new_n726), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT29), .Z(new_n781));
  INV_X1    g356(.A(G2090), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(G4), .A2(G16), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n602), .B2(G16), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n785), .A2(G1348), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n694), .A2(G20), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT23), .Z(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G299), .B2(G16), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G1956), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n726), .A2(G26), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT28), .Z(new_n792));
  NAND2_X1  g367(.A1(new_n498), .A2(G140), .ZN(new_n793));
  OAI21_X1  g368(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n794));
  INV_X1    g369(.A(G116), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(G2105), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(new_n493), .B2(G128), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n793), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n792), .B1(new_n798), .B2(G29), .ZN(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT96), .B(G2067), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n785), .A2(G1348), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n786), .A2(new_n790), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  NOR4_X1   g378(.A1(new_n738), .A2(new_n778), .A3(new_n783), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n781), .A2(new_n782), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT101), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n771), .A2(new_n772), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT99), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n804), .A2(new_n806), .A3(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n724), .A2(new_n809), .ZN(G311));
  INV_X1    g385(.A(G311), .ZN(G150));
  AOI22_X1  g386(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n812), .A2(new_n551), .ZN(new_n813));
  INV_X1    g388(.A(G55), .ZN(new_n814));
  INV_X1    g389(.A(G93), .ZN(new_n815));
  OAI221_X1 g390(.A(new_n813), .B1(new_n538), .B2(new_n814), .C1(new_n581), .C2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n816), .A2(G860), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT37), .Z(new_n818));
  NAND2_X1  g393(.A1(new_n602), .A2(G559), .ZN(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n560), .B(new_n816), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n824), .A2(KEYINPUT39), .ZN(new_n825));
  INV_X1    g400(.A(G860), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n824), .B2(KEYINPUT39), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n818), .B1(new_n825), .B2(new_n827), .ZN(G145));
  MUX2_X1   g403(.A(new_n770), .B(new_n769), .S(new_n748), .Z(new_n829));
  XNOR2_X1  g404(.A(new_n798), .B(new_n513), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n829), .B(new_n830), .Z(new_n831));
  OAI21_X1  g406(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n832));
  INV_X1    g407(.A(G118), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n832), .B1(new_n833), .B2(G2105), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(new_n493), .B2(G130), .ZN(new_n835));
  INV_X1    g410(.A(G142), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n835), .B1(new_n623), .B2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT103), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(new_n616), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(new_n717), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT104), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n831), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n491), .B(new_n625), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(G162), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n829), .B(new_n830), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(new_n841), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n843), .A2(new_n845), .A3(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(G37), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n842), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(new_n846), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n845), .B1(new_n852), .B2(new_n843), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT40), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(G395));
  NAND2_X1  g431(.A1(new_n816), .A2(new_n605), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n611), .B(new_n822), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n601), .B(G299), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(KEYINPUT105), .Z(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(KEYINPUT41), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT41), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n859), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n862), .B1(new_n858), .B2(new_n866), .ZN(new_n867));
  XOR2_X1   g442(.A(G303), .B(KEYINPUT106), .Z(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(G290), .ZN(new_n869));
  XNOR2_X1  g444(.A(G288), .B(new_n703), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n869), .B(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT42), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n867), .B(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n857), .B1(new_n873), .B2(new_n605), .ZN(G295));
  OAI21_X1  g449(.A(new_n857), .B1(new_n873), .B2(new_n605), .ZN(G331));
  INV_X1    g450(.A(KEYINPUT43), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n822), .B(G301), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(G168), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n822), .B(G171), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(G286), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(new_n860), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n863), .A2(new_n878), .A3(new_n880), .A4(new_n865), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n882), .A2(new_n883), .A3(new_n871), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(new_n849), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n871), .B1(new_n882), .B2(new_n883), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n876), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n885), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT108), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  AOI211_X1 g465(.A(KEYINPUT108), .B(new_n871), .C1(new_n882), .C2(new_n883), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n888), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n887), .B1(new_n892), .B2(new_n876), .ZN(new_n893));
  OAI21_X1  g468(.A(KEYINPUT43), .B1(new_n885), .B2(new_n886), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(KEYINPUT107), .ZN(new_n895));
  OAI211_X1 g470(.A(new_n888), .B(new_n876), .C1(new_n890), .C2(new_n891), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT107), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n897), .B(KEYINPUT43), .C1(new_n885), .C2(new_n886), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n895), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT44), .ZN(new_n900));
  MUX2_X1   g475(.A(new_n893), .B(new_n899), .S(new_n900), .Z(G397));
  NAND2_X1  g476(.A1(new_n489), .A2(G137), .ZN(new_n902));
  OAI211_X1 g477(.A(G40), .B(new_n902), .C1(new_n482), .C2(new_n484), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  AOI22_X1  g479(.A1(new_n465), .A2(KEYINPUT68), .B1(G113), .B2(G2104), .ZN(new_n905));
  AOI211_X1 g480(.A(KEYINPUT69), .B(new_n479), .C1(new_n905), .C2(new_n468), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n473), .B1(new_n470), .B2(G2105), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n904), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(KEYINPUT110), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT110), .ZN(new_n910));
  OAI211_X1 g485(.A(new_n904), .B(new_n910), .C1(new_n906), .C2(new_n907), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  XOR2_X1   g487(.A(KEYINPUT109), .B(G1384), .Z(new_n913));
  AOI21_X1  g488(.A(KEYINPUT45), .B1(new_n513), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(G1996), .ZN(new_n917));
  AOI21_X1  g492(.A(KEYINPUT46), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n918), .A2(KEYINPUT126), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n918), .A2(KEYINPUT126), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n798), .A2(G2067), .ZN(new_n921));
  INV_X1    g496(.A(G2067), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n793), .A2(new_n922), .A3(new_n797), .ZN(new_n923));
  AND2_X1   g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  AOI211_X1 g500(.A(new_n769), .B(new_n925), .C1(KEYINPUT46), .C2(new_n917), .ZN(new_n926));
  OAI22_X1  g501(.A1(new_n919), .A2(new_n920), .B1(new_n915), .B2(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n927), .B(KEYINPUT47), .ZN(new_n928));
  NOR3_X1   g503(.A1(new_n915), .A2(G1986), .A3(G290), .ZN(new_n929));
  XOR2_X1   g504(.A(new_n929), .B(KEYINPUT48), .Z(new_n930));
  NAND2_X1  g505(.A1(new_n770), .A2(new_n917), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n925), .B1(G1996), .B2(new_n769), .ZN(new_n932));
  OR2_X1    g507(.A1(new_n717), .A2(new_n720), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n717), .A2(new_n720), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n931), .A2(new_n932), .A3(new_n933), .A4(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n930), .B1(new_n936), .B2(new_n915), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n931), .A2(new_n932), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n923), .B1(new_n938), .B2(new_n934), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(new_n916), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n928), .A2(new_n937), .A3(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT63), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT118), .ZN(new_n943));
  AOI21_X1  g518(.A(G1384), .B1(new_n508), .B2(new_n512), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT50), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n910), .B1(new_n475), .B2(new_n904), .ZN(new_n948));
  INV_X1    g523(.A(new_n911), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n943), .B(new_n947), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n944), .A2(new_n945), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n946), .B1(new_n909), .B2(new_n911), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n953), .A2(new_n943), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n952), .A2(new_n954), .A3(G2090), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT111), .B1(new_n944), .B2(KEYINPUT45), .ZN(new_n956));
  INV_X1    g531(.A(G1384), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n489), .A2(G138), .ZN(new_n958));
  AOI22_X1  g533(.A1(new_n958), .A2(KEYINPUT4), .B1(new_n502), .B2(new_n503), .ZN(new_n959));
  INV_X1    g534(.A(new_n512), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n957), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT111), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT45), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n961), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n513), .A2(KEYINPUT45), .A3(new_n913), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n956), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(G1971), .B1(new_n966), .B2(new_n912), .ZN(new_n967));
  OAI21_X1  g542(.A(G8), .B1(new_n955), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(G303), .A2(G8), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT55), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OR2_X1    g546(.A1(new_n971), .A2(KEYINPUT113), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n969), .A2(new_n970), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n971), .A2(KEYINPUT113), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n968), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(G1981), .ZN(new_n978));
  OAI21_X1  g553(.A(KEYINPUT116), .B1(new_n703), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT116), .ZN(new_n980));
  NAND3_X1  g555(.A1(G305), .A2(new_n980), .A3(G1981), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n586), .A2(new_n587), .A3(new_n978), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT115), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n983), .B(new_n984), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n982), .A2(KEYINPUT49), .A3(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT49), .B1(new_n982), .B2(new_n985), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n912), .A2(new_n944), .ZN(new_n989));
  AOI21_X1  g564(.A(KEYINPUT114), .B1(new_n989), .B2(G8), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n961), .B1(new_n909), .B2(new_n911), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT114), .ZN(new_n992));
  INV_X1    g567(.A(G8), .ZN(new_n993));
  NOR3_X1   g568(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n988), .B1(new_n990), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(KEYINPUT117), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n989), .A2(KEYINPUT114), .A3(G8), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n992), .B1(new_n991), .B2(new_n993), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT117), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n999), .A2(new_n1000), .A3(new_n988), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n996), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n1003));
  INV_X1    g578(.A(G1976), .ZN(new_n1004));
  NOR2_X1   g579(.A1(G288), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1003), .B1(new_n999), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G288), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1003), .B1(new_n1008), .B2(G1976), .ZN(new_n1009));
  AOI211_X1 g584(.A(new_n1005), .B(new_n1009), .C1(new_n997), .C2(new_n998), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n953), .A2(new_n782), .A3(new_n951), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT112), .B1(new_n1013), .B2(new_n967), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT112), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n956), .A2(new_n964), .A3(new_n965), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1016), .B1(new_n911), .B2(new_n909), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n1015), .B(new_n1012), .C1(new_n1017), .C2(G1971), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1014), .A2(G8), .A3(new_n1018), .A4(new_n975), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n977), .A2(new_n1002), .A3(new_n1011), .A4(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n961), .B(KEYINPUT45), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n912), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(G1966), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G2084), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n953), .A2(new_n1025), .A3(new_n951), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1027), .A2(G8), .A3(G168), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n942), .B1(new_n1020), .B2(new_n1028), .ZN(new_n1029));
  AND2_X1   g604(.A1(new_n1002), .A2(new_n1011), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1014), .A2(G8), .A3(new_n1018), .ZN(new_n1031));
  AOI211_X1 g606(.A(new_n942), .B(new_n1028), .C1(new_n1031), .C2(new_n976), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1030), .A2(new_n1032), .A3(new_n1019), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1029), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n966), .A2(new_n912), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1035), .B1(new_n1036), .B2(G2078), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1035), .A2(G2078), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n912), .A2(new_n1021), .A3(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n912), .A2(new_n947), .A3(new_n951), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(new_n733), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1037), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(G171), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1020), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(G8), .B1(new_n1027), .B2(G286), .ZN(new_n1045));
  AOI21_X1  g620(.A(G168), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT51), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT62), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT51), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1049), .B(G8), .C1(new_n1027), .C2(G286), .ZN(new_n1050));
  AND3_X1   g625(.A1(new_n1047), .A2(new_n1048), .A3(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1048), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1044), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1002), .A2(new_n1004), .A3(new_n1008), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(new_n985), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1019), .ZN(new_n1057));
  AOI22_X1  g632(.A1(new_n1056), .A2(new_n999), .B1(new_n1030), .B2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1034), .A2(new_n1054), .A3(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT61), .ZN(new_n1060));
  INV_X1    g635(.A(G1956), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1061), .B1(new_n952), .B2(new_n954), .ZN(new_n1062));
  XNOR2_X1  g637(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(G299), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n574), .A2(new_n576), .A3(new_n1063), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  XOR2_X1   g642(.A(KEYINPUT56), .B(G2072), .Z(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1067), .B1(new_n1017), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1060), .B1(new_n1062), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n951), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1072), .B1(new_n953), .B2(new_n943), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT118), .ZN(new_n1075));
  AOI21_X1  g650(.A(G1956), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n966), .A2(new_n912), .A3(new_n1069), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1067), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  AND3_X1   g654(.A1(new_n1071), .A2(new_n1079), .A3(KEYINPUT121), .ZN(new_n1080));
  AOI21_X1  g655(.A(KEYINPUT121), .B1(new_n1071), .B2(new_n1079), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1067), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1083), .B1(new_n1062), .B2(new_n1077), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1077), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1076), .A2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1060), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1036), .A2(G1996), .ZN(new_n1088));
  XNOR2_X1  g663(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n1089));
  XNOR2_X1  g664(.A(new_n1089), .B(new_n741), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n991), .A2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n561), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(KEYINPUT59), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1094), .B(new_n561), .C1(new_n1088), .C2(new_n1091), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1087), .A2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(KEYINPUT122), .B1(new_n1082), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT121), .ZN(new_n1099));
  OAI21_X1  g674(.A(KEYINPUT61), .B1(new_n1076), .B2(new_n1085), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1099), .B1(new_n1084), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1071), .A2(new_n1079), .A3(KEYINPUT121), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT122), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1103), .A2(new_n1104), .A3(new_n1087), .A4(new_n1096), .ZN(new_n1105));
  INV_X1    g680(.A(G1348), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1040), .A2(new_n1106), .B1(new_n922), .B2(new_n991), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(KEYINPUT60), .ZN(new_n1108));
  XNOR2_X1  g683(.A(new_n1108), .B(new_n602), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1109), .B1(KEYINPUT60), .B2(new_n1107), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1098), .A2(new_n1105), .A3(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1079), .B1(new_n601), .B2(new_n1107), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1112), .B1(new_n1076), .B2(new_n1085), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n903), .B1(G2105), .B2(new_n470), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n914), .B1(KEYINPUT123), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT124), .ZN(new_n1117));
  OR2_X1    g692(.A1(new_n1115), .A2(KEYINPUT123), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1116), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1117), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n965), .B(new_n1038), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1121), .A2(new_n1037), .A3(new_n1041), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1043), .B1(new_n1122), .B2(G171), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT54), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1047), .A2(new_n1050), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1042), .A2(G171), .ZN(new_n1128));
  XOR2_X1   g703(.A(new_n1128), .B(KEYINPUT125), .Z(new_n1129));
  AOI21_X1  g704(.A(new_n1124), .B1(new_n1122), .B2(G171), .ZN(new_n1130));
  AOI211_X1 g705(.A(new_n1020), .B(new_n1127), .C1(new_n1129), .C2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1059), .B1(new_n1114), .B2(new_n1131), .ZN(new_n1132));
  XOR2_X1   g707(.A(G290), .B(G1986), .Z(new_n1133));
  AOI21_X1  g708(.A(new_n915), .B1(new_n936), .B2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n941), .B1(new_n1132), .B2(new_n1134), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g710(.A(KEYINPUT127), .ZN(new_n1137));
  NAND2_X1  g711(.A1(new_n643), .A2(new_n459), .ZN(new_n1138));
  NOR2_X1   g712(.A1(G227), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g713(.A(new_n1137), .B1(new_n692), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g714(.A(new_n1139), .ZN(new_n1141));
  AOI211_X1 g715(.A(KEYINPUT127), .B(new_n1141), .C1(new_n690), .C2(new_n691), .ZN(new_n1142));
  OAI22_X1  g716(.A1(new_n1140), .A2(new_n1142), .B1(new_n850), .B2(new_n853), .ZN(new_n1143));
  AND2_X1   g717(.A1(new_n895), .A2(new_n896), .ZN(new_n1144));
  AOI21_X1  g718(.A(new_n1143), .B1(new_n1144), .B2(new_n898), .ZN(G308));
  OAI221_X1 g719(.A(new_n899), .B1(new_n853), .B2(new_n850), .C1(new_n1140), .C2(new_n1142), .ZN(G225));
endmodule


