//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 1 1 1 1 0 1 1 0 0 0 0 0 0 0 0 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 1 1 1 1 0 0 0 0 0 1 1 0 0 1 1 0 0 1 0 0 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:19 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n815,
    new_n816, new_n817, new_n818, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT77), .B(G125), .ZN(new_n190));
  NOR3_X1   g004(.A1(new_n190), .A2(KEYINPUT16), .A3(G140), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G140), .ZN(new_n193));
  INV_X1    g007(.A(G125), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT77), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT77), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G125), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n193), .B1(new_n195), .B2(new_n197), .ZN(new_n198));
  NOR2_X1   g012(.A1(G125), .A2(G140), .ZN(new_n199));
  OAI211_X1 g013(.A(KEYINPUT78), .B(KEYINPUT16), .C1(new_n198), .C2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(new_n199), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n202), .B1(new_n190), .B2(new_n193), .ZN(new_n203));
  AOI21_X1  g017(.A(KEYINPUT78), .B1(new_n203), .B2(KEYINPUT16), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n192), .B1(new_n201), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OAI211_X1 g021(.A(G146), .B(new_n192), .C1(new_n201), .C2(new_n204), .ZN(new_n208));
  NOR2_X1   g022(.A1(G237), .A2(G953), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G214), .ZN(new_n210));
  INV_X1    g024(.A(G143), .ZN(new_n211));
  XNOR2_X1  g025(.A(new_n210), .B(new_n211), .ZN(new_n212));
  AOI21_X1  g026(.A(KEYINPUT95), .B1(new_n212), .B2(G131), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n210), .A2(new_n211), .ZN(new_n214));
  AOI21_X1  g028(.A(G143), .B1(new_n209), .B2(G214), .ZN(new_n215));
  OAI21_X1  g029(.A(G131), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT95), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT17), .B1(new_n213), .B2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n212), .A2(KEYINPUT95), .A3(G131), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n216), .A2(new_n217), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n214), .A2(new_n215), .ZN(new_n222));
  INV_X1    g036(.A(G131), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT17), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n220), .A2(new_n221), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n207), .A2(new_n208), .A3(new_n219), .A4(new_n226), .ZN(new_n227));
  XNOR2_X1  g041(.A(G113), .B(G122), .ZN(new_n228));
  INV_X1    g042(.A(G104), .ZN(new_n229));
  XNOR2_X1  g043(.A(new_n228), .B(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT18), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n222), .B1(new_n231), .B2(new_n223), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n212), .A2(KEYINPUT18), .A3(G131), .ZN(new_n233));
  NAND2_X1  g047(.A1(G125), .A2(G140), .ZN(new_n234));
  AND3_X1   g048(.A1(new_n202), .A2(KEYINPUT79), .A3(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(KEYINPUT79), .B1(new_n202), .B2(new_n234), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT65), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(new_n206), .ZN(new_n239));
  NAND2_X1  g053(.A1(KEYINPUT65), .A2(G146), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n237), .A2(new_n241), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n203), .A2(new_n206), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n232), .B(new_n233), .C1(new_n242), .C2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n227), .A2(new_n230), .A3(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n220), .A2(new_n221), .A3(new_n224), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n247), .B1(new_n235), .B2(new_n236), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n195), .A2(new_n197), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n199), .B1(new_n249), .B2(G140), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT19), .ZN(new_n251));
  INV_X1    g065(.A(new_n240), .ZN(new_n252));
  NOR2_X1   g066(.A1(KEYINPUT65), .A2(G146), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n248), .A2(new_n251), .A3(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n208), .A2(new_n246), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(new_n244), .ZN(new_n257));
  INV_X1    g071(.A(new_n230), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n245), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(G475), .A2(G902), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT20), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n245), .A2(new_n259), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT20), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n264), .A2(new_n265), .A3(new_n261), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(G902), .ZN(new_n268));
  XNOR2_X1  g082(.A(G128), .B(G143), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT13), .ZN(new_n270));
  INV_X1    g084(.A(G128), .ZN(new_n271));
  NOR3_X1   g085(.A1(new_n271), .A2(KEYINPUT13), .A3(G143), .ZN(new_n272));
  INV_X1    g086(.A(G134), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI22_X1  g088(.A1(new_n270), .A2(new_n274), .B1(new_n273), .B2(new_n269), .ZN(new_n275));
  INV_X1    g089(.A(G116), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n276), .A2(G122), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  AND2_X1   g092(.A1(KEYINPUT69), .A2(G116), .ZN(new_n279));
  NOR2_X1   g093(.A1(KEYINPUT69), .A2(G116), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(KEYINPUT97), .B1(new_n281), .B2(G122), .ZN(new_n282));
  OR2_X1    g096(.A1(KEYINPUT69), .A2(G116), .ZN(new_n283));
  NAND2_X1  g097(.A1(KEYINPUT69), .A2(G116), .ZN(new_n284));
  AND4_X1   g098(.A1(KEYINPUT97), .A2(new_n283), .A3(G122), .A4(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n278), .B1(new_n282), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(G107), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n283), .A2(G122), .A3(new_n284), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT97), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n281), .A2(KEYINPUT97), .A3(G122), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G107), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n292), .A2(new_n293), .A3(new_n278), .ZN(new_n294));
  AND3_X1   g108(.A1(new_n287), .A2(KEYINPUT98), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(KEYINPUT98), .B1(new_n287), .B2(new_n294), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n275), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G217), .ZN(new_n298));
  NOR3_X1   g112(.A1(new_n187), .A2(new_n298), .A3(G953), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n277), .B1(new_n292), .B2(KEYINPUT14), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT14), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n290), .A2(new_n291), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n293), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT99), .ZN(new_n304));
  XNOR2_X1  g118(.A(new_n269), .B(new_n273), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n294), .A2(new_n305), .ZN(new_n306));
  NOR3_X1   g120(.A1(new_n303), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(KEYINPUT14), .B1(new_n282), .B2(new_n285), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(new_n302), .A3(new_n278), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G107), .ZN(new_n310));
  AND2_X1   g124(.A1(new_n294), .A2(new_n305), .ZN(new_n311));
  AOI21_X1  g125(.A(KEYINPUT99), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  OAI211_X1 g126(.A(new_n297), .B(new_n299), .C1(new_n307), .C2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n304), .B1(new_n303), .B2(new_n306), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n310), .A2(new_n311), .A3(KEYINPUT99), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n299), .B1(new_n317), .B2(new_n297), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n268), .B1(new_n314), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G478), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n320), .A2(KEYINPUT15), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n245), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n230), .B1(new_n227), .B2(new_n244), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n268), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G475), .ZN(new_n326));
  OAI221_X1 g140(.A(new_n268), .B1(KEYINPUT15), .B2(new_n320), .C1(new_n314), .C2(new_n318), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n267), .A2(new_n322), .A3(new_n326), .A4(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT11), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n329), .B1(new_n273), .B2(G137), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n273), .A2(G137), .ZN(new_n331));
  INV_X1    g145(.A(G137), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(KEYINPUT11), .A3(G134), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n330), .A2(new_n331), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G131), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n330), .A2(new_n333), .A3(new_n223), .A4(new_n331), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT86), .B1(new_n293), .B2(G104), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT86), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n340), .A2(new_n229), .A3(G107), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n293), .A2(G104), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n339), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G101), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT87), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n293), .A2(G104), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT3), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n348), .A2(KEYINPUT83), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n347), .B1(new_n349), .B2(new_n342), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT83), .ZN(new_n351));
  OAI22_X1  g165(.A1(new_n351), .A2(KEYINPUT3), .B1(new_n229), .B2(G107), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(KEYINPUT3), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G101), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n350), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n343), .A2(KEYINPUT87), .A3(G101), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n346), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n239), .A2(G143), .A3(new_n240), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(KEYINPUT1), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G128), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n211), .A2(G146), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n363), .B1(new_n254), .B2(G143), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n211), .A2(G146), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n359), .A2(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n271), .A2(KEYINPUT1), .ZN(new_n367));
  AOI22_X1  g181(.A1(new_n361), .A2(new_n364), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n358), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n359), .A2(new_n365), .A3(new_n367), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n271), .B1(new_n363), .B2(KEYINPUT1), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n370), .B1(new_n366), .B2(new_n371), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n372), .A2(new_n356), .A3(new_n357), .A4(new_n346), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n338), .B1(new_n369), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(KEYINPUT89), .B1(new_n374), .B2(KEYINPUT12), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NOR3_X1   g190(.A1(new_n374), .A2(KEYINPUT89), .A3(KEYINPUT12), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n374), .A2(KEYINPUT88), .A3(KEYINPUT12), .ZN(new_n378));
  AOI21_X1  g192(.A(KEYINPUT88), .B1(new_n374), .B2(KEYINPUT12), .ZN(new_n379));
  OAI22_X1  g193(.A1(new_n376), .A2(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n348), .A2(KEYINPUT83), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n349), .B1(new_n342), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n229), .A2(G107), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n229), .A2(G107), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n383), .B1(new_n384), .B2(new_n353), .ZN(new_n385));
  OAI21_X1  g199(.A(KEYINPUT84), .B1(new_n382), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT84), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n350), .A2(new_n354), .A3(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT4), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n386), .A2(new_n388), .A3(new_n389), .A4(G101), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(KEYINPUT85), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n349), .A2(new_n342), .ZN(new_n392));
  AOI22_X1  g206(.A1(KEYINPUT83), .A2(new_n348), .B1(new_n293), .B2(G104), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n392), .B(new_n383), .C1(new_n393), .C2(new_n349), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n355), .B1(new_n394), .B2(KEYINPUT84), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT85), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n395), .A2(new_n396), .A3(new_n389), .A4(new_n388), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n391), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n359), .A2(KEYINPUT0), .A3(G128), .A4(new_n365), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n362), .B1(new_n241), .B2(new_n211), .ZN(new_n400));
  NAND2_X1  g214(.A1(KEYINPUT0), .A2(G128), .ZN(new_n401));
  OAI21_X1  g215(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NOR3_X1   g217(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n401), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n399), .B1(new_n400), .B2(new_n405), .ZN(new_n406));
  AND2_X1   g220(.A1(new_n356), .A2(KEYINPUT4), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n386), .A2(new_n388), .A3(G101), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n406), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n398), .A2(new_n409), .ZN(new_n410));
  AND3_X1   g224(.A1(new_n346), .A2(new_n356), .A3(new_n357), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n271), .B1(new_n359), .B2(KEYINPUT1), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n370), .B1(new_n412), .B2(new_n400), .ZN(new_n413));
  AND2_X1   g227(.A1(new_n413), .A2(KEYINPUT10), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT10), .ZN(new_n415));
  AOI22_X1  g229(.A1(new_n411), .A2(new_n414), .B1(new_n373), .B2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n410), .A2(new_n416), .A3(new_n338), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n380), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(G110), .B(G140), .ZN(new_n419));
  INV_X1    g233(.A(G953), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n420), .A2(G227), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n419), .B(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n410), .A2(new_n416), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n337), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT90), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n423), .A2(KEYINPUT90), .A3(new_n337), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n422), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n417), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  AOI22_X1  g245(.A1(new_n418), .A2(new_n422), .B1(new_n428), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(G469), .B1(new_n432), .B2(G902), .ZN(new_n433));
  INV_X1    g247(.A(G469), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n429), .B1(new_n428), .B2(new_n417), .ZN(new_n435));
  OR2_X1    g249(.A1(new_n378), .A2(new_n379), .ZN(new_n436));
  INV_X1    g250(.A(new_n377), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n375), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n430), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n434), .B(new_n268), .C1(new_n435), .C2(new_n439), .ZN(new_n440));
  AOI211_X1 g254(.A(new_n189), .B(new_n328), .C1(new_n433), .C2(new_n440), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n338), .A2(new_n406), .ZN(new_n442));
  XNOR2_X1  g256(.A(KEYINPUT2), .B(G113), .ZN(new_n443));
  INV_X1    g257(.A(G119), .ZN(new_n444));
  NOR3_X1   g258(.A1(new_n279), .A2(new_n280), .A3(new_n444), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n276), .A2(G119), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n443), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  XOR2_X1   g261(.A(KEYINPUT2), .B(G113), .Z(new_n448));
  NAND3_X1  g262(.A1(new_n283), .A2(G119), .A3(new_n284), .ZN(new_n449));
  INV_X1    g263(.A(new_n446), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n447), .A2(KEYINPUT70), .A3(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT70), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n453), .B(new_n443), .C1(new_n445), .C2(new_n446), .ZN(new_n454));
  AND2_X1   g268(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(KEYINPUT67), .B1(new_n273), .B2(G137), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT67), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n457), .A2(new_n332), .A3(G134), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n456), .A2(new_n458), .A3(new_n331), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(G131), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT68), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n459), .A2(KEYINPUT68), .A3(G131), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n462), .A2(new_n336), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n368), .B1(KEYINPUT71), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT71), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n462), .A2(new_n466), .A3(new_n336), .A4(new_n463), .ZN(new_n467));
  AOI211_X1 g281(.A(new_n442), .B(new_n455), .C1(new_n465), .C2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n452), .A2(new_n454), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n464), .A2(KEYINPUT71), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n470), .A2(new_n467), .A3(new_n413), .ZN(new_n471));
  INV_X1    g285(.A(new_n442), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(KEYINPUT28), .B1(new_n468), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n442), .B1(new_n465), .B2(new_n467), .ZN(new_n475));
  AOI21_X1  g289(.A(KEYINPUT28), .B1(new_n475), .B2(new_n469), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n209), .A2(G210), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT27), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n479), .B(new_n480), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(KEYINPUT26), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(G101), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT26), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n481), .B(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n355), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT29), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n268), .B1(new_n478), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(KEYINPUT76), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT76), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n492), .B(new_n268), .C1(new_n478), .C2(new_n489), .ZN(new_n493));
  OAI21_X1  g307(.A(KEYINPUT66), .B1(new_n338), .B2(new_n406), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n413), .A2(new_n336), .A3(new_n463), .A4(new_n462), .ZN(new_n495));
  OR2_X1    g309(.A1(new_n400), .A2(new_n405), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT66), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n496), .A2(new_n497), .A3(new_n337), .A4(new_n399), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n494), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT30), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n469), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n471), .A2(KEYINPUT30), .A3(new_n472), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n471), .A2(new_n472), .A3(new_n469), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n505), .A2(KEYINPUT75), .A3(new_n487), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT75), .ZN(new_n507));
  AOI22_X1  g321(.A1(new_n501), .A2(new_n502), .B1(new_n475), .B2(new_n469), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n507), .B1(new_n508), .B2(new_n488), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n499), .A2(new_n455), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n504), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT73), .B(KEYINPUT28), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n513), .A2(new_n477), .A3(new_n488), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT29), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n506), .A2(new_n509), .A3(new_n514), .A4(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n491), .A2(new_n493), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(G472), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT32), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n487), .B1(new_n475), .B2(new_n469), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n503), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(KEYINPUT31), .ZN(new_n522));
  INV_X1    g336(.A(new_n512), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n523), .B1(new_n504), .B2(new_n510), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n487), .B1(new_n524), .B2(new_n476), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT72), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT31), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n503), .A2(new_n520), .A3(new_n527), .A4(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n503), .A2(new_n520), .A3(new_n528), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT72), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n526), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(G472), .A2(G902), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n533), .B(KEYINPUT74), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n519), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n513), .A2(new_n477), .ZN(new_n536));
  AOI22_X1  g350(.A1(new_n536), .A2(new_n487), .B1(KEYINPUT31), .B2(new_n521), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n531), .A2(new_n529), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n534), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n539), .A2(KEYINPUT32), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n518), .A2(new_n535), .A3(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(G214), .B1(G237), .B2(G902), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(G952), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n545), .A2(G953), .ZN(new_n546));
  NAND2_X1  g360(.A1(G234), .A2(G237), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(KEYINPUT21), .B(G898), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n547), .A2(G902), .A3(G953), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n548), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n449), .A2(KEYINPUT5), .A3(new_n450), .ZN(new_n554));
  INV_X1    g368(.A(G113), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT5), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n555), .B1(new_n446), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n451), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n411), .A2(new_n560), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n391), .A2(new_n397), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n407), .A2(new_n408), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n455), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n561), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(G110), .B(G122), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n566), .B(new_n561), .C1(new_n562), .C2(new_n564), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n568), .A2(KEYINPUT6), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n413), .A2(new_n190), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n571), .B1(new_n406), .B2(new_n190), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n420), .A2(G224), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n572), .B(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT91), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n469), .B1(new_n408), .B2(new_n407), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n398), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n566), .B1(new_n577), .B2(new_n561), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT6), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n575), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  AOI22_X1  g394(.A1(new_n576), .A2(new_n398), .B1(new_n411), .B2(new_n560), .ZN(new_n581));
  NOR4_X1   g395(.A1(new_n581), .A2(KEYINPUT91), .A3(KEYINPUT6), .A4(new_n566), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n570), .B(new_n574), .C1(new_n580), .C2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT93), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT92), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n554), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n449), .A2(KEYINPUT92), .A3(KEYINPUT5), .A4(new_n450), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n586), .A2(new_n557), .A3(new_n587), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n411), .A2(new_n584), .A3(new_n451), .A4(new_n588), .ZN(new_n589));
  AND3_X1   g403(.A1(new_n586), .A2(new_n557), .A3(new_n587), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n346), .A2(new_n451), .A3(new_n356), .A4(new_n357), .ZN(new_n591));
  OAI21_X1  g405(.A(KEYINPUT93), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n358), .A2(new_n559), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n589), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n566), .B(KEYINPUT8), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT7), .ZN(new_n597));
  INV_X1    g411(.A(new_n573), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n572), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n598), .A2(new_n597), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n571), .B(new_n600), .C1(new_n406), .C2(new_n190), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n596), .A2(new_n569), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(KEYINPUT94), .B1(new_n603), .B2(new_n268), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n603), .A2(KEYINPUT94), .A3(new_n268), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n583), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(G210), .B1(G237), .B2(G902), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n583), .B(new_n607), .C1(new_n604), .C2(new_n605), .ZN(new_n610));
  AOI211_X1 g424(.A(new_n544), .B(new_n553), .C1(new_n609), .C2(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n298), .B1(G234), .B2(new_n268), .ZN(new_n612));
  NOR2_X1   g426(.A1(KEYINPUT81), .A2(KEYINPUT25), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT22), .B(G137), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(KEYINPUT80), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n420), .A2(G221), .A3(G234), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT23), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n620), .B1(new_n444), .B2(G128), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n271), .A2(KEYINPUT23), .A3(G119), .ZN(new_n622));
  OAI211_X1 g436(.A(new_n621), .B(new_n622), .C1(G119), .C2(new_n271), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(G110), .ZN(new_n624));
  XOR2_X1   g438(.A(KEYINPUT24), .B(G110), .Z(new_n625));
  XNOR2_X1  g439(.A(G119), .B(G128), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n628), .B1(new_n207), .B2(new_n208), .ZN(new_n629));
  OAI22_X1  g443(.A1(new_n623), .A2(G110), .B1(new_n626), .B2(new_n625), .ZN(new_n630));
  INV_X1    g444(.A(new_n242), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n208), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n619), .B1(new_n629), .B2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n628), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT78), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT16), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n636), .B1(new_n250), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n200), .ZN(new_n639));
  AOI21_X1  g453(.A(G146), .B1(new_n639), .B2(new_n192), .ZN(new_n640));
  AOI211_X1 g454(.A(new_n206), .B(new_n191), .C1(new_n638), .C2(new_n200), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n635), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n642), .A2(new_n632), .A3(new_n618), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n634), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n614), .B1(new_n644), .B2(new_n268), .ZN(new_n645));
  AOI211_X1 g459(.A(G902), .B(new_n613), .C1(new_n634), .C2(new_n643), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n612), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n612), .A2(G902), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n648), .B(KEYINPUT82), .Z(new_n649));
  NAND2_X1  g463(.A1(new_n644), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n441), .A2(new_n542), .A3(new_n611), .A4(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G101), .ZN(G3));
  AOI211_X1 g468(.A(new_n651), .B(new_n189), .C1(new_n433), .C2(new_n440), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n539), .A2(new_n268), .ZN(new_n656));
  AOI22_X1  g470(.A1(new_n656), .A2(G472), .B1(new_n540), .B2(new_n539), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n611), .ZN(new_n659));
  INV_X1    g473(.A(new_n318), .ZN(new_n660));
  AOI21_X1  g474(.A(KEYINPUT33), .B1(new_n660), .B2(new_n313), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT33), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n297), .B1(new_n307), .B2(new_n312), .ZN(new_n663));
  INV_X1    g477(.A(new_n299), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT100), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n313), .A2(new_n666), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n317), .A2(KEYINPUT100), .A3(new_n297), .A4(new_n299), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n665), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(KEYINPUT101), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT101), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n665), .A2(new_n667), .A3(new_n671), .A4(new_n668), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n661), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n320), .A2(G902), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n319), .A2(new_n320), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI22_X1  g491(.A1(new_n263), .A2(new_n266), .B1(G475), .B2(new_n325), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n658), .A2(new_n659), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT34), .B(G104), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G6));
  INV_X1    g497(.A(KEYINPUT103), .ZN(new_n684));
  INV_X1    g498(.A(new_n610), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n603), .A2(new_n268), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT94), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n603), .A2(KEYINPUT94), .A3(new_n268), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n607), .B1(new_n690), .B2(new_n583), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n543), .B1(new_n685), .B2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT102), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n263), .A2(new_n693), .A3(new_n266), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n265), .B1(new_n264), .B2(new_n261), .ZN(new_n695));
  AOI211_X1 g509(.A(KEYINPUT20), .B(new_n262), .C1(new_n245), .C2(new_n259), .ZN(new_n696));
  OAI21_X1  g510(.A(KEYINPUT102), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n322), .A2(new_n327), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n698), .A2(new_n552), .A3(new_n326), .A4(new_n699), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n684), .B1(new_n692), .B2(new_n700), .ZN(new_n701));
  OR3_X1    g515(.A1(new_n692), .A2(new_n684), .A3(new_n700), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n658), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT35), .B(G107), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G9));
  NAND2_X1  g519(.A1(new_n642), .A2(new_n632), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n618), .A2(KEYINPUT36), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n649), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n647), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n441), .A2(new_n611), .A3(new_n657), .A4(new_n710), .ZN(new_n711));
  XOR2_X1   g525(.A(KEYINPUT37), .B(G110), .Z(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G12));
  INV_X1    g527(.A(KEYINPUT105), .ZN(new_n714));
  XOR2_X1   g528(.A(KEYINPUT104), .B(G900), .Z(new_n715));
  OR2_X1    g529(.A1(new_n715), .A2(new_n551), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n548), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n698), .A2(new_n326), .A3(new_n699), .A4(new_n717), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n714), .B1(new_n692), .B2(new_n718), .ZN(new_n719));
  AND4_X1   g533(.A1(new_n326), .A2(new_n698), .A3(new_n699), .A4(new_n717), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n544), .B1(new_n609), .B2(new_n610), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n720), .A2(new_n721), .A3(KEYINPUT105), .ZN(new_n722));
  AND2_X1   g536(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n189), .B1(new_n433), .B2(new_n440), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n542), .A2(new_n724), .A3(new_n710), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G128), .ZN(G30));
  XOR2_X1   g542(.A(new_n717), .B(KEYINPUT107), .Z(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(KEYINPUT39), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n724), .A2(new_n730), .ZN(new_n731));
  XOR2_X1   g545(.A(new_n731), .B(KEYINPUT40), .Z(new_n732));
  NAND2_X1  g546(.A1(new_n609), .A2(new_n610), .ZN(new_n733));
  XOR2_X1   g547(.A(new_n733), .B(KEYINPUT38), .Z(new_n734));
  AOI21_X1  g548(.A(KEYINPUT32), .B1(new_n539), .B2(new_n540), .ZN(new_n735));
  AOI211_X1 g549(.A(new_n519), .B(new_n534), .C1(new_n537), .C2(new_n538), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n505), .A2(new_n488), .ZN(new_n738));
  OR2_X1    g552(.A1(new_n468), .A2(new_n473), .ZN(new_n739));
  OAI211_X1 g553(.A(new_n738), .B(new_n268), .C1(new_n488), .C2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(G472), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT106), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n741), .B(new_n742), .ZN(new_n743));
  AND2_X1   g557(.A1(new_n737), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n678), .B1(new_n322), .B2(new_n327), .ZN(new_n745));
  INV_X1    g559(.A(new_n710), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n745), .A2(new_n543), .A3(new_n746), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n734), .A2(new_n744), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n732), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G143), .ZN(G45));
  INV_X1    g564(.A(KEYINPUT108), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n677), .A2(new_n721), .A3(new_n679), .A4(new_n717), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n751), .B1(new_n725), .B2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(new_n674), .ZN(new_n754));
  AOI211_X1 g568(.A(new_n661), .B(new_n754), .C1(new_n670), .C2(new_n672), .ZN(new_n755));
  INV_X1    g569(.A(new_n676), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n679), .B(new_n717), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n757), .A2(new_n692), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n746), .B1(new_n737), .B2(new_n518), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n758), .A2(new_n759), .A3(KEYINPUT108), .A4(new_n724), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n753), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G146), .ZN(G48));
  AOI21_X1  g576(.A(KEYINPUT90), .B1(new_n423), .B2(new_n337), .ZN(new_n763));
  AOI211_X1 g577(.A(new_n425), .B(new_n338), .C1(new_n410), .C2(new_n416), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n417), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  AOI22_X1  g579(.A1(new_n765), .A2(new_n422), .B1(new_n431), .B2(new_n380), .ZN(new_n766));
  OAI21_X1  g580(.A(G469), .B1(new_n766), .B2(G902), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n767), .A2(new_n440), .A3(new_n188), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(KEYINPUT109), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT109), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n767), .A2(new_n440), .A3(new_n770), .A4(new_n188), .ZN(new_n771));
  AND4_X1   g585(.A1(new_n542), .A2(new_n769), .A3(new_n652), .A4(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n659), .A2(new_n680), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(KEYINPUT41), .B(G113), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n774), .B(new_n775), .ZN(G15));
  NAND2_X1  g590(.A1(new_n702), .A2(new_n701), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n772), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G116), .ZN(G18));
  NOR4_X1   g593(.A1(new_n692), .A2(new_n768), .A3(new_n553), .A4(new_n328), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n759), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G119), .ZN(G21));
  XOR2_X1   g596(.A(KEYINPUT110), .B(G472), .Z(new_n783));
  AOI21_X1  g597(.A(new_n783), .B1(new_n539), .B2(new_n268), .ZN(new_n784));
  AOI22_X1  g598(.A1(new_n478), .A2(new_n487), .B1(KEYINPUT31), .B2(new_n521), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n534), .B1(new_n785), .B2(new_n538), .ZN(new_n786));
  NOR4_X1   g600(.A1(new_n784), .A2(new_n651), .A3(new_n786), .A4(new_n553), .ZN(new_n787));
  AND3_X1   g601(.A1(new_n787), .A2(new_n769), .A3(new_n771), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n679), .A2(new_n699), .ZN(new_n789));
  OAI21_X1  g603(.A(KEYINPUT111), .B1(new_n692), .B2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT111), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n721), .A2(new_n791), .A3(new_n745), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n788), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G122), .ZN(G24));
  NOR2_X1   g609(.A1(new_n692), .A2(new_n768), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n756), .B1(new_n673), .B2(new_n674), .ZN(new_n797));
  INV_X1    g611(.A(new_n717), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n797), .A2(new_n678), .A3(new_n798), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n784), .A2(new_n746), .A3(new_n786), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n796), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G125), .ZN(G27));
  INV_X1    g616(.A(KEYINPUT42), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n685), .A2(new_n691), .A3(new_n544), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n542), .A2(new_n652), .A3(new_n724), .A4(new_n804), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n803), .B1(new_n805), .B2(new_n757), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n433), .A2(new_n440), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(new_n188), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n609), .A2(new_n543), .A3(new_n610), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n651), .B1(new_n737), .B2(new_n518), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n810), .A2(new_n811), .A3(KEYINPUT42), .A4(new_n799), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n806), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(G131), .ZN(G33));
  INV_X1    g628(.A(KEYINPUT112), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n815), .B1(new_n805), .B2(new_n718), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n810), .A2(new_n811), .A3(KEYINPUT112), .A4(new_n720), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(G134), .ZN(G36));
  NOR2_X1   g633(.A1(new_n797), .A2(new_n679), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(KEYINPUT43), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n657), .A2(new_n746), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT44), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n821), .A2(KEYINPUT44), .A3(new_n822), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n825), .A2(new_n804), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(G469), .A2(G902), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n431), .B1(new_n763), .B2(new_n764), .ZN(new_n829));
  INV_X1    g643(.A(new_n417), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n830), .B1(new_n436), .B2(new_n438), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n829), .B(KEYINPUT45), .C1(new_n831), .C2(new_n429), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(KEYINPUT113), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT113), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n432), .A2(new_n834), .A3(KEYINPUT45), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n432), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT45), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n434), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT114), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n836), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n840), .B1(new_n836), .B2(new_n839), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n828), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT46), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI211_X1 g659(.A(KEYINPUT46), .B(new_n828), .C1(new_n841), .C2(new_n842), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n845), .A2(new_n440), .A3(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n847), .A2(new_n188), .A3(new_n730), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n827), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(new_n332), .ZN(G39));
  NAND2_X1  g664(.A1(new_n847), .A2(new_n188), .ZN(new_n851));
  XNOR2_X1  g665(.A(KEYINPUT115), .B(KEYINPUT47), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n847), .A2(new_n188), .A3(new_n852), .ZN(new_n855));
  NOR4_X1   g669(.A1(new_n542), .A2(new_n757), .A3(new_n652), .A4(new_n809), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(G140), .ZN(G42));
  AND2_X1   g672(.A1(new_n744), .A2(new_n652), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n768), .A2(new_n809), .A3(new_n548), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n796), .ZN(new_n862));
  NOR4_X1   g676(.A1(new_n784), .A2(new_n651), .A3(new_n786), .A4(new_n548), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n821), .A2(new_n863), .ZN(new_n864));
  OAI221_X1 g678(.A(new_n546), .B1(new_n861), .B2(new_n680), .C1(new_n862), .C2(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n821), .A2(new_n811), .A3(new_n860), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT48), .ZN(new_n867));
  OR2_X1    g681(.A1(new_n866), .A2(KEYINPUT48), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n865), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n767), .A2(new_n440), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n871), .A2(new_n188), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n872), .B1(new_n854), .B2(new_n855), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n864), .A2(new_n809), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n870), .A2(new_n544), .A3(new_n188), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT120), .ZN(new_n878));
  OR2_X1    g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n877), .A2(new_n878), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n879), .A2(new_n734), .A3(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n864), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT50), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n821), .A2(new_n800), .A3(new_n860), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n859), .A2(new_n678), .A3(new_n797), .A4(new_n860), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT121), .ZN(new_n886));
  OR2_X1    g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n885), .A2(new_n886), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n884), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n883), .A2(KEYINPUT51), .A3(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n869), .B1(new_n876), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(KEYINPUT119), .B1(new_n873), .B2(new_n875), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT119), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n847), .A2(new_n188), .A3(new_n852), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n852), .B1(new_n847), .B2(new_n188), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n893), .B(new_n874), .C1(new_n896), .C2(new_n872), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n892), .A2(new_n897), .A3(new_n883), .A4(new_n889), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT51), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n891), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n719), .A2(new_n722), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n801), .B1(new_n901), .B2(new_n725), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n902), .B1(new_n753), .B2(new_n760), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n724), .A2(new_n746), .A3(new_n717), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n744), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(new_n793), .ZN(new_n906));
  AOI21_X1  g720(.A(KEYINPUT52), .B1(new_n903), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n784), .A2(new_n786), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(new_n710), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n909), .A2(new_n757), .ZN(new_n910));
  AOI22_X1  g724(.A1(new_n723), .A2(new_n726), .B1(new_n796), .B2(new_n910), .ZN(new_n911));
  AND4_X1   g725(.A1(KEYINPUT52), .A2(new_n911), .A3(new_n761), .A4(new_n906), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n907), .A2(new_n912), .ZN(new_n913));
  AOI22_X1  g727(.A1(new_n777), .A2(new_n772), .B1(new_n788), .B2(new_n793), .ZN(new_n914));
  AOI22_X1  g728(.A1(new_n772), .A2(new_n773), .B1(new_n780), .B2(new_n759), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n914), .A2(new_n813), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(KEYINPUT117), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT117), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n914), .A2(new_n813), .A3(new_n915), .A4(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(new_n328), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n920), .B1(new_n797), .B2(new_n679), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n921), .A2(new_n655), .A3(new_n611), .A4(new_n657), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n922), .A2(new_n653), .A3(new_n711), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n542), .A2(new_n710), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT116), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n698), .A2(new_n326), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n322), .A2(new_n327), .A3(new_n717), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(new_n927), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n929), .A2(KEYINPUT116), .A3(new_n326), .A4(new_n698), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n924), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n810), .B1(new_n932), .B2(new_n910), .ZN(new_n933));
  AND4_X1   g747(.A1(KEYINPUT53), .A2(new_n818), .A3(new_n923), .A4(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n917), .A2(new_n919), .A3(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n913), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n903), .A2(KEYINPUT52), .A3(new_n906), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n911), .A2(new_n761), .A3(new_n906), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT52), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n818), .A2(new_n923), .A3(new_n933), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n916), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(KEYINPUT53), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n936), .A2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT118), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT54), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n943), .B1(new_n907), .B2(new_n912), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT53), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(KEYINPUT54), .B1(new_n951), .B2(new_n944), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n949), .A2(new_n950), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n941), .A2(new_n919), .A3(new_n917), .A4(new_n934), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n953), .A2(new_n954), .A3(new_n947), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(KEYINPUT118), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n900), .A2(new_n948), .A3(new_n952), .A4(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n545), .A2(new_n420), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT122), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n871), .A2(KEYINPUT49), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n871), .A2(KEYINPUT49), .ZN(new_n962));
  NOR4_X1   g776(.A1(new_n961), .A2(new_n962), .A3(new_n544), .A4(new_n189), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n963), .A2(new_n734), .A3(new_n820), .A4(new_n859), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n960), .A2(new_n964), .ZN(G75));
  NAND2_X1  g779(.A1(new_n953), .A2(new_n954), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n966), .A2(G210), .A3(G902), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT56), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n570), .B1(new_n580), .B2(new_n582), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(new_n574), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT55), .ZN(new_n971));
  AND3_X1   g785(.A1(new_n967), .A2(new_n968), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n971), .B1(new_n967), .B2(new_n968), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n420), .A2(G952), .ZN(new_n974));
  NOR3_X1   g788(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(G51));
  XOR2_X1   g789(.A(new_n828), .B(KEYINPUT57), .Z(new_n976));
  AOI21_X1  g790(.A(new_n947), .B1(new_n953), .B2(new_n954), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT123), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n955), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n978), .B(KEYINPUT54), .C1(new_n936), .C2(new_n944), .ZN(new_n980));
  INV_X1    g794(.A(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n976), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(new_n766), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n966), .A2(G902), .ZN(new_n985));
  OR3_X1    g799(.A1(new_n985), .A2(new_n841), .A3(new_n842), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n974), .B1(new_n984), .B2(new_n986), .ZN(G54));
  NAND2_X1  g801(.A1(KEYINPUT58), .A2(G475), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n260), .B1(new_n985), .B2(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(new_n974), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NOR3_X1   g805(.A1(new_n985), .A2(new_n260), .A3(new_n988), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n991), .A2(new_n992), .ZN(G60));
  NAND2_X1  g807(.A1(G478), .A2(G902), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n994), .B(KEYINPUT59), .ZN(new_n995));
  OAI211_X1 g809(.A(new_n673), .B(new_n995), .C1(new_n979), .C2(new_n981), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(new_n990), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n948), .A2(new_n952), .A3(new_n956), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n673), .B1(new_n998), .B2(new_n995), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n997), .A2(new_n999), .ZN(G63));
  NAND2_X1  g814(.A1(G217), .A2(G902), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1001), .B(KEYINPUT60), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n966), .A2(new_n708), .A3(new_n1003), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n945), .A2(new_n1002), .ZN(new_n1005));
  OAI211_X1 g819(.A(new_n990), .B(new_n1004), .C1(new_n1005), .C2(new_n644), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT61), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1006), .B(new_n1007), .ZN(G66));
  NAND3_X1  g822(.A1(new_n550), .A2(G224), .A3(G953), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n914), .A2(new_n915), .A3(new_n923), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1009), .B1(new_n1010), .B2(G953), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n969), .B1(G898), .B2(new_n420), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1011), .B(new_n1012), .Z(G69));
  INV_X1    g827(.A(KEYINPUT125), .ZN(new_n1014));
  AND2_X1   g828(.A1(new_n793), .A2(new_n811), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n847), .A2(new_n188), .A3(new_n730), .A4(new_n1015), .ZN(new_n1016));
  AND4_X1   g830(.A1(new_n813), .A2(new_n1016), .A3(new_n818), .A4(new_n903), .ZN(new_n1017));
  INV_X1    g831(.A(new_n849), .ZN(new_n1018));
  NAND4_X1  g832(.A1(new_n1017), .A2(new_n1018), .A3(new_n420), .A4(new_n857), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n499), .A2(new_n500), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n502), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n248), .A2(new_n251), .ZN(new_n1022));
  XOR2_X1   g836(.A(new_n1021), .B(new_n1022), .Z(new_n1023));
  AOI21_X1  g837(.A(new_n1023), .B1(G900), .B2(G953), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1019), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n921), .A2(new_n730), .ZN(new_n1026));
  NOR2_X1   g840(.A1(new_n805), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n903), .A2(new_n749), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1027), .B1(new_n1028), .B2(KEYINPUT62), .ZN(new_n1029));
  INV_X1    g843(.A(KEYINPUT62), .ZN(new_n1030));
  NAND3_X1  g844(.A1(new_n903), .A2(new_n1030), .A3(new_n749), .ZN(new_n1031));
  AND2_X1   g845(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n849), .B1(new_n896), .B2(new_n856), .ZN(new_n1033));
  AOI21_X1  g847(.A(G953), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  XOR2_X1   g848(.A(new_n1023), .B(KEYINPUT124), .Z(new_n1035));
  INV_X1    g849(.A(new_n1035), .ZN(new_n1036));
  OAI211_X1 g850(.A(new_n1014), .B(new_n1025), .C1(new_n1034), .C2(new_n1036), .ZN(new_n1037));
  INV_X1    g851(.A(KEYINPUT126), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n420), .B1(G227), .B2(G900), .ZN(new_n1039));
  INV_X1    g853(.A(new_n1039), .ZN(new_n1040));
  NAND3_X1  g854(.A1(new_n1037), .A2(new_n1038), .A3(new_n1040), .ZN(new_n1041));
  NAND4_X1  g855(.A1(new_n1018), .A2(new_n857), .A3(new_n1029), .A4(new_n1031), .ZN(new_n1042));
  NAND2_X1  g856(.A1(new_n1042), .A2(new_n420), .ZN(new_n1043));
  AOI22_X1  g857(.A1(new_n1043), .A2(new_n1035), .B1(new_n1019), .B2(new_n1024), .ZN(new_n1044));
  AOI21_X1  g858(.A(KEYINPUT126), .B1(new_n1044), .B2(new_n1014), .ZN(new_n1045));
  OAI211_X1 g859(.A(KEYINPUT126), .B(new_n1025), .C1(new_n1034), .C2(new_n1036), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n1046), .A2(new_n1039), .ZN(new_n1047));
  OAI21_X1  g861(.A(new_n1041), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g862(.A(new_n1048), .ZN(G72));
  NAND2_X1  g863(.A1(G472), .A2(G902), .ZN(new_n1050));
  XOR2_X1   g864(.A(new_n1050), .B(KEYINPUT63), .Z(new_n1051));
  NAND3_X1  g865(.A1(new_n506), .A2(new_n509), .A3(new_n521), .ZN(new_n1052));
  OAI211_X1 g866(.A(new_n1051), .B(new_n1052), .C1(new_n951), .C2(new_n944), .ZN(new_n1053));
  NAND2_X1  g867(.A1(new_n1053), .A2(new_n990), .ZN(new_n1054));
  INV_X1    g868(.A(new_n1010), .ZN(new_n1055));
  NAND3_X1  g869(.A1(new_n1033), .A2(new_n1055), .A3(new_n1017), .ZN(new_n1056));
  AOI211_X1 g870(.A(new_n488), .B(new_n505), .C1(new_n1056), .C2(new_n1051), .ZN(new_n1057));
  OAI21_X1  g871(.A(new_n1051), .B1(new_n1042), .B2(new_n1010), .ZN(new_n1058));
  INV_X1    g872(.A(KEYINPUT127), .ZN(new_n1059));
  OR2_X1    g873(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g874(.A(new_n738), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1061));
  AOI211_X1 g875(.A(new_n1054), .B(new_n1057), .C1(new_n1060), .C2(new_n1061), .ZN(G57));
endmodule


