//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 1 0 1 0 0 0 1 1 1 0 0 1 1 1 0 1 1 0 1 1 1 0 0 0 1 0 1 0 0 1 0 1 1 0 1 0 0 1 0 1 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:17 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n438, new_n445, new_n450, new_n452, new_n453,
    new_n456, new_n457, new_n458, new_n459, new_n460, new_n461, new_n464,
    new_n465, new_n466, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n536, new_n537, new_n538, new_n539, new_n540, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n555, new_n556, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n628, new_n629, new_n632,
    new_n633, new_n635, new_n636, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n847, new_n848, new_n849, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1189, new_n1190,
    new_n1191;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  OR2_X1    g011(.A1(new_n436), .A2(KEYINPUT66), .ZN(new_n437));
  NAND2_X1  g012(.A1(new_n436), .A2(KEYINPUT66), .ZN(new_n438));
  NAND2_X1  g013(.A1(new_n437), .A2(new_n438), .ZN(G220));
  INV_X1    g014(.A(G96), .ZN(G221));
  INV_X1    g015(.A(G69), .ZN(G235));
  INV_X1    g016(.A(G120), .ZN(G236));
  INV_X1    g017(.A(G57), .ZN(G237));
  INV_X1    g018(.A(G108), .ZN(G238));
  NAND4_X1  g019(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT67), .Z(G158));
  NAND3_X1  g021(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  INV_X1    g026(.A(G567), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT68), .ZN(G234));
  NAND3_X1  g029(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR3_X1   g030(.A1(G219), .A2(G218), .A3(G221), .ZN(new_n456));
  NAND3_X1  g031(.A1(new_n456), .A2(new_n438), .A3(new_n437), .ZN(new_n457));
  XNOR2_X1  g032(.A(KEYINPUT69), .B(KEYINPUT2), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n457), .B(new_n458), .ZN(new_n459));
  NOR4_X1   g034(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n459), .A2(new_n461), .ZN(G325));
  INV_X1    g037(.A(G325), .ZN(G261));
  NAND2_X1  g038(.A1(new_n459), .A2(G2106), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n464), .B1(new_n452), .B2(new_n460), .ZN(new_n465));
  XOR2_X1   g040(.A(new_n465), .B(KEYINPUT70), .Z(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(G319));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  AND2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  OAI21_X1  g045(.A(G125), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n468), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI211_X1 g048(.A(G137), .B(new_n468), .C1(new_n469), .C2(new_n470), .ZN(new_n474));
  INV_X1    g049(.A(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G101), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n473), .A2(new_n478), .ZN(G160));
  OAI21_X1  g054(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(G112), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n480), .B1(new_n481), .B2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT3), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(new_n475), .ZN(new_n484));
  NAND2_X1  g059(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n485));
  AOI21_X1  g060(.A(G2105), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n482), .B1(G136), .B2(new_n486), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n468), .B1(new_n484), .B2(new_n485), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT71), .ZN(new_n489));
  OR2_X1    g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n489), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G124), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n487), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  XNOR2_X1  g069(.A(new_n494), .B(KEYINPUT72), .ZN(G162));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n497), .B1(new_n469), .B2(new_n470), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n484), .A2(new_n485), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n501), .A2(G126), .A3(G2105), .ZN(new_n502));
  OR2_X1    g077(.A1(G102), .A2(G2105), .ZN(new_n503));
  OAI211_X1 g078(.A(new_n503), .B(G2104), .C1(G114), .C2(new_n468), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n497), .B(KEYINPUT4), .C1(new_n470), .C2(new_n469), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n500), .A2(new_n502), .A3(new_n504), .A4(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  XNOR2_X1  g082(.A(KEYINPUT5), .B(G543), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n508), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g086(.A(new_n511), .B(KEYINPUT75), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  OAI21_X1  g088(.A(KEYINPUT73), .B1(new_n510), .B2(KEYINPUT6), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT73), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n515), .A2(new_n516), .A3(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n510), .A2(KEYINPUT6), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n518), .A2(G543), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n518), .A2(new_n508), .A3(new_n519), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT74), .B(G88), .ZN(new_n522));
  OAI22_X1  g097(.A1(new_n513), .A2(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n512), .A2(new_n523), .ZN(G166));
  INV_X1    g099(.A(new_n521), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G89), .ZN(new_n526));
  INV_X1    g101(.A(new_n520), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G51), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n529), .A2(KEYINPUT7), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(KEYINPUT7), .ZN(new_n531));
  AND2_X1   g106(.A1(G63), .A2(G651), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n530), .A2(new_n531), .B1(new_n508), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n526), .A2(new_n528), .A3(new_n533), .ZN(G286));
  INV_X1    g109(.A(G286), .ZN(G168));
  NAND2_X1  g110(.A1(new_n527), .A2(G52), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n537), .A2(new_n510), .ZN(new_n538));
  XNOR2_X1  g113(.A(KEYINPUT76), .B(G90), .ZN(new_n539));
  OAI211_X1 g114(.A(new_n536), .B(new_n538), .C1(new_n521), .C2(new_n539), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT77), .ZN(G171));
  NAND2_X1  g116(.A1(G68), .A2(G543), .ZN(new_n542));
  AND2_X1   g117(.A1(KEYINPUT5), .A2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(KEYINPUT5), .A2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(G56), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n542), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G651), .ZN(new_n548));
  INV_X1    g123(.A(G81), .ZN(new_n549));
  INV_X1    g124(.A(G43), .ZN(new_n550));
  OAI221_X1 g125(.A(new_n548), .B1(new_n521), .B2(new_n549), .C1(new_n550), .C2(new_n520), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  INV_X1    g132(.A(G65), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(KEYINPUT79), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT79), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G65), .ZN(new_n561));
  OAI211_X1 g136(.A(new_n559), .B(new_n561), .C1(new_n543), .C2(new_n544), .ZN(new_n562));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n510), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AND2_X1   g139(.A1(G53), .A2(G543), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n515), .B1(new_n516), .B2(G651), .ZN(new_n566));
  NOR3_X1   g141(.A1(new_n510), .A2(KEYINPUT73), .A3(KEYINPUT6), .ZN(new_n567));
  OAI211_X1 g142(.A(new_n519), .B(new_n565), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(KEYINPUT9), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n514), .A2(new_n517), .B1(KEYINPUT6), .B2(new_n510), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT9), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n570), .A2(new_n571), .A3(new_n565), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n564), .B1(new_n569), .B2(new_n572), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n518), .A2(G91), .A3(new_n508), .A4(new_n519), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT78), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n570), .A2(KEYINPUT78), .A3(G91), .A4(new_n508), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n573), .A2(new_n578), .ZN(G299));
  INV_X1    g154(.A(G171), .ZN(G301));
  OR2_X1    g155(.A1(new_n512), .A2(new_n523), .ZN(G303));
  OAI21_X1  g156(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n582));
  INV_X1    g157(.A(G87), .ZN(new_n583));
  INV_X1    g158(.A(G49), .ZN(new_n584));
  OAI221_X1 g159(.A(new_n582), .B1(new_n521), .B2(new_n583), .C1(new_n584), .C2(new_n520), .ZN(G288));
  INV_X1    g160(.A(KEYINPUT80), .ZN(new_n586));
  INV_X1    g161(.A(G61), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n545), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n508), .A2(KEYINPUT80), .A3(G61), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(G651), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT81), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI211_X1 g170(.A(KEYINPUT81), .B(G651), .C1(new_n590), .C2(new_n592), .ZN(new_n596));
  AND2_X1   g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(G48), .ZN(new_n598));
  INV_X1    g173(.A(G86), .ZN(new_n599));
  OAI22_X1  g174(.A1(new_n598), .A2(new_n520), .B1(new_n521), .B2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n597), .A2(new_n601), .ZN(G305));
  AOI22_X1  g177(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n603), .A2(new_n510), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT82), .ZN(new_n605));
  AOI22_X1  g180(.A1(G47), .A2(new_n527), .B1(new_n525), .B2(G85), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(G290));
  INV_X1    g182(.A(KEYINPUT10), .ZN(new_n608));
  INV_X1    g183(.A(G92), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n521), .B2(new_n609), .ZN(new_n610));
  NAND4_X1  g185(.A1(new_n570), .A2(KEYINPUT10), .A3(G92), .A4(new_n508), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(G79), .A2(G543), .ZN(new_n613));
  INV_X1    g188(.A(G66), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n545), .B2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT84), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  OAI211_X1 g192(.A(KEYINPUT84), .B(new_n613), .C1(new_n545), .C2(new_n614), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n617), .A2(G651), .A3(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT83), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n520), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n570), .A2(KEYINPUT83), .A3(G543), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n621), .A2(G54), .A3(new_n622), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n612), .A2(new_n619), .A3(new_n623), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n624), .A2(G868), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n625), .B1(G171), .B2(G868), .ZN(G284));
  XNOR2_X1  g201(.A(G284), .B(KEYINPUT85), .ZN(G321));
  INV_X1    g202(.A(G868), .ZN(new_n628));
  NAND2_X1  g203(.A1(G299), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(G168), .B2(new_n628), .ZN(G297));
  OAI21_X1  g205(.A(new_n629), .B1(G168), .B2(new_n628), .ZN(G280));
  AND3_X1   g206(.A1(new_n612), .A2(new_n619), .A3(new_n623), .ZN(new_n632));
  INV_X1    g207(.A(G559), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n632), .B1(new_n633), .B2(G860), .ZN(G148));
  NAND2_X1  g209(.A1(new_n551), .A2(new_n628), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n624), .A2(G559), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n635), .B1(new_n636), .B2(new_n628), .ZN(G323));
  XNOR2_X1  g212(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g213(.A1(new_n501), .A2(new_n476), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT86), .B(KEYINPUT12), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT13), .Z(new_n642));
  NOR2_X1   g217(.A1(new_n642), .A2(G2100), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT87), .ZN(new_n644));
  INV_X1    g219(.A(new_n492), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n645), .A2(G123), .ZN(new_n646));
  OAI21_X1  g221(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n647), .A2(KEYINPUT88), .ZN(new_n648));
  INV_X1    g223(.A(G111), .ZN(new_n649));
  AOI22_X1  g224(.A1(new_n647), .A2(KEYINPUT88), .B1(new_n649), .B2(G2105), .ZN(new_n650));
  AOI22_X1  g225(.A1(new_n648), .A2(new_n650), .B1(new_n486), .B2(G135), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n646), .A2(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(G2096), .ZN(new_n654));
  AOI22_X1  g229(.A1(G2100), .A2(new_n642), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  OAI211_X1 g230(.A(new_n644), .B(new_n655), .C1(new_n654), .C2(new_n653), .ZN(G156));
  XNOR2_X1  g231(.A(G2427), .B(G2438), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2430), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT15), .B(G2435), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n660), .A2(KEYINPUT14), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2451), .B(G2454), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT16), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n662), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2443), .B(G2446), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1341), .B(G1348), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(KEYINPUT89), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  OAI21_X1  g246(.A(G14), .B1(new_n667), .B2(new_n668), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(G401));
  XOR2_X1   g248(.A(G2072), .B(G2078), .Z(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2067), .B(G2678), .ZN(new_n676));
  XOR2_X1   g251(.A(G2084), .B(G2090), .Z(new_n677));
  NAND3_X1  g252(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT18), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT90), .B(KEYINPUT17), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n674), .B(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n677), .ZN(new_n682));
  NOR3_X1   g257(.A1(new_n681), .A2(new_n676), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n682), .B1(new_n675), .B2(new_n676), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(new_n681), .B2(new_n676), .ZN(new_n685));
  NOR3_X1   g260(.A1(new_n679), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G2096), .B(G2100), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(G227));
  XNOR2_X1  g263(.A(G1971), .B(G1976), .ZN(new_n689));
  INV_X1    g264(.A(KEYINPUT19), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(G1956), .B(G2474), .Z(new_n692));
  XOR2_X1   g267(.A(G1961), .B(G1966), .Z(new_n693));
  AND2_X1   g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT20), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n692), .A2(new_n693), .ZN(new_n697));
  NOR3_X1   g272(.A1(new_n691), .A2(new_n694), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(new_n691), .B2(new_n697), .ZN(new_n699));
  AND2_X1   g274(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(G1991), .B(G1996), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1981), .B(G1986), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n702), .A2(new_n703), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n702), .A2(new_n703), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n705), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n707), .A2(new_n710), .ZN(G229));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G26), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT28), .Z(new_n714));
  NAND2_X1  g289(.A1(new_n486), .A2(G140), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n468), .A2(G116), .ZN(new_n716));
  OAI21_X1  g291(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n717));
  INV_X1    g292(.A(G128), .ZN(new_n718));
  OAI221_X1 g293(.A(new_n715), .B1(new_n716), .B2(new_n717), .C1(new_n492), .C2(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n714), .B1(new_n719), .B2(G29), .ZN(new_n720));
  INV_X1    g295(.A(G2067), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n551), .A2(G16), .ZN(new_n723));
  INV_X1    g298(.A(G16), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G19), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n722), .B1(G1341), .B2(new_n727), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n712), .A2(G32), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n468), .A2(G105), .A3(G2104), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT95), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  AND3_X1   g307(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT26), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n486), .A2(G141), .ZN(new_n735));
  AND3_X1   g310(.A1(new_n732), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(G129), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n736), .B1(new_n492), .B2(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT96), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n738), .A2(new_n739), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n729), .B1(new_n742), .B2(G29), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT27), .B(G1996), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT31), .B(G11), .ZN(new_n746));
  INV_X1    g321(.A(G28), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n747), .A2(KEYINPUT30), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT30), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n712), .B1(new_n749), .B2(G28), .ZN(new_n750));
  OAI221_X1 g325(.A(new_n746), .B1(new_n748), .B2(new_n750), .C1(new_n652), .C2(new_n712), .ZN(new_n751));
  NOR2_X1   g326(.A1(G27), .A2(G29), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G164), .B2(G29), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT99), .B(G2078), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n751), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n753), .A2(new_n754), .ZN(new_n756));
  NAND2_X1  g331(.A1(G160), .A2(G29), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT24), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n758), .A2(G34), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n712), .B1(new_n758), .B2(G34), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n757), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(G2084), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(G2072), .ZN(new_n764));
  OR2_X1    g339(.A1(G29), .A2(G33), .ZN(new_n765));
  XOR2_X1   g340(.A(KEYINPUT93), .B(KEYINPUT25), .Z(new_n766));
  NAND3_X1  g341(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n486), .A2(G139), .ZN(new_n769));
  AOI22_X1  g344(.A1(new_n501), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n768), .B(new_n769), .C1(new_n468), .C2(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n765), .B1(new_n771), .B2(new_n712), .ZN(new_n772));
  AOI211_X1 g347(.A(new_n756), .B(new_n763), .C1(new_n764), .C2(new_n772), .ZN(new_n773));
  NAND4_X1  g348(.A1(new_n728), .A2(new_n745), .A3(new_n755), .A4(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n724), .A2(G20), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT23), .Z(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G299), .B2(G16), .ZN(new_n777));
  INV_X1    g352(.A(G1956), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n772), .A2(new_n764), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT94), .ZN(new_n781));
  INV_X1    g356(.A(G1341), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n724), .A2(G21), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G168), .B2(new_n724), .ZN(new_n784));
  XOR2_X1   g359(.A(KEYINPUT97), .B(G1966), .Z(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  AOI22_X1  g361(.A1(new_n782), .A2(new_n726), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n781), .B(new_n787), .C1(new_n784), .C2(new_n786), .ZN(new_n788));
  NOR3_X1   g363(.A1(new_n774), .A2(new_n779), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n761), .A2(new_n762), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n724), .A2(G5), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G171), .B2(new_n724), .ZN(new_n792));
  OAI221_X1 g367(.A(new_n790), .B1(new_n792), .B2(G1961), .C1(new_n743), .C2(new_n744), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT98), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(G4), .A2(G16), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(new_n632), .B2(G16), .ZN(new_n797));
  AND2_X1   g372(.A1(new_n797), .A2(G1348), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n792), .B2(G1961), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G1348), .B2(new_n797), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n795), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(G29), .A2(G35), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G162), .B2(G29), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT29), .ZN(new_n804));
  INV_X1    g379(.A(G2090), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n793), .A2(new_n794), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n789), .A2(new_n801), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n724), .A2(G23), .ZN(new_n809));
  INV_X1    g384(.A(G288), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n809), .B1(new_n810), .B2(new_n724), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT33), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G1976), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n724), .A2(G6), .ZN(new_n814));
  INV_X1    g389(.A(G305), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n814), .B1(new_n815), .B2(new_n724), .ZN(new_n816));
  XNOR2_X1  g391(.A(KEYINPUT32), .B(G1981), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n816), .A2(new_n817), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n724), .A2(G22), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT92), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(G166), .B2(new_n724), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(G1971), .Z(new_n823));
  NAND4_X1  g398(.A1(new_n813), .A2(new_n818), .A3(new_n819), .A4(new_n823), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n824), .A2(KEYINPUT34), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(KEYINPUT34), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n712), .A2(G25), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n645), .A2(G119), .ZN(new_n828));
  NOR2_X1   g403(.A1(G95), .A2(G2105), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(KEYINPUT91), .Z(new_n830));
  INV_X1    g405(.A(G107), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n475), .B1(new_n831), .B2(G2105), .ZN(new_n832));
  AOI22_X1  g407(.A1(new_n830), .A2(new_n832), .B1(G131), .B2(new_n486), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n828), .A2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n827), .B1(new_n835), .B2(new_n712), .ZN(new_n836));
  XOR2_X1   g411(.A(KEYINPUT35), .B(G1991), .Z(new_n837));
  XOR2_X1   g412(.A(new_n836), .B(new_n837), .Z(new_n838));
  MUX2_X1   g413(.A(G24), .B(G290), .S(G16), .Z(new_n839));
  NOR2_X1   g414(.A1(new_n839), .A2(G1986), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n839), .A2(G1986), .ZN(new_n841));
  NOR3_X1   g416(.A1(new_n838), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n825), .A2(new_n826), .A3(new_n842), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n843), .A2(KEYINPUT36), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(KEYINPUT36), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n808), .B1(new_n844), .B2(new_n845), .ZN(G311));
  INV_X1    g421(.A(new_n808), .ZN(new_n847));
  INV_X1    g422(.A(new_n845), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n843), .A2(KEYINPUT36), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n847), .B1(new_n848), .B2(new_n849), .ZN(G150));
  INV_X1    g425(.A(G860), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT39), .ZN(new_n852));
  AOI22_X1  g427(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n853), .A2(new_n510), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n518), .A2(G55), .A3(G543), .A4(new_n519), .ZN(new_n855));
  NAND4_X1  g430(.A1(new_n518), .A2(G93), .A3(new_n508), .A4(new_n519), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT100), .ZN(new_n857));
  AND3_X1   g432(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n857), .B1(new_n855), .B2(new_n856), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n854), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(KEYINPUT101), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT101), .ZN(new_n862));
  OAI211_X1 g437(.A(new_n862), .B(new_n854), .C1(new_n858), .C2(new_n859), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n861), .A2(new_n551), .A3(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n860), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n865), .A2(new_n862), .A3(new_n552), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT38), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n632), .A2(G559), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n868), .B(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(new_n852), .ZN(new_n871));
  AND2_X1   g446(.A1(new_n871), .A2(KEYINPUT102), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n871), .A2(KEYINPUT102), .ZN(new_n873));
  OAI221_X1 g448(.A(new_n851), .B1(new_n852), .B2(new_n870), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n860), .A2(G860), .ZN(new_n875));
  XOR2_X1   g450(.A(new_n875), .B(KEYINPUT37), .Z(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(G145));
  NAND2_X1  g452(.A1(new_n486), .A2(G142), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n468), .A2(G118), .ZN(new_n879));
  OAI21_X1  g454(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n881), .B1(new_n645), .B2(G130), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n834), .B(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n771), .A2(KEYINPUT104), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(G164), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n883), .B(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n742), .B(new_n719), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(new_n641), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n888), .A2(new_n641), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n887), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n891), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n893), .A2(new_n886), .A3(new_n889), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(G162), .B(G160), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(KEYINPUT103), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(new_n653), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT103), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n896), .B(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(new_n652), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n895), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(G37), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n898), .A2(new_n892), .A3(new_n894), .A4(new_n901), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g482(.A1(new_n815), .A2(G288), .ZN(new_n908));
  XNOR2_X1  g483(.A(G166), .B(G290), .ZN(new_n909));
  NOR2_X1   g484(.A1(G305), .A2(new_n810), .ZN(new_n910));
  NOR3_X1   g485(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n909), .B1(new_n908), .B2(new_n910), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(KEYINPUT107), .A2(KEYINPUT42), .ZN(new_n915));
  OR2_X1    g490(.A1(KEYINPUT107), .A2(KEYINPUT42), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n912), .A2(new_n913), .A3(KEYINPUT107), .A4(KEYINPUT42), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(G299), .A2(KEYINPUT105), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT105), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n573), .A2(new_n578), .A3(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n920), .A2(new_n632), .A3(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n624), .A2(KEYINPUT105), .A3(G299), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT106), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT41), .ZN(new_n927));
  AOI211_X1 g502(.A(new_n926), .B(new_n927), .C1(new_n923), .C2(new_n924), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n923), .A2(new_n927), .A3(new_n924), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n927), .B1(new_n923), .B2(new_n924), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n928), .B1(new_n931), .B2(new_n926), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n867), .B(new_n636), .ZN(new_n933));
  MUX2_X1   g508(.A(new_n925), .B(new_n932), .S(new_n933), .Z(new_n934));
  AND2_X1   g509(.A1(new_n919), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n919), .A2(new_n934), .ZN(new_n936));
  OAI21_X1  g511(.A(G868), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n937), .B1(G868), .B2(new_n865), .ZN(G295));
  OAI21_X1  g513(.A(new_n937), .B1(G868), .B2(new_n865), .ZN(G331));
  AND3_X1   g514(.A1(G171), .A2(new_n864), .A3(new_n866), .ZN(new_n940));
  AOI21_X1  g515(.A(G171), .B1(new_n864), .B2(new_n866), .ZN(new_n941));
  OAI21_X1  g516(.A(G286), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n867), .A2(G301), .ZN(new_n943));
  NAND3_X1  g518(.A1(G171), .A2(new_n864), .A3(new_n866), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n943), .A2(G168), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(new_n932), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n942), .A2(new_n945), .A3(new_n925), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n913), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n950), .A2(new_n911), .ZN(new_n951));
  AOI21_X1  g526(.A(G37), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n947), .A2(new_n914), .A3(new_n948), .ZN(new_n953));
  AOI21_X1  g528(.A(KEYINPUT43), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n948), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n931), .B1(new_n942), .B2(new_n945), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n951), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  AND4_X1   g532(.A1(KEYINPUT43), .A2(new_n957), .A3(new_n953), .A4(new_n904), .ZN(new_n958));
  OAI21_X1  g533(.A(KEYINPUT44), .B1(new_n954), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT44), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT43), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n961), .B1(new_n952), .B2(new_n953), .ZN(new_n962));
  AND4_X1   g537(.A1(new_n961), .A2(new_n957), .A3(new_n953), .A4(new_n904), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n960), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n959), .A2(new_n964), .ZN(G397));
  INV_X1    g540(.A(KEYINPUT109), .ZN(new_n966));
  INV_X1    g541(.A(G1384), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n506), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT45), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(G125), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n971), .B1(new_n484), .B2(new_n485), .ZN(new_n972));
  INV_X1    g547(.A(new_n472), .ZN(new_n973));
  OAI21_X1  g548(.A(G2105), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  XOR2_X1   g549(.A(KEYINPUT108), .B(G40), .Z(new_n975));
  NAND4_X1  g550(.A1(new_n974), .A2(new_n477), .A3(new_n474), .A4(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n966), .B1(new_n970), .B2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(KEYINPUT45), .B1(new_n506), .B2(new_n967), .ZN(new_n978));
  INV_X1    g553(.A(new_n976), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n978), .A2(new_n979), .A3(KEYINPUT109), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G1996), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OR3_X1    g559(.A1(new_n984), .A2(KEYINPUT110), .A3(new_n742), .ZN(new_n985));
  OAI21_X1  g560(.A(KEYINPUT110), .B1(new_n984), .B2(new_n742), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n983), .B1(new_n740), .B2(new_n741), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n719), .B(G2067), .ZN(new_n988));
  OR2_X1    g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  AOI22_X1  g564(.A1(new_n985), .A2(new_n986), .B1(new_n982), .B2(new_n989), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n834), .B(new_n837), .ZN(new_n991));
  OR2_X1    g566(.A1(new_n991), .A2(new_n981), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g568(.A(G290), .B(G1986), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n993), .B1(new_n982), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT53), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n506), .A2(KEYINPUT45), .A3(new_n967), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n970), .A2(new_n979), .A3(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n996), .B1(new_n998), .B2(G2078), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n968), .A2(KEYINPUT50), .ZN(new_n1000));
  XOR2_X1   g575(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n1000), .B(new_n979), .C1(new_n968), .C2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G1961), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AND2_X1   g580(.A1(new_n999), .A2(new_n1005), .ZN(new_n1006));
  AND3_X1   g581(.A1(new_n506), .A2(KEYINPUT45), .A3(new_n967), .ZN(new_n1007));
  NOR3_X1   g582(.A1(new_n1007), .A2(new_n978), .A3(new_n976), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n996), .A2(G2078), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1006), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(G171), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1007), .A2(new_n978), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1013), .A2(G40), .A3(G160), .A4(new_n1009), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n999), .A2(new_n1005), .A3(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1012), .B1(G171), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT124), .ZN(new_n1019));
  AOI21_X1  g594(.A(G301), .B1(new_n1015), .B2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1020), .B1(new_n1019), .B2(new_n1015), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n1021), .B(KEYINPUT54), .C1(G171), .C2(new_n1011), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT115), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n600), .B(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n597), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(G1981), .ZN(new_n1026));
  XNOR2_X1  g601(.A(KEYINPUT114), .B(G1981), .ZN(new_n1027));
  AND4_X1   g602(.A1(new_n596), .A2(new_n595), .A3(new_n601), .A4(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1026), .A2(new_n1029), .A3(KEYINPUT49), .ZN(new_n1030));
  NAND4_X1  g605(.A1(G160), .A2(new_n506), .A3(new_n967), .A4(new_n975), .ZN(new_n1031));
  XOR2_X1   g606(.A(KEYINPUT113), .B(G8), .Z(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT49), .ZN(new_n1036));
  INV_X1    g611(.A(G1981), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1037), .B1(new_n597), .B2(new_n1024), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1036), .B1(new_n1038), .B2(new_n1028), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1030), .A2(new_n1035), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(G1976), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1035), .B1(new_n1041), .B2(G288), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT52), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT52), .B1(G288), .B2(new_n1041), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1044), .B1(new_n1042), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1040), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n1049));
  INV_X1    g624(.A(G8), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1049), .B1(G166), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1048), .A2(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g627(.A(KEYINPUT111), .B(G1971), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n998), .A2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1054), .B1(new_n1003), .B2(G2090), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1052), .A2(G8), .A3(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n976), .B1(new_n968), .B2(new_n1002), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT50), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n506), .A2(new_n1058), .A3(new_n967), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1057), .A2(new_n805), .A3(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1032), .B1(new_n1054), .B2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1056), .B1(new_n1052), .B2(new_n1061), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1047), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT51), .ZN(new_n1064));
  XOR2_X1   g639(.A(KEYINPUT116), .B(G2084), .Z(new_n1065));
  OAI22_X1  g640(.A1(new_n1003), .A2(new_n1065), .B1(new_n1008), .B2(new_n786), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(G8), .ZN(new_n1067));
  NAND2_X1  g642(.A1(G286), .A2(new_n1033), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1064), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1066), .A2(G286), .A3(new_n1033), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1066), .A2(new_n1033), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT51), .B1(G286), .B2(new_n1033), .ZN(new_n1072));
  AOI22_X1  g647(.A1(new_n1069), .A2(new_n1070), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1018), .A2(new_n1022), .A3(new_n1063), .A4(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT61), .ZN(new_n1075));
  NOR2_X1   g650(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n1076));
  XOR2_X1   g651(.A(new_n1076), .B(KEYINPUT118), .Z(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT117), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT57), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1078), .B1(G299), .B2(new_n1082), .ZN(new_n1083));
  AOI211_X1 g658(.A(new_n1081), .B(new_n1077), .C1(new_n573), .C2(new_n578), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(G1956), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1086));
  XOR2_X1   g661(.A(KEYINPUT56), .B(G2072), .Z(new_n1087));
  NOR4_X1   g662(.A1(new_n1007), .A2(new_n978), .A3(new_n976), .A4(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1086), .B1(new_n1088), .B2(KEYINPUT119), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1090), .B1(new_n998), .B2(new_n1087), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1085), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n778), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1087), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1013), .A2(KEYINPUT119), .A3(new_n979), .A4(new_n1095), .ZN(new_n1096));
  AND4_X1   g671(.A1(new_n1085), .A2(new_n1091), .A3(new_n1094), .A4(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1075), .B1(new_n1092), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT59), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n970), .A2(new_n983), .A3(new_n979), .A4(new_n997), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT121), .ZN(new_n1101));
  XOR2_X1   g676(.A(KEYINPUT58), .B(G1341), .Z(new_n1102));
  AND3_X1   g677(.A1(new_n1031), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1101), .B1(new_n1031), .B2(new_n1102), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1100), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT122), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  OAI211_X1 g682(.A(KEYINPUT122), .B(new_n1100), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1099), .B1(new_n1109), .B2(new_n552), .ZN(new_n1110));
  AOI211_X1 g685(.A(KEYINPUT59), .B(new_n551), .C1(new_n1107), .C2(new_n1108), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1098), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1089), .A2(new_n1085), .A3(new_n1091), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(KEYINPUT61), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT120), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1089), .A2(new_n1115), .A3(new_n1091), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1091), .A2(new_n1094), .A3(new_n1096), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1085), .B1(new_n1117), .B2(KEYINPUT120), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1114), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(KEYINPUT123), .B1(new_n1112), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1118), .A2(new_n1116), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1121), .A2(KEYINPUT61), .A3(new_n1113), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1031), .A2(new_n1102), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(KEYINPUT121), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1031), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT122), .B1(new_n1126), .B2(new_n1100), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1108), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n552), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(KEYINPUT59), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1109), .A2(new_n1099), .A3(new_n552), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT123), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1122), .A2(new_n1132), .A3(new_n1133), .A4(new_n1098), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1031), .A2(G2067), .ZN(new_n1135));
  INV_X1    g710(.A(G1348), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1135), .B1(new_n1003), .B2(new_n1136), .ZN(new_n1137));
  AND3_X1   g712(.A1(new_n1137), .A2(KEYINPUT60), .A3(new_n624), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n624), .B1(new_n1137), .B2(KEYINPUT60), .ZN(new_n1139));
  OAI22_X1  g714(.A1(new_n1138), .A2(new_n1139), .B1(KEYINPUT60), .B2(new_n1137), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1120), .A2(new_n1134), .A3(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1121), .B1(new_n624), .B2(new_n1137), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(new_n1113), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1074), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT63), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1047), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1052), .B1(G8), .B2(new_n1055), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1066), .A2(G168), .A3(new_n1033), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1145), .B1(new_n1146), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1148), .ZN(new_n1151));
  OAI211_X1 g726(.A(new_n1151), .B(new_n1145), .C1(new_n1052), .C2(new_n1061), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1047), .B1(new_n1152), .B2(new_n1056), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1040), .A2(new_n1041), .A3(new_n810), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1034), .B1(new_n1154), .B2(new_n1029), .ZN(new_n1155));
  NOR3_X1   g730(.A1(new_n1150), .A2(new_n1153), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT62), .ZN(new_n1160));
  OAI21_X1  g735(.A(KEYINPUT125), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT125), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1073), .A2(new_n1162), .A3(KEYINPUT62), .ZN(new_n1163));
  NOR3_X1   g738(.A1(new_n1047), .A2(new_n1062), .A3(new_n1012), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1161), .A2(new_n1163), .A3(new_n1164), .A4(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1156), .A2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n995), .B1(new_n1144), .B2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n719), .A2(G2067), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n835), .A2(new_n837), .ZN(new_n1170));
  XOR2_X1   g745(.A(new_n1170), .B(KEYINPUT126), .Z(new_n1171));
  AOI21_X1  g746(.A(new_n1169), .B1(new_n990), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT127), .ZN(new_n1173));
  OR3_X1    g748(.A1(new_n1172), .A2(new_n1173), .A3(new_n981), .ZN(new_n1174));
  INV_X1    g749(.A(new_n993), .ZN(new_n1175));
  NOR3_X1   g750(.A1(new_n981), .A2(G1986), .A3(G290), .ZN(new_n1176));
  XOR2_X1   g751(.A(new_n1176), .B(KEYINPUT48), .Z(new_n1177));
  OAI21_X1  g752(.A(new_n982), .B1(new_n988), .B2(new_n742), .ZN(new_n1178));
  AND2_X1   g753(.A1(new_n984), .A2(KEYINPUT46), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n984), .A2(KEYINPUT46), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1178), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1181), .A2(KEYINPUT47), .ZN(new_n1182));
  OR2_X1    g757(.A1(new_n1181), .A2(KEYINPUT47), .ZN(new_n1183));
  AOI22_X1  g758(.A1(new_n1175), .A2(new_n1177), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1173), .B1(new_n1172), .B2(new_n981), .ZN(new_n1185));
  AND3_X1   g760(.A1(new_n1174), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1168), .A2(new_n1186), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g762(.A1(new_n466), .A2(G227), .ZN(new_n1189));
  OAI21_X1  g763(.A(new_n1189), .B1(new_n707), .B2(new_n710), .ZN(new_n1190));
  NOR2_X1   g764(.A1(new_n1190), .A2(G401), .ZN(new_n1191));
  OAI211_X1 g765(.A(new_n906), .B(new_n1191), .C1(new_n962), .C2(new_n963), .ZN(G225));
  INV_X1    g766(.A(G225), .ZN(G308));
endmodule


