//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 1 0 0 0 1 1 1 1 0 0 0 1 0 0 0 1 1 1 1 0 1 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 1 0 0 1 0 1 0 0 0 1 0 0 1 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:36 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n565, new_n566, new_n567, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n618,
    new_n620, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1152, new_n1153, new_n1154;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT66), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(KEYINPUT68), .B(KEYINPUT2), .Z(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(KEYINPUT70), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n463), .B1(new_n464), .B2(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n467), .A2(KEYINPUT70), .A3(G2104), .ZN(new_n468));
  AND3_X1   g043(.A1(new_n465), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n469), .A2(KEYINPUT71), .A3(G137), .A4(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT71), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n465), .A2(new_n468), .A3(new_n470), .A4(new_n466), .ZN(new_n473));
  INV_X1    g048(.A(G137), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n464), .A2(G2105), .ZN(new_n476));
  AOI22_X1  g051(.A1(new_n471), .A2(new_n475), .B1(G101), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  XNOR2_X1  g053(.A(KEYINPUT3), .B(G2104), .ZN(new_n479));
  AOI21_X1  g054(.A(KEYINPUT69), .B1(new_n479), .B2(G125), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n467), .A2(G2104), .ZN(new_n481));
  AND4_X1   g056(.A1(KEYINPUT69), .A2(new_n466), .A3(new_n481), .A4(G125), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n478), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n477), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G160));
  NAND2_X1  g061(.A1(new_n469), .A2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G124), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n470), .A2(G112), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n490));
  OAI22_X1  g065(.A1(new_n487), .A2(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n473), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n491), .B1(G136), .B2(new_n492), .ZN(new_n493));
  XOR2_X1   g068(.A(new_n493), .B(KEYINPUT72), .Z(G162));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n465), .A2(new_n468), .A3(new_n496), .A4(new_n466), .ZN(new_n497));
  NOR3_X1   g072(.A1(new_n495), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n498));
  AOI22_X1  g073(.A1(new_n497), .A2(KEYINPUT4), .B1(new_n479), .B2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT74), .ZN(new_n500));
  AND2_X1   g075(.A1(G126), .A2(G2105), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n465), .A2(new_n468), .A3(new_n466), .A4(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  OAI21_X1  g078(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT73), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n505), .B1(new_n470), .B2(G114), .ZN(new_n506));
  INV_X1    g081(.A(G114), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(KEYINPUT73), .A3(G2105), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n504), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n500), .B1(new_n503), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n504), .ZN(new_n511));
  AND3_X1   g086(.A1(new_n507), .A2(KEYINPUT73), .A3(G2105), .ZN(new_n512));
  AOI21_X1  g087(.A(KEYINPUT73), .B1(new_n507), .B2(G2105), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n514), .A2(KEYINPUT74), .A3(new_n502), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n499), .B1(new_n510), .B2(new_n515), .ZN(G164));
  AND2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G543), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G50), .ZN(new_n522));
  INV_X1    g097(.A(G88), .ZN(new_n523));
  INV_X1    g098(.A(new_n519), .ZN(new_n524));
  NAND2_X1  g099(.A1(KEYINPUT75), .A2(KEYINPUT5), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(new_n520), .ZN(new_n526));
  NAND3_X1  g101(.A1(KEYINPUT75), .A2(KEYINPUT5), .A3(G543), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n524), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n522), .B1(new_n523), .B2(new_n529), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n528), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n531));
  INV_X1    g106(.A(G651), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n530), .A2(new_n533), .ZN(G166));
  INV_X1    g109(.A(new_n527), .ZN(new_n535));
  AOI21_X1  g110(.A(G543), .B1(KEYINPUT75), .B2(KEYINPUT5), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(KEYINPUT76), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT76), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n528), .A2(new_n539), .ZN(new_n540));
  AND2_X1   g115(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  AND3_X1   g116(.A1(new_n541), .A2(G63), .A3(G651), .ZN(new_n542));
  NAND3_X1  g117(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n543));
  XOR2_X1   g118(.A(new_n543), .B(KEYINPUT7), .Z(new_n544));
  AOI21_X1  g119(.A(new_n544), .B1(G51), .B2(new_n521), .ZN(new_n545));
  INV_X1    g120(.A(G89), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n546), .B2(new_n529), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n542), .A2(new_n547), .ZN(G168));
  NAND2_X1  g123(.A1(new_n541), .A2(G64), .ZN(new_n549));
  NAND2_X1  g124(.A1(G77), .A2(G543), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n532), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n521), .A2(G52), .ZN(new_n552));
  INV_X1    g127(.A(G90), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n553), .B2(new_n529), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n551), .A2(new_n554), .ZN(G171));
  NAND2_X1  g130(.A1(new_n541), .A2(G56), .ZN(new_n556));
  NAND2_X1  g131(.A1(G68), .A2(G543), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n532), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n521), .A2(G43), .ZN(new_n559));
  INV_X1    g134(.A(G81), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n560), .B2(new_n529), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  NAND4_X1  g138(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT77), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  AOI22_X1  g143(.A1(new_n528), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n569), .A2(new_n532), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n537), .A2(new_n519), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n570), .B1(G91), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n521), .A2(G53), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT9), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n572), .A2(new_n574), .ZN(G299));
  OR2_X1    g150(.A1(new_n551), .A2(new_n554), .ZN(G301));
  OR2_X1    g151(.A1(new_n542), .A2(new_n547), .ZN(G286));
  INV_X1    g152(.A(G166), .ZN(G303));
  AOI22_X1  g153(.A1(new_n571), .A2(G87), .B1(G49), .B2(new_n521), .ZN(new_n579));
  AOI21_X1  g154(.A(G74), .B1(new_n538), .B2(new_n540), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n580), .B2(new_n532), .ZN(G288));
  INV_X1    g156(.A(G61), .ZN(new_n582));
  NOR3_X1   g157(.A1(new_n537), .A2(KEYINPUT78), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n582), .B1(new_n526), .B2(new_n527), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT78), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n583), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n571), .A2(G86), .B1(G48), .B2(new_n521), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(G305));
  NAND2_X1  g165(.A1(G72), .A2(G543), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n538), .A2(new_n540), .ZN(new_n592));
  INV_X1    g167(.A(G60), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(G651), .ZN(new_n595));
  XOR2_X1   g170(.A(KEYINPUT79), .B(G85), .Z(new_n596));
  AOI22_X1  g171(.A1(new_n571), .A2(new_n596), .B1(new_n521), .B2(G47), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n595), .A2(new_n597), .ZN(G290));
  INV_X1    g173(.A(G868), .ZN(new_n599));
  OR3_X1    g174(.A1(G171), .A2(KEYINPUT80), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(KEYINPUT80), .B1(G171), .B2(new_n599), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n571), .A2(G92), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n602), .B(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(G79), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n537), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n607), .A2(G651), .B1(new_n521), .B2(G54), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT81), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n609), .B(new_n610), .ZN(new_n611));
  OAI211_X1 g186(.A(new_n600), .B(new_n601), .C1(new_n611), .C2(G868), .ZN(G284));
  OAI211_X1 g187(.A(new_n600), .B(new_n601), .C1(new_n611), .C2(G868), .ZN(G321));
  NOR2_X1   g188(.A1(G286), .A2(new_n599), .ZN(new_n614));
  XNOR2_X1  g189(.A(G299), .B(KEYINPUT82), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(new_n599), .ZN(G297));
  XOR2_X1   g191(.A(G297), .B(KEYINPUT83), .Z(G280));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n611), .B1(new_n618), .B2(G860), .ZN(G148));
  INV_X1    g194(.A(new_n562), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(new_n599), .ZN(new_n621));
  AND2_X1   g196(.A1(new_n611), .A2(new_n618), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(new_n599), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g199(.A1(new_n479), .A2(new_n476), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT12), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT13), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2100), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n492), .A2(G135), .ZN(new_n629));
  NOR3_X1   g204(.A1(new_n470), .A2(KEYINPUT84), .A3(G111), .ZN(new_n630));
  OAI21_X1  g205(.A(KEYINPUT84), .B1(new_n470), .B2(G111), .ZN(new_n631));
  OR2_X1    g206(.A1(G99), .A2(G2105), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n631), .A2(G2104), .A3(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(G123), .ZN(new_n634));
  OAI221_X1 g209(.A(new_n629), .B1(new_n630), .B2(new_n633), .C1(new_n634), .C2(new_n487), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n635), .A2(G2096), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(G2096), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n628), .A2(new_n636), .A3(new_n637), .ZN(G156));
  INV_X1    g213(.A(KEYINPUT14), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2427), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT15), .B(G2435), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n639), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n643), .B1(new_n642), .B2(new_n641), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2451), .B(G2454), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1341), .B(G1348), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n644), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2443), .B(G2446), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  AND3_X1   g227(.A1(new_n651), .A2(G14), .A3(new_n652), .ZN(G401));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  XNOR2_X1  g229(.A(G2067), .B(G2678), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2072), .B(G2078), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n654), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT85), .B(KEYINPUT17), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n657), .B(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n659), .B1(new_n662), .B2(new_n656), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n654), .A2(new_n655), .A3(new_n657), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT18), .Z(new_n665));
  NAND3_X1  g240(.A1(new_n662), .A2(new_n656), .A3(new_n654), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n663), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2096), .B(G2100), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(G227));
  XOR2_X1   g244(.A(G1971), .B(G1976), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT19), .ZN(new_n671));
  XOR2_X1   g246(.A(G1956), .B(G2474), .Z(new_n672));
  XOR2_X1   g247(.A(G1961), .B(G1966), .Z(new_n673));
  AND2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT20), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n672), .A2(new_n673), .ZN(new_n677));
  NOR3_X1   g252(.A1(new_n671), .A2(new_n674), .A3(new_n677), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n678), .B1(new_n671), .B2(new_n677), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(G1991), .B(G1996), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT86), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n682), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1981), .B(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(G229));
  INV_X1    g262(.A(G16), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(G23), .ZN(new_n689));
  INV_X1    g264(.A(G288), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n689), .B1(new_n690), .B2(new_n688), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT33), .B(G1976), .Z(new_n692));
  OR2_X1    g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n688), .A2(G22), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(G166), .B2(new_n688), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n696), .A2(G1971), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(G1971), .ZN(new_n698));
  NAND4_X1  g273(.A1(new_n693), .A2(new_n694), .A3(new_n697), .A4(new_n698), .ZN(new_n699));
  MUX2_X1   g274(.A(G6), .B(G305), .S(G16), .Z(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT32), .B(G1981), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT34), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n688), .A2(G24), .ZN(new_n706));
  INV_X1    g281(.A(G290), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n706), .B1(new_n707), .B2(new_n688), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(G1986), .ZN(new_n709));
  INV_X1    g284(.A(G29), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G25), .ZN(new_n711));
  INV_X1    g286(.A(G119), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n470), .A2(G107), .ZN(new_n713));
  OAI21_X1  g288(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n714));
  OAI22_X1  g289(.A1(new_n487), .A2(new_n712), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(G131), .B2(new_n492), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n711), .B1(new_n716), .B2(new_n710), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT35), .B(G1991), .Z(new_n718));
  XOR2_X1   g293(.A(new_n717), .B(new_n718), .Z(new_n719));
  NOR2_X1   g294(.A1(new_n709), .A2(new_n719), .ZN(new_n720));
  AND3_X1   g295(.A1(new_n705), .A2(KEYINPUT87), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(KEYINPUT87), .B1(new_n705), .B2(new_n720), .ZN(new_n722));
  OAI22_X1  g297(.A1(new_n721), .A2(new_n722), .B1(new_n704), .B2(new_n703), .ZN(new_n723));
  AND2_X1   g298(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n723), .A2(new_n724), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n710), .B1(KEYINPUT24), .B2(G34), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(KEYINPUT24), .B2(G34), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n485), .B2(G29), .ZN(new_n730));
  INV_X1    g305(.A(G2084), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT99), .Z(new_n733));
  NOR2_X1   g308(.A1(G29), .A2(G35), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(G162), .B2(G29), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT29), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n733), .B1(new_n736), .B2(G2090), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n688), .A2(G4), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(new_n611), .B2(new_n688), .ZN(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT89), .B(G1348), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n740), .A2(new_n741), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n742), .B(new_n743), .C1(new_n731), .C2(new_n730), .ZN(new_n744));
  AOI211_X1 g319(.A(new_n737), .B(new_n744), .C1(G2090), .C2(new_n736), .ZN(new_n745));
  NAND2_X1  g320(.A1(G168), .A2(G16), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n746), .B(KEYINPUT96), .C1(G16), .C2(G21), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(KEYINPUT96), .B2(new_n746), .ZN(new_n748));
  INV_X1    g323(.A(G1966), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT30), .B(G28), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(new_n710), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT31), .B(G11), .ZN(new_n753));
  OAI211_X1 g328(.A(new_n752), .B(new_n753), .C1(new_n635), .C2(new_n710), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT97), .Z(new_n755));
  NAND2_X1  g330(.A1(new_n688), .A2(G5), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G171), .B2(new_n688), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n755), .B1(G1961), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n750), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT98), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n492), .A2(G141), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT94), .ZN(new_n762));
  NAND3_X1  g337(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT95), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT26), .ZN(new_n765));
  INV_X1    g340(.A(new_n487), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n766), .A2(G129), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n476), .A2(G105), .ZN(new_n768));
  NAND4_X1  g343(.A1(new_n762), .A2(new_n765), .A3(new_n767), .A4(new_n768), .ZN(new_n769));
  MUX2_X1   g344(.A(G32), .B(new_n769), .S(G29), .Z(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT27), .ZN(new_n771));
  INV_X1    g346(.A(G1996), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT93), .B(KEYINPUT28), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n710), .A2(G26), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(G104), .A2(G2105), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT91), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n778), .B(G2104), .C1(G116), .C2(new_n470), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT92), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G128), .B2(new_n766), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n492), .A2(G140), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n776), .B1(new_n783), .B2(G29), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G2067), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G1961), .B2(new_n757), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n710), .A2(G27), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G164), .B2(new_n710), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G2078), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n688), .A2(G19), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT90), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(new_n562), .B2(new_n688), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(G1341), .Z(new_n793));
  AOI21_X1  g368(.A(KEYINPUT23), .B1(new_n688), .B2(G20), .ZN(new_n794));
  AND3_X1   g369(.A1(new_n688), .A2(KEYINPUT23), .A3(G20), .ZN(new_n795));
  AOI211_X1 g370(.A(new_n794), .B(new_n795), .C1(G299), .C2(G16), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  XOR2_X1   g372(.A(KEYINPUT100), .B(G1956), .Z(new_n798));
  OR2_X1    g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n797), .A2(new_n798), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT25), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(G139), .ZN(new_n804));
  AOI22_X1  g379(.A1(new_n479), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n805));
  OAI221_X1 g380(.A(new_n803), .B1(new_n473), .B2(new_n804), .C1(new_n805), .C2(new_n470), .ZN(new_n806));
  MUX2_X1   g381(.A(G33), .B(new_n806), .S(G29), .Z(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(G2072), .Z(new_n808));
  NAND4_X1  g383(.A1(new_n793), .A2(new_n799), .A3(new_n800), .A4(new_n808), .ZN(new_n809));
  NOR4_X1   g384(.A1(new_n773), .A2(new_n786), .A3(new_n789), .A4(new_n809), .ZN(new_n810));
  AND2_X1   g385(.A1(new_n760), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n727), .A2(new_n745), .A3(new_n811), .ZN(G150));
  INV_X1    g387(.A(G150), .ZN(G311));
  NAND2_X1  g388(.A1(new_n611), .A2(G559), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT38), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n541), .A2(G67), .ZN(new_n817));
  NAND2_X1  g392(.A1(G80), .A2(G543), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n532), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n521), .A2(G55), .ZN(new_n820));
  INV_X1    g395(.A(G93), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n820), .B1(new_n821), .B2(new_n529), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n620), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n819), .A2(new_n822), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n562), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n816), .B(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT39), .ZN(new_n830));
  AOI21_X1  g405(.A(G860), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(new_n830), .B2(new_n829), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n823), .A2(G860), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT101), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT37), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(KEYINPUT102), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT102), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n832), .A2(new_n838), .A3(new_n835), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n837), .A2(new_n839), .ZN(G145));
  XNOR2_X1  g415(.A(new_n485), .B(new_n635), .ZN(new_n841));
  XNOR2_X1  g416(.A(G162), .B(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n783), .B(new_n806), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(new_n769), .Z(new_n844));
  INV_X1    g419(.A(G130), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n470), .A2(G118), .ZN(new_n846));
  OAI21_X1  g421(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n847));
  OAI22_X1  g422(.A1(new_n487), .A2(new_n845), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(G142), .B2(new_n492), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n626), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n716), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n479), .A2(new_n498), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n509), .B1(new_n469), .B2(new_n501), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n851), .B(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n844), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n844), .A2(new_n857), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n842), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n844), .A2(new_n857), .ZN(new_n862));
  INV_X1    g437(.A(new_n842), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n862), .A2(new_n863), .A3(new_n858), .ZN(new_n864));
  INV_X1    g439(.A(G37), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n861), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g442(.A(G290), .B(G305), .Z(new_n868));
  XNOR2_X1  g443(.A(G166), .B(G288), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n868), .B(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT42), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n622), .B(new_n827), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n609), .B(G299), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT41), .ZN(new_n874));
  AOI21_X1  g449(.A(KEYINPUT103), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n872), .A2(new_n873), .ZN(new_n876));
  OR2_X1    g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  OR3_X1    g452(.A1(new_n872), .A2(KEYINPUT103), .A3(new_n873), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n871), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI211_X1 g454(.A(new_n878), .B(new_n871), .C1(new_n876), .C2(new_n875), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  OAI21_X1  g456(.A(G868), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n882), .B1(G868), .B2(new_n825), .ZN(G295));
  OAI21_X1  g458(.A(new_n882), .B1(G868), .B2(new_n825), .ZN(G331));
  XNOR2_X1  g459(.A(G171), .B(G168), .ZN(new_n885));
  AND2_X1   g460(.A1(new_n827), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n886), .A2(new_n873), .ZN(new_n887));
  OAI21_X1  g462(.A(KEYINPUT104), .B1(new_n827), .B2(new_n885), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n827), .A2(new_n885), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT104), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n887), .A2(new_n888), .A3(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n874), .B1(new_n886), .B2(new_n889), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n892), .A2(new_n893), .A3(new_n870), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(new_n865), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n892), .A2(new_n893), .ZN(new_n897));
  INV_X1    g472(.A(new_n870), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(KEYINPUT43), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n891), .A2(new_n888), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n874), .B1(new_n901), .B2(new_n886), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n887), .B1(new_n827), .B2(new_n885), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n870), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT43), .ZN(new_n905));
  NOR3_X1   g480(.A1(new_n895), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(KEYINPUT44), .B1(new_n900), .B2(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n905), .B1(new_n896), .B2(new_n899), .ZN(new_n908));
  NOR3_X1   g483(.A1(new_n895), .A2(new_n904), .A3(KEYINPUT43), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n907), .B1(new_n910), .B2(KEYINPUT44), .ZN(G397));
  NAND3_X1  g486(.A1(new_n477), .A2(G40), .A3(new_n484), .ZN(new_n912));
  INV_X1    g487(.A(G1384), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n514), .A2(new_n502), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n913), .B1(new_n499), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT45), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n912), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n769), .B(new_n772), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n783), .A2(G2067), .ZN(new_n920));
  INV_X1    g495(.A(G2067), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n781), .A2(new_n921), .A3(new_n782), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n919), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n716), .B(new_n718), .ZN(new_n924));
  OR2_X1    g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(G290), .A2(G1986), .ZN(new_n926));
  XOR2_X1   g501(.A(new_n926), .B(KEYINPUT106), .Z(new_n927));
  NOR2_X1   g502(.A1(G290), .A2(G1986), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n928), .B(KEYINPUT105), .ZN(new_n929));
  OR2_X1    g504(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n918), .B1(new_n925), .B2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT54), .ZN(new_n932));
  XOR2_X1   g507(.A(new_n477), .B(KEYINPUT123), .Z(new_n933));
  AOI21_X1  g508(.A(new_n470), .B1(new_n483), .B2(KEYINPUT124), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n934), .B1(KEYINPUT124), .B2(new_n483), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT53), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n936), .A2(G2078), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n935), .A2(G40), .A3(new_n917), .A4(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n933), .A2(new_n938), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n856), .A2(KEYINPUT108), .A3(KEYINPUT45), .A4(new_n913), .ZN(new_n940));
  OAI211_X1 g515(.A(KEYINPUT45), .B(new_n913), .C1(new_n499), .C2(new_n914), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT108), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT50), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n514), .A2(KEYINPUT74), .A3(new_n502), .ZN(new_n946));
  AOI21_X1  g521(.A(KEYINPUT74), .B1(new_n514), .B2(new_n502), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n854), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n945), .B1(new_n948), .B2(new_n913), .ZN(new_n949));
  XNOR2_X1  g524(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n913), .B(new_n950), .C1(new_n499), .C2(new_n914), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n477), .A2(new_n951), .A3(G40), .A4(new_n484), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(G1961), .ZN(new_n955));
  AOI22_X1  g530(.A1(new_n939), .A2(new_n944), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT109), .ZN(new_n957));
  INV_X1    g532(.A(new_n912), .ZN(new_n958));
  AOI21_X1  g533(.A(KEYINPUT45), .B1(new_n948), .B2(new_n913), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT107), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n958), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n960), .B(new_n916), .C1(G164), .C2(G1384), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n944), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n957), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  AOI22_X1  g539(.A1(new_n959), .A2(new_n960), .B1(new_n943), .B2(new_n940), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n916), .B1(G164), .B2(G1384), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n912), .B1(new_n966), .B2(KEYINPUT107), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n965), .A2(new_n967), .A3(KEYINPUT109), .ZN(new_n968));
  AOI21_X1  g543(.A(G2078), .B1(new_n964), .B2(new_n968), .ZN(new_n969));
  OAI211_X1 g544(.A(new_n956), .B(G301), .C1(new_n969), .C2(KEYINPUT53), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n954), .A2(new_n955), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT45), .B1(new_n856), .B2(new_n913), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n912), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n948), .A2(KEYINPUT45), .A3(new_n913), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n973), .A2(new_n974), .A3(new_n937), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n971), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(G2078), .ZN(new_n977));
  NOR3_X1   g552(.A1(new_n961), .A2(new_n963), .A3(new_n957), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT109), .B1(new_n965), .B2(new_n967), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n977), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n976), .B1(new_n980), .B2(new_n936), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n970), .B1(new_n981), .B2(G301), .ZN(new_n982));
  NAND2_X1  g557(.A1(G286), .A2(G8), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n917), .A2(G40), .A3(new_n484), .A4(new_n477), .ZN(new_n985));
  NOR3_X1   g560(.A1(G164), .A2(new_n916), .A3(G1384), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n749), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n988));
  XNOR2_X1  g563(.A(KEYINPUT117), .B(G2084), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n958), .A2(new_n988), .A3(new_n951), .A4(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  AOI211_X1 g566(.A(KEYINPUT51), .B(new_n984), .C1(new_n991), .C2(G8), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n983), .B(KEYINPUT122), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT121), .ZN(new_n995));
  AOI21_X1  g570(.A(G1966), .B1(new_n973), .B2(new_n974), .ZN(new_n996));
  INV_X1    g571(.A(new_n989), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n949), .A2(new_n952), .A3(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n995), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n987), .A2(new_n990), .A3(KEYINPUT121), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n994), .B1(new_n1001), .B2(G8), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT51), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n993), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1001), .A2(new_n984), .ZN(new_n1005));
  AOI22_X1  g580(.A1(new_n932), .A2(new_n982), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(G1971), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n964), .A2(new_n968), .A3(new_n1007), .ZN(new_n1008));
  OR2_X1    g583(.A1(new_n954), .A2(G2090), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(G8), .ZN(new_n1011));
  NOR2_X1   g586(.A1(G166), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT111), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1012), .B1(new_n1013), .B2(KEYINPUT55), .ZN(new_n1014));
  XNOR2_X1  g589(.A(KEYINPUT111), .B(KEYINPUT55), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1014), .B1(new_n1012), .B2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1010), .A2(G8), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n915), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1018), .A2(new_n477), .A3(G40), .A4(new_n484), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(G8), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n579), .B(G1976), .C1(new_n532), .C2(new_n580), .ZN(new_n1022));
  OR2_X1    g597(.A1(new_n1022), .A2(KEYINPUT112), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(KEYINPUT112), .ZN(new_n1024));
  INV_X1    g599(.A(G1976), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT52), .B1(G288), .B2(new_n1025), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1021), .A2(new_n1023), .A3(new_n1024), .A4(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1028));
  OAI21_X1  g603(.A(KEYINPUT52), .B1(new_n1028), .B2(new_n1020), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT113), .ZN(new_n1031));
  INV_X1    g606(.A(G1981), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n588), .A2(new_n1032), .A3(new_n589), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1032), .B1(new_n588), .B2(new_n589), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1031), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1020), .B1(new_n1036), .B2(KEYINPUT49), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1035), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT113), .B1(new_n1038), .B2(new_n1033), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT49), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1037), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT114), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1037), .A2(KEYINPUT114), .A3(new_n1041), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1030), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1017), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1016), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n958), .B1(new_n1018), .B2(new_n950), .ZN(new_n1049));
  NOR3_X1   g624(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1050));
  OR3_X1    g625(.A1(new_n1049), .A2(G2090), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1008), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(KEYINPUT116), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT116), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1008), .A2(new_n1051), .A3(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1053), .A2(G8), .A3(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1047), .B1(new_n1048), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G1956), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1058), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1059));
  XOR2_X1   g634(.A(G299), .B(KEYINPUT57), .Z(new_n1060));
  XNOR2_X1  g635(.A(KEYINPUT56), .B(G2072), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n965), .A2(new_n967), .A3(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1059), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1060), .B1(new_n1059), .B2(new_n1062), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT120), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n958), .A2(new_n1065), .A3(new_n921), .A4(new_n1018), .ZN(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT120), .B1(new_n1019), .B2(G2067), .ZN(new_n1067));
  INV_X1    g642(.A(G1348), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1068), .B1(new_n949), .B2(new_n952), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1066), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n609), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1063), .B1(new_n1064), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1064), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1074), .A2(KEYINPUT61), .A3(new_n1063), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT61), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1063), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1076), .B1(new_n1077), .B2(new_n1064), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1071), .A2(KEYINPUT60), .ZN(new_n1080));
  XNOR2_X1  g655(.A(new_n1070), .B(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1071), .A2(KEYINPUT60), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT59), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n965), .A2(new_n967), .A3(new_n772), .ZN(new_n1084));
  XOR2_X1   g659(.A(KEYINPUT58), .B(G1341), .Z(new_n1085));
  NAND2_X1  g660(.A1(new_n1019), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1083), .B1(new_n1087), .B2(new_n562), .ZN(new_n1088));
  AOI211_X1 g663(.A(KEYINPUT59), .B(new_n620), .C1(new_n1084), .C2(new_n1086), .ZN(new_n1089));
  OAI22_X1  g664(.A1(new_n1081), .A2(new_n1082), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1073), .B1(new_n1079), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n939), .A2(new_n944), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(new_n971), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1093), .B1(new_n980), .B2(new_n936), .ZN(new_n1094));
  OAI21_X1  g669(.A(KEYINPUT125), .B1(new_n1094), .B2(G301), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n932), .B1(new_n981), .B2(G301), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n956), .B1(new_n969), .B2(KEYINPUT53), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT125), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1097), .A2(new_n1098), .A3(G171), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1095), .A2(new_n1096), .A3(new_n1099), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1006), .A2(new_n1057), .A3(new_n1091), .A4(new_n1100), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n987), .A2(KEYINPUT121), .A3(new_n990), .ZN(new_n1102));
  AOI21_X1  g677(.A(KEYINPUT121), .B1(new_n987), .B2(new_n990), .ZN(new_n1103));
  OAI21_X1  g678(.A(G8), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n994), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1003), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1005), .B1(new_n1106), .B2(new_n992), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(KEYINPUT62), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT62), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1004), .A2(new_n1109), .A3(new_n1005), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n981), .A2(G301), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1057), .A2(new_n1108), .A3(new_n1110), .A4(new_n1111), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1113));
  NOR3_X1   g688(.A1(new_n1017), .A2(new_n1113), .A3(new_n1030), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n690), .A2(new_n1025), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1033), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  XOR2_X1   g691(.A(new_n1020), .B(KEYINPUT115), .Z(new_n1117));
  AOI21_X1  g692(.A(new_n1114), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1101), .A2(new_n1112), .A3(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n991), .A2(G8), .A3(G168), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT118), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n991), .A2(KEYINPUT118), .A3(G8), .A4(G168), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(KEYINPUT63), .B1(new_n1057), .B2(new_n1124), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1017), .A2(new_n1046), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT119), .ZN(new_n1127));
  AND2_X1   g702(.A1(new_n1124), .A2(KEYINPUT63), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1011), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1129));
  OR2_X1    g704(.A1(new_n1129), .A2(new_n1016), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1126), .A2(new_n1127), .A3(new_n1128), .A4(new_n1130), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1124), .B(KEYINPUT63), .C1(new_n1129), .C2(new_n1016), .ZN(new_n1132));
  OAI21_X1  g707(.A(KEYINPUT119), .B1(new_n1132), .B2(new_n1047), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1125), .A2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n931), .B1(new_n1119), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(KEYINPUT48), .B1(new_n929), .B2(new_n918), .ZN(new_n1137));
  AND3_X1   g712(.A1(new_n929), .A2(KEYINPUT48), .A3(new_n918), .ZN(new_n1138));
  AOI211_X1 g713(.A(new_n1137), .B(new_n1138), .C1(new_n918), .C2(new_n925), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n920), .A2(new_n922), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n918), .B1(new_n1140), .B2(new_n769), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT46), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1142), .B1(new_n918), .B2(new_n772), .ZN(new_n1143));
  NOR4_X1   g718(.A1(new_n912), .A2(new_n917), .A3(KEYINPUT46), .A4(G1996), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1141), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  XOR2_X1   g720(.A(new_n1145), .B(KEYINPUT47), .Z(new_n1146));
  NAND2_X1  g721(.A1(new_n716), .A2(new_n718), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n922), .B1(new_n923), .B2(new_n1147), .ZN(new_n1148));
  AOI211_X1 g723(.A(new_n1139), .B(new_n1146), .C1(new_n918), .C2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1136), .A2(new_n1149), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g725(.A1(G401), .A2(new_n461), .A3(G227), .ZN(new_n1152));
  XOR2_X1   g726(.A(new_n1152), .B(KEYINPUT126), .Z(new_n1153));
  NOR2_X1   g727(.A1(new_n1153), .A2(G229), .ZN(new_n1154));
  OAI211_X1 g728(.A(new_n866), .B(new_n1154), .C1(new_n908), .C2(new_n909), .ZN(G225));
  INV_X1    g729(.A(G225), .ZN(G308));
endmodule


