//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 1 0 1 1 0 1 1 0 0 1 0 0 0 1 0 1 1 0 1 0 0 1 0 1 1 0 1 0 1 0 1 0 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:42 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(G237), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(new_n189), .A3(G214), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  NOR2_X1   g006(.A1(G237), .A2(G953), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(G143), .A3(G214), .ZN(new_n194));
  NAND2_X1  g008(.A1(KEYINPUT18), .A2(G131), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n192), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(G125), .B(G140), .ZN(new_n197));
  INV_X1    g011(.A(G146), .ZN(new_n198));
  XNOR2_X1  g012(.A(new_n197), .B(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT88), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n192), .A2(new_n194), .ZN(new_n201));
  INV_X1    g015(.A(new_n195), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n200), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  AOI211_X1 g017(.A(KEYINPUT88), .B(new_n195), .C1(new_n192), .C2(new_n194), .ZN(new_n204));
  OAI211_X1 g018(.A(new_n196), .B(new_n199), .C1(new_n203), .C2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G125), .ZN(new_n206));
  NOR3_X1   g020(.A1(new_n206), .A2(KEYINPUT16), .A3(G140), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n207), .B1(new_n197), .B2(KEYINPUT16), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT75), .B1(new_n208), .B2(G146), .ZN(new_n209));
  INV_X1    g023(.A(G140), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G125), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n206), .A2(G140), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n211), .A2(new_n212), .A3(KEYINPUT16), .ZN(new_n213));
  OR3_X1    g027(.A1(new_n206), .A2(KEYINPUT16), .A3(G140), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT75), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n215), .A2(new_n216), .A3(new_n198), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT74), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n218), .B1(new_n208), .B2(G146), .ZN(new_n219));
  AND4_X1   g033(.A1(new_n218), .A2(new_n213), .A3(G146), .A4(new_n214), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n209), .B(new_n217), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G131), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n222), .B1(new_n192), .B2(new_n194), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(KEYINPUT17), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n193), .A2(G143), .A3(G214), .ZN(new_n225));
  AOI21_X1  g039(.A(G143), .B1(new_n193), .B2(G214), .ZN(new_n226));
  OAI21_X1  g040(.A(G131), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n192), .A2(new_n222), .A3(new_n194), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n224), .B1(new_n229), .B2(KEYINPUT17), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n205), .B1(new_n221), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g045(.A(G113), .B(G122), .ZN(new_n232));
  INV_X1    g046(.A(G104), .ZN(new_n233));
  XNOR2_X1  g047(.A(new_n232), .B(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  AND2_X1   g049(.A1(new_n231), .A2(new_n235), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n234), .B(new_n205), .C1(new_n221), .C2(new_n230), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n187), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G475), .ZN(new_n240));
  NOR2_X1   g054(.A1(G475), .A2(G902), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT91), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n211), .A2(new_n212), .A3(KEYINPUT90), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT19), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n211), .A2(new_n212), .A3(KEYINPUT90), .A4(KEYINPUT19), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n243), .B1(new_n248), .B2(new_n198), .ZN(new_n249));
  AOI211_X1 g063(.A(KEYINPUT91), .B(G146), .C1(new_n246), .C2(new_n247), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NOR3_X1   g065(.A1(new_n225), .A2(new_n226), .A3(G131), .ZN(new_n252));
  OAI21_X1  g066(.A(KEYINPUT89), .B1(new_n252), .B2(new_n223), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n215), .A2(new_n198), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT89), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n227), .A2(new_n256), .A3(new_n228), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n253), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n205), .B1(new_n251), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(new_n235), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n242), .B1(new_n260), .B2(new_n237), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT20), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT92), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n254), .B1(new_n229), .B2(KEYINPUT89), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n264), .B(new_n257), .C1(new_n250), .C2(new_n249), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n234), .B1(new_n265), .B2(new_n205), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n241), .B1(new_n266), .B2(new_n238), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT92), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n267), .A2(new_n268), .A3(KEYINPUT20), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n262), .B(new_n241), .C1(new_n266), .C2(new_n238), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT93), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n260), .A2(new_n237), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n273), .A2(KEYINPUT93), .A3(new_n262), .A4(new_n241), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n263), .A2(new_n269), .A3(new_n272), .A4(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G478), .ZN(new_n276));
  XNOR2_X1  g090(.A(KEYINPUT9), .B(G234), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n278), .A2(G217), .A3(new_n189), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT13), .ZN(new_n280));
  INV_X1    g094(.A(G128), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n280), .B1(new_n281), .B2(G143), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(G143), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n191), .A2(G128), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n285), .A2(new_n280), .ZN(new_n286));
  OAI21_X1  g100(.A(G134), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G134), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n285), .A2(new_n283), .A3(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G122), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G116), .ZN(new_n291));
  INV_X1    g105(.A(G116), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G122), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(KEYINPUT78), .B(G107), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n296), .A2(new_n291), .A3(new_n293), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n287), .B(new_n289), .C1(new_n297), .C2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT94), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n285), .A2(new_n283), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G134), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n289), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n292), .A2(KEYINPUT14), .A3(G122), .ZN(new_n304));
  OAI211_X1 g118(.A(G107), .B(new_n304), .C1(new_n294), .C2(KEYINPUT14), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n295), .A2(new_n296), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n303), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n299), .A2(new_n300), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n300), .B1(new_n299), .B2(new_n307), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n279), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n299), .A2(new_n307), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(KEYINPUT94), .ZN(new_n313));
  INV_X1    g127(.A(new_n279), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n313), .A2(new_n314), .A3(new_n308), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  AOI211_X1 g130(.A(KEYINPUT15), .B(new_n276), .C1(new_n316), .C2(new_n187), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n187), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n276), .A2(KEYINPUT15), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n189), .A2(G952), .ZN(new_n322));
  NAND2_X1  g136(.A1(G234), .A2(G237), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  XOR2_X1   g138(.A(new_n324), .B(KEYINPUT95), .Z(new_n325));
  AND3_X1   g139(.A1(new_n323), .A2(G902), .A3(G953), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT21), .B(G898), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AND2_X1   g142(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  AND4_X1   g144(.A1(new_n240), .A2(new_n275), .A3(new_n321), .A4(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(G221), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n332), .B1(new_n278), .B2(new_n187), .ZN(new_n333));
  INV_X1    g147(.A(G469), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n334), .A2(new_n187), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n198), .A2(G143), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n191), .A2(G146), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT1), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n336), .A2(new_n337), .A3(new_n338), .A4(G128), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(KEYINPUT79), .ZN(new_n340));
  XNOR2_X1  g154(.A(G143), .B(G146), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT79), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n341), .A2(new_n342), .A3(new_n338), .A4(G128), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n336), .A2(new_n337), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(new_n281), .ZN(new_n345));
  INV_X1    g159(.A(new_n337), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT1), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n340), .A2(new_n343), .A3(new_n345), .A4(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n233), .A2(KEYINPUT3), .ZN(new_n349));
  INV_X1    g163(.A(G107), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT78), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT78), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(G107), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n349), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G101), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n233), .A2(G107), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n350), .A2(G104), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(KEYINPUT3), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n354), .A2(new_n355), .A3(new_n356), .A4(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(G104), .B1(new_n351), .B2(new_n353), .ZN(new_n360));
  INV_X1    g174(.A(new_n357), .ZN(new_n361));
  OAI21_X1  g175(.A(G101), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n348), .A2(new_n359), .A3(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n354), .A2(new_n356), .A3(new_n358), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G101), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n367), .A2(KEYINPUT4), .A3(new_n359), .ZN(new_n368));
  NAND2_X1  g182(.A1(KEYINPUT0), .A2(G128), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n336), .A2(new_n337), .A3(new_n369), .ZN(new_n370));
  XOR2_X1   g184(.A(KEYINPUT0), .B(G128), .Z(new_n371));
  OAI21_X1  g185(.A(new_n370), .B1(new_n371), .B2(new_n341), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n355), .A2(KEYINPUT4), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n366), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n368), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n362), .A2(new_n359), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n345), .A2(new_n347), .A3(new_n339), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(KEYINPUT10), .A3(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT11), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n380), .B1(new_n288), .B2(G137), .ZN(new_n381));
  INV_X1    g195(.A(G137), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(KEYINPUT11), .A3(G134), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n288), .A2(G137), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n381), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G131), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n381), .A2(new_n383), .A3(new_n222), .A4(new_n384), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(KEYINPUT64), .A3(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT64), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n385), .A2(new_n389), .A3(G131), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n365), .A2(new_n375), .A3(new_n379), .A4(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n378), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n376), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n391), .B1(new_n363), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT12), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT80), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n396), .B1(new_n391), .B2(new_n397), .ZN(new_n398));
  AND2_X1   g212(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n395), .A2(new_n398), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n392), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(G110), .B(G140), .ZN(new_n402));
  AND2_X1   g216(.A1(new_n189), .A2(G227), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n402), .B(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  AND2_X1   g219(.A1(new_n392), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n365), .A2(new_n375), .A3(new_n379), .ZN(new_n407));
  INV_X1    g221(.A(new_n391), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI22_X1  g223(.A1(new_n401), .A2(new_n404), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n335), .B1(new_n410), .B2(G469), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n392), .A2(new_n405), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n395), .A2(new_n398), .ZN(new_n413));
  OR2_X1    g227(.A1(new_n395), .A2(new_n398), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n405), .B1(new_n409), .B2(new_n392), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n334), .B(new_n187), .C1(new_n415), .C2(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n333), .B1(new_n411), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n331), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(G210), .B1(G237), .B2(G902), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n420), .B(KEYINPUT86), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n370), .B(G125), .C1(new_n371), .C2(new_n341), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n423), .B1(new_n378), .B2(G125), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n189), .A2(G224), .ZN(new_n425));
  XOR2_X1   g239(.A(new_n424), .B(new_n425), .Z(new_n426));
  INV_X1    g240(.A(G119), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT65), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT65), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(G119), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n428), .A2(new_n430), .A3(G116), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n292), .A2(G119), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n431), .A2(KEYINPUT5), .A3(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(KEYINPUT65), .B(G119), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT5), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n434), .A2(new_n435), .A3(G116), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n433), .A2(G113), .A3(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(G113), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(KEYINPUT2), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT2), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(G113), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n431), .A2(new_n432), .A3(new_n442), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n437), .A2(new_n443), .A3(new_n359), .A4(new_n362), .ZN(new_n444));
  XNOR2_X1  g258(.A(G110), .B(G122), .ZN(new_n445));
  AOI22_X1  g259(.A1(new_n296), .A2(new_n349), .B1(KEYINPUT3), .B2(new_n357), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n355), .B1(new_n446), .B2(new_n356), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n359), .A2(KEYINPUT4), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n443), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n442), .B1(new_n431), .B2(new_n432), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n374), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n444), .B(new_n445), .C1(new_n449), .C2(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n444), .B1(new_n449), .B2(new_n452), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n445), .B(KEYINPUT81), .ZN(new_n455));
  AOI22_X1  g269(.A1(new_n453), .A2(KEYINPUT6), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  AND3_X1   g270(.A1(new_n454), .A2(KEYINPUT6), .A3(new_n455), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n426), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n425), .A2(KEYINPUT7), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT84), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n459), .B1(new_n423), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n424), .A2(new_n461), .ZN(new_n462));
  OAI221_X1 g276(.A(new_n423), .B1(new_n460), .B2(new_n459), .C1(new_n378), .C2(G125), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n451), .ZN(new_n465));
  AOI22_X1  g279(.A1(new_n465), .A2(new_n443), .B1(new_n366), .B2(new_n373), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n362), .A2(new_n359), .A3(new_n443), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  AOI22_X1  g282(.A1(new_n466), .A2(new_n368), .B1(new_n468), .B2(new_n437), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n464), .B1(new_n469), .B2(new_n445), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n445), .B(KEYINPUT8), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n436), .A2(KEYINPUT83), .A3(G113), .ZN(new_n472));
  AOI21_X1  g286(.A(KEYINPUT83), .B1(new_n436), .B2(G113), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n433), .B(KEYINPUT82), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n467), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n377), .B1(new_n443), .B2(new_n437), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n471), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(G902), .B1(new_n470), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n458), .A2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT85), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n422), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n458), .A2(KEYINPUT85), .A3(new_n479), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT87), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n485), .B1(new_n480), .B2(new_n421), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n482), .A2(KEYINPUT87), .A3(new_n483), .ZN(new_n489));
  OAI21_X1  g303(.A(G214), .B1(G237), .B2(G902), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n419), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(G472), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n388), .A2(new_n390), .A3(new_n372), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n288), .A2(G137), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n382), .A2(G134), .ZN(new_n496));
  OAI21_X1  g310(.A(G131), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  AND2_X1   g311(.A1(new_n387), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n378), .ZN(new_n499));
  AOI21_X1  g313(.A(KEYINPUT30), .B1(new_n494), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n465), .A2(new_n443), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT30), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n503), .B1(new_n498), .B2(new_n378), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n494), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n501), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT66), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n507), .B1(new_n450), .B2(new_n451), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n465), .A2(KEYINPUT66), .A3(new_n443), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n494), .A2(new_n499), .A3(new_n508), .A4(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n193), .A2(G210), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n511), .B(KEYINPUT27), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT26), .B(G101), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n512), .B(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n506), .A2(new_n510), .A3(new_n515), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n516), .A2(KEYINPUT29), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n517), .A2(G902), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT28), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n494), .A2(new_n499), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n508), .A2(new_n509), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n519), .B1(new_n522), .B2(new_n510), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n510), .A2(new_n519), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(KEYINPUT29), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  XOR2_X1   g340(.A(KEYINPUT68), .B(KEYINPUT28), .Z(new_n527));
  AND4_X1   g341(.A1(new_n494), .A2(new_n499), .A3(new_n508), .A4(new_n509), .ZN(new_n528));
  AOI22_X1  g342(.A1(new_n494), .A2(new_n499), .B1(new_n465), .B2(new_n443), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n524), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n526), .B(new_n514), .C1(KEYINPUT29), .C2(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n493), .B1(new_n518), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT67), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n505), .A2(new_n502), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n510), .B(new_n514), .C1(new_n535), .C2(new_n500), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n534), .B1(new_n536), .B2(KEYINPUT31), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n528), .A2(new_n515), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT31), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n506), .A2(new_n538), .A3(KEYINPUT67), .A4(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n531), .A2(new_n515), .B1(KEYINPUT31), .B2(new_n536), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT69), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n541), .A2(new_n542), .A3(KEYINPUT69), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(G472), .A2(G902), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT32), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n533), .B1(new_n547), .B2(new_n551), .ZN(new_n552));
  AND3_X1   g366(.A1(new_n541), .A2(new_n542), .A3(KEYINPUT69), .ZN(new_n553));
  AOI21_X1  g367(.A(KEYINPUT69), .B1(new_n541), .B2(new_n542), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n548), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n550), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT77), .ZN(new_n558));
  INV_X1    g372(.A(G234), .ZN(new_n559));
  OAI21_X1  g373(.A(G217), .B1(new_n559), .B2(G902), .ZN(new_n560));
  XOR2_X1   g374(.A(new_n560), .B(KEYINPUT70), .Z(new_n561));
  NAND3_X1  g375(.A1(new_n428), .A2(new_n430), .A3(G128), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n562), .B1(new_n427), .B2(G128), .ZN(new_n563));
  XNOR2_X1  g377(.A(KEYINPUT24), .B(G110), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT23), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(KEYINPUT71), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT71), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(KEYINPUT23), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n562), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(KEYINPUT72), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT72), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n562), .A2(new_n572), .A3(new_n569), .ZN(new_n573));
  OAI21_X1  g387(.A(KEYINPUT73), .B1(new_n434), .B2(G128), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n428), .A2(new_n430), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT73), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n575), .A2(new_n576), .A3(new_n281), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n571), .A2(new_n573), .A3(new_n574), .A4(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n281), .A2(KEYINPUT23), .A3(G119), .ZN(new_n579));
  AND2_X1   g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(G110), .ZN(new_n581));
  OAI221_X1 g395(.A(new_n221), .B1(new_n563), .B2(new_n564), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT76), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n578), .A2(new_n581), .A3(new_n579), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n563), .A2(new_n564), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n197), .A2(new_n198), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n255), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n583), .B1(new_n586), .B2(new_n589), .ZN(new_n590));
  AOI211_X1 g404(.A(KEYINPUT76), .B(new_n588), .C1(new_n584), .C2(new_n585), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n582), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(KEYINPUT22), .B(G137), .ZN(new_n593));
  NOR3_X1   g407(.A1(new_n332), .A2(new_n559), .A3(G953), .ZN(new_n594));
  XOR2_X1   g408(.A(new_n593), .B(new_n594), .Z(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n582), .B(new_n595), .C1(new_n590), .C2(new_n591), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n597), .A2(new_n187), .A3(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT25), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n597), .A2(KEYINPUT25), .A3(new_n187), .A4(new_n598), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n561), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n597), .A2(new_n598), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n560), .A2(new_n187), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n557), .A2(new_n558), .A3(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n558), .B1(new_n557), .B2(new_n607), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n492), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(G101), .ZN(G3));
  INV_X1    g426(.A(new_n607), .ZN(new_n613));
  AOI21_X1  g427(.A(G902), .B1(new_n545), .B2(new_n546), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n555), .B1(new_n614), .B2(new_n493), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n406), .A2(new_n409), .ZN(new_n616));
  INV_X1    g430(.A(new_n407), .ZN(new_n617));
  AOI22_X1  g431(.A1(new_n413), .A2(new_n414), .B1(new_n617), .B2(new_n391), .ZN(new_n618));
  OAI211_X1 g432(.A(new_n616), .B(G469), .C1(new_n618), .C2(new_n405), .ZN(new_n619));
  INV_X1    g433(.A(new_n335), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n417), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n333), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n613), .A2(new_n615), .A3(new_n623), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n458), .A2(new_n479), .A3(new_n422), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n422), .B1(new_n458), .B2(new_n479), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n490), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT96), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OAI211_X1 g443(.A(KEYINPUT96), .B(new_n490), .C1(new_n625), .C2(new_n626), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n318), .A2(new_n276), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n276), .A2(G902), .ZN(new_n633));
  AOI21_X1  g447(.A(KEYINPUT33), .B1(new_n316), .B2(KEYINPUT97), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT97), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT33), .ZN(new_n636));
  AOI211_X1 g450(.A(new_n635), .B(new_n636), .C1(new_n311), .C2(new_n315), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n633), .B1(new_n634), .B2(new_n637), .ZN(new_n638));
  AOI22_X1  g452(.A1(new_n275), .A2(new_n240), .B1(new_n632), .B2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n631), .A2(new_n640), .A3(new_n329), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n624), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT34), .B(G104), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G6));
  NAND3_X1  g458(.A1(new_n263), .A2(new_n269), .A3(new_n270), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n240), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n646), .A2(new_n321), .ZN(new_n647));
  AND4_X1   g461(.A1(new_n330), .A2(new_n647), .A3(new_n629), .A4(new_n630), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n624), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT35), .B(G107), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G9));
  NOR3_X1   g465(.A1(new_n615), .A2(new_n419), .A3(new_n491), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n601), .A2(new_n602), .ZN(new_n653));
  INV_X1    g467(.A(new_n561), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  OR2_X1    g469(.A1(new_n596), .A2(KEYINPUT36), .ZN(new_n656));
  OR2_X1    g470(.A1(new_n592), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n592), .A2(new_n656), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n659), .A2(new_n605), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n655), .A2(KEYINPUT98), .A3(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT98), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n663), .B1(new_n603), .B2(new_n660), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n652), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT37), .B(G110), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT99), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n666), .B(new_n668), .ZN(G12));
  NAND3_X1  g483(.A1(new_n629), .A2(new_n418), .A3(new_n630), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n670), .B1(new_n556), .B2(new_n552), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n325), .B(KEYINPUT101), .ZN(new_n672));
  INV_X1    g486(.A(G900), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(KEYINPUT100), .ZN(new_n674));
  OR2_X1    g488(.A1(new_n673), .A2(KEYINPUT100), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n326), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(KEYINPUT102), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n646), .A2(new_n321), .A3(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n671), .A2(new_n665), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G128), .ZN(G30));
  INV_X1    g495(.A(new_n489), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n486), .B1(new_n483), .B2(new_n482), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n685));
  XOR2_X1   g499(.A(new_n684), .B(new_n685), .Z(new_n686));
  NAND2_X1  g500(.A1(new_n506), .A2(new_n510), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n514), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n522), .A2(new_n510), .ZN(new_n689));
  AOI21_X1  g503(.A(G902), .B1(new_n689), .B2(new_n515), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n493), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n691), .B1(new_n547), .B2(new_n551), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT104), .ZN(new_n693));
  AND3_X1   g507(.A1(new_n692), .A2(new_n693), .A3(new_n556), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n693), .B1(new_n692), .B2(new_n556), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XOR2_X1   g510(.A(new_n678), .B(KEYINPUT39), .Z(new_n697));
  NAND2_X1  g511(.A1(new_n418), .A2(new_n697), .ZN(new_n698));
  OR2_X1    g512(.A1(new_n698), .A2(KEYINPUT40), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(KEYINPUT40), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n275), .A2(new_n240), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(new_n490), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n702), .A2(new_n703), .A3(new_n321), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n699), .A2(new_n700), .A3(new_n704), .ZN(new_n705));
  OR4_X1    g519(.A1(new_n665), .A2(new_n686), .A3(new_n696), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G143), .ZN(G45));
  NAND2_X1  g521(.A1(new_n638), .A2(new_n632), .ZN(new_n708));
  INV_X1    g522(.A(new_n678), .ZN(new_n709));
  AND4_X1   g523(.A1(KEYINPUT105), .A2(new_n701), .A3(new_n708), .A4(new_n709), .ZN(new_n710));
  AOI21_X1  g524(.A(KEYINPUT105), .B1(new_n639), .B2(new_n709), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n671), .A2(new_n665), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT106), .B(G146), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G48));
  OAI21_X1  g529(.A(new_n187), .B1(new_n415), .B2(new_n416), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(G469), .ZN(new_n717));
  AND3_X1   g531(.A1(new_n717), .A2(new_n622), .A3(new_n417), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n641), .A2(new_n557), .A3(new_n607), .A4(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(KEYINPUT41), .B(G113), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G15));
  NAND4_X1  g535(.A1(new_n648), .A2(new_n557), .A3(new_n607), .A4(new_n718), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G116), .ZN(G18));
  AND4_X1   g537(.A1(new_n331), .A2(new_n629), .A3(new_n630), .A4(new_n718), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n665), .A2(new_n557), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G119), .ZN(G21));
  AND4_X1   g540(.A1(new_n330), .A2(new_n718), .A3(new_n629), .A4(new_n630), .ZN(new_n727));
  INV_X1    g541(.A(new_n321), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n701), .A2(KEYINPUT107), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(KEYINPUT107), .B1(new_n701), .B2(new_n728), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n524), .B1(new_n689), .B2(new_n519), .ZN(new_n732));
  AOI22_X1  g546(.A1(new_n732), .A2(new_n515), .B1(KEYINPUT31), .B2(new_n536), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n549), .B1(new_n733), .B2(new_n541), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n547), .A2(new_n187), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n734), .B1(new_n735), .B2(G472), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n727), .A2(new_n731), .A3(new_n736), .A4(new_n607), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G122), .ZN(G24));
  AND3_X1   g552(.A1(new_n718), .A2(new_n629), .A3(new_n630), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n665), .A2(new_n712), .A3(new_n739), .A4(new_n736), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G125), .ZN(G27));
  INV_X1    g555(.A(KEYINPUT42), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT108), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n623), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n418), .A2(KEYINPUT108), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n703), .B1(new_n488), .B2(new_n489), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n747), .A2(new_n557), .A3(new_n607), .A4(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n712), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n742), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n557), .A2(new_n607), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n490), .B1(new_n682), .B2(new_n683), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n746), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n753), .A2(KEYINPUT42), .A3(new_n712), .A4(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n751), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(KEYINPUT109), .B(G131), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n757), .B(new_n758), .ZN(G33));
  NAND4_X1  g573(.A1(new_n755), .A2(new_n557), .A3(new_n607), .A4(new_n679), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G134), .ZN(G36));
  NAND2_X1  g575(.A1(new_n702), .A2(new_n708), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(KEYINPUT43), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT43), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n702), .A2(new_n764), .A3(new_n708), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n665), .A2(new_n615), .A3(new_n763), .A4(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT44), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT111), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n766), .A2(KEYINPUT111), .A3(new_n767), .ZN(new_n771));
  OR2_X1    g585(.A1(new_n766), .A2(new_n767), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n770), .A2(new_n748), .A3(new_n771), .A4(new_n772), .ZN(new_n773));
  OR2_X1    g587(.A1(new_n773), .A2(KEYINPUT112), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(KEYINPUT112), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n616), .B1(new_n618), .B2(new_n405), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT45), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n334), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n410), .A2(KEYINPUT45), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n335), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g594(.A(KEYINPUT110), .B1(new_n780), .B2(KEYINPUT46), .ZN(new_n781));
  OR3_X1    g595(.A1(new_n780), .A2(KEYINPUT110), .A3(KEYINPUT46), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n780), .A2(KEYINPUT46), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n781), .A2(new_n417), .A3(new_n782), .A4(new_n783), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n784), .A2(new_n622), .A3(new_n697), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n774), .A2(new_n775), .A3(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G137), .ZN(G39));
  NOR4_X1   g601(.A1(new_n750), .A2(new_n557), .A3(new_n607), .A4(new_n754), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n784), .A2(KEYINPUT47), .A3(new_n622), .ZN(new_n789));
  AOI21_X1  g603(.A(KEYINPUT47), .B1(new_n784), .B2(new_n622), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G140), .ZN(G42));
  NAND3_X1  g606(.A1(new_n655), .A2(new_n661), .A3(new_n709), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n670), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n794), .B(new_n731), .C1(new_n694), .C2(new_n695), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n671), .B(new_n665), .C1(new_n712), .C2(new_n679), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n795), .A2(new_n796), .A3(new_n740), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT116), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n795), .A2(new_n796), .A3(new_n740), .A4(KEYINPUT116), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT52), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n702), .A2(new_n728), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n491), .A2(new_n804), .A3(new_n329), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n624), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n639), .A2(new_n330), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n808), .A2(new_n684), .A3(new_n809), .A4(new_n490), .ZN(new_n810));
  OAI21_X1  g624(.A(KEYINPUT114), .B1(new_n491), .B2(new_n807), .ZN(new_n811));
  INV_X1    g625(.A(new_n615), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n603), .A2(new_n623), .A3(new_n606), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n810), .A2(new_n811), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n806), .A2(new_n814), .A3(new_n666), .ZN(new_n815));
  INV_X1    g629(.A(new_n492), .ZN(new_n816));
  INV_X1    g630(.A(new_n610), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n816), .B1(new_n817), .B2(new_n608), .ZN(new_n818));
  OAI21_X1  g632(.A(KEYINPUT115), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  AOI22_X1  g633(.A1(new_n624), .A2(new_n805), .B1(new_n652), .B2(new_n665), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT115), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n611), .A2(new_n820), .A3(new_n821), .A4(new_n814), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n755), .A2(new_n665), .A3(new_n712), .A4(new_n736), .ZN(new_n824));
  NOR4_X1   g638(.A1(new_n623), .A2(new_n646), .A3(new_n728), .A4(new_n678), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n665), .A2(new_n825), .A3(new_n557), .A4(new_n748), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n824), .A2(new_n760), .A3(new_n826), .ZN(new_n827));
  AND4_X1   g641(.A1(new_n719), .A2(new_n725), .A3(new_n737), .A4(new_n722), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n757), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n799), .A2(KEYINPUT52), .A3(new_n800), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n803), .A2(new_n823), .A3(new_n830), .A4(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT53), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT54), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n829), .B1(new_n822), .B2(new_n819), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n797), .A2(KEYINPUT52), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n836), .A2(KEYINPUT53), .A3(new_n803), .A4(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n834), .A2(new_n835), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(KEYINPUT117), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n836), .A2(KEYINPUT53), .A3(new_n803), .A4(new_n831), .ZN(new_n841));
  AND4_X1   g655(.A1(new_n803), .A2(new_n823), .A3(new_n830), .A4(new_n837), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n841), .B1(new_n842), .B2(KEYINPUT53), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(KEYINPUT54), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT117), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n834), .A2(new_n845), .A3(new_n838), .A4(new_n835), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n840), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n672), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n763), .A2(new_n765), .A3(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT118), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n849), .B(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n748), .A2(new_n718), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n852), .B(KEYINPUT120), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n854), .A2(new_n665), .A3(new_n736), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n613), .A2(new_n325), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n696), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(new_n853), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n701), .A2(new_n708), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(KEYINPUT121), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT121), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n857), .A2(new_n862), .A3(new_n853), .A4(new_n859), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n855), .A2(new_n861), .A3(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT122), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n855), .A2(new_n861), .A3(KEYINPUT122), .A4(new_n863), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT119), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n736), .A2(new_n607), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n851), .A2(new_n870), .A3(new_n748), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n789), .A2(new_n790), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n717), .A2(new_n417), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(new_n333), .ZN(new_n874));
  AOI22_X1  g688(.A1(new_n869), .A2(new_n871), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n851), .A2(KEYINPUT119), .A3(new_n870), .A4(new_n748), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n686), .A2(new_n703), .A3(new_n718), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n877), .A2(new_n851), .A3(new_n870), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT50), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n877), .A2(KEYINPUT50), .A3(new_n870), .A4(new_n851), .ZN(new_n881));
  AOI22_X1  g695(.A1(new_n875), .A2(new_n876), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n868), .A2(KEYINPUT51), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n854), .A2(new_n753), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(KEYINPUT48), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n851), .A2(new_n739), .A3(new_n870), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n322), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n858), .A2(new_n640), .ZN(new_n888));
  OR3_X1    g702(.A1(new_n887), .A2(new_n888), .A3(KEYINPUT123), .ZN(new_n889));
  OAI21_X1  g703(.A(KEYINPUT123), .B1(new_n887), .B2(new_n888), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n885), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n864), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n882), .A2(new_n892), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n883), .B(new_n891), .C1(KEYINPUT51), .C2(new_n893), .ZN(new_n894));
  OAI22_X1  g708(.A1(new_n847), .A2(new_n894), .B1(G952), .B2(G953), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n873), .B(KEYINPUT49), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n686), .A2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT113), .ZN(new_n898));
  OR4_X1    g712(.A1(new_n613), .A2(new_n703), .A3(new_n333), .A4(new_n762), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n900), .B(new_n696), .C1(new_n898), .C2(new_n899), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n895), .A2(new_n901), .ZN(G75));
  NAND2_X1  g716(.A1(new_n834), .A2(new_n838), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n903), .A2(G902), .A3(new_n421), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT56), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n456), .A2(new_n457), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(new_n426), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT55), .ZN(new_n908));
  AND3_X1   g722(.A1(new_n904), .A2(new_n905), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n908), .B1(new_n904), .B2(new_n905), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n189), .A2(G952), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(G51));
  XNOR2_X1  g726(.A(new_n335), .B(KEYINPUT57), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n834), .A2(new_n835), .A3(new_n838), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n835), .B1(new_n834), .B2(new_n838), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n916), .B1(new_n416), .B2(new_n415), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n903), .A2(G902), .A3(new_n779), .A4(new_n778), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n911), .B1(new_n917), .B2(new_n918), .ZN(G54));
  INV_X1    g733(.A(KEYINPUT124), .ZN(new_n920));
  INV_X1    g734(.A(new_n911), .ZN(new_n921));
  NAND2_X1  g735(.A1(KEYINPUT58), .A2(G475), .ZN(new_n922));
  AOI211_X1 g736(.A(new_n187), .B(new_n922), .C1(new_n834), .C2(new_n838), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n921), .B1(new_n923), .B2(new_n273), .ZN(new_n924));
  INV_X1    g738(.A(new_n922), .ZN(new_n925));
  AND4_X1   g739(.A1(G902), .A2(new_n903), .A3(new_n273), .A4(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n920), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n903), .A2(G902), .A3(new_n925), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n928), .A2(new_n237), .A3(new_n260), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n923), .A2(new_n273), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n929), .A2(new_n930), .A3(KEYINPUT124), .A4(new_n921), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n927), .A2(new_n931), .ZN(G60));
  NOR2_X1   g746(.A1(new_n634), .A2(new_n637), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(G478), .A2(G902), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT59), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n934), .B1(new_n847), .B2(new_n936), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n934), .B(new_n936), .C1(new_n914), .C2(new_n915), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n921), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n937), .A2(new_n939), .ZN(G63));
  NAND2_X1  g754(.A1(G217), .A2(G902), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT60), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n903), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n911), .B1(new_n944), .B2(new_n604), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n945), .B(KEYINPUT61), .C1(new_n659), .C2(new_n944), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT61), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n944), .A2(new_n659), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n942), .B1(new_n834), .B2(new_n838), .ZN(new_n949));
  INV_X1    g763(.A(new_n604), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n921), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n947), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n946), .A2(new_n952), .ZN(G66));
  INV_X1    g767(.A(G224), .ZN(new_n954));
  OAI21_X1  g768(.A(G953), .B1(new_n327), .B2(new_n954), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n823), .A2(new_n828), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n955), .B1(new_n956), .B2(G953), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n906), .B1(G898), .B2(new_n189), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n957), .B(new_n958), .ZN(G69));
  AOI21_X1  g773(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n796), .A2(new_n740), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT125), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n962), .B(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n760), .ZN(new_n965));
  NOR4_X1   g779(.A1(new_n752), .A2(new_n631), .A3(new_n730), .A4(new_n729), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n965), .B1(new_n785), .B2(new_n966), .ZN(new_n967));
  AND4_X1   g781(.A1(new_n757), .A2(new_n964), .A3(new_n791), .A4(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n786), .A2(new_n189), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n500), .B1(new_n494), .B2(new_n504), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(new_n248), .Z(new_n971));
  AOI21_X1  g785(.A(new_n971), .B1(G900), .B2(G953), .ZN(new_n972));
  AOI21_X1  g786(.A(KEYINPUT127), .B1(new_n969), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n964), .A2(new_n706), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT62), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n974), .B(new_n975), .ZN(new_n976));
  AOI211_X1 g790(.A(new_n698), .B(new_n754), .C1(new_n640), .C2(new_n804), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n977), .B1(new_n609), .B2(new_n610), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n791), .B1(KEYINPUT126), .B2(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n979), .B1(KEYINPUT126), .B2(new_n978), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n976), .A2(new_n980), .A3(new_n786), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n981), .A2(new_n189), .ZN(new_n982));
  INV_X1    g796(.A(new_n971), .ZN(new_n983));
  OAI211_X1 g797(.A(new_n961), .B(new_n973), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n983), .B1(new_n981), .B2(new_n189), .ZN(new_n985));
  INV_X1    g799(.A(new_n973), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n960), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n984), .A2(new_n987), .ZN(G72));
  NAND2_X1  g802(.A1(G472), .A2(G902), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT63), .Z(new_n990));
  AND4_X1   g804(.A1(new_n516), .A2(new_n843), .A3(new_n688), .A4(new_n990), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n976), .A2(new_n980), .A3(new_n786), .A4(new_n956), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n688), .B1(new_n992), .B2(new_n990), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n786), .A2(new_n956), .A3(new_n968), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n516), .B1(new_n994), .B2(new_n990), .ZN(new_n995));
  NOR4_X1   g809(.A1(new_n991), .A2(new_n993), .A3(new_n911), .A4(new_n995), .ZN(G57));
endmodule


