//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 0 1 1 0 1 0 1 0 0 1 0 1 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 0 1 1 1 0 1 0 0 0 0 0 1 1 1 1 0 0 1 1 0 1 0 1 0 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:09 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n537, new_n538, new_n539, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n550, new_n551, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n560, new_n561, new_n562,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n589, new_n590, new_n591, new_n592, new_n595, new_n597, new_n598,
    new_n599, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1108;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT65), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  NAND2_X1  g029(.A1(new_n451), .A2(G2106), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n452), .A2(G567), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT66), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  NAND3_X1  g035(.A1(new_n460), .A2(G101), .A3(G2104), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n461), .B(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G137), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(new_n460), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n463), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  AOI22_X1  g042(.A1(new_n465), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(new_n460), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n467), .A2(new_n469), .ZN(G160));
  NAND2_X1  g045(.A1(new_n465), .A2(G2105), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G124), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n460), .A2(G112), .ZN(new_n474));
  OAI21_X1  g049(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n466), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n476), .B1(G136), .B2(new_n477), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT68), .ZN(G162));
  INV_X1    g054(.A(KEYINPUT71), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n460), .A2(G138), .ZN(new_n481));
  OR2_X1    g056(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n482));
  NAND2_X1  g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n480), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT70), .ZN(new_n487));
  OAI21_X1  g062(.A(KEYINPUT4), .B1(new_n484), .B2(new_n487), .ZN(new_n488));
  AND2_X1   g063(.A1(new_n460), .A2(G138), .ZN(new_n489));
  NOR2_X1   g064(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n490));
  INV_X1    g065(.A(new_n483), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n489), .B(new_n487), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n486), .B1(new_n488), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n465), .A2(new_n489), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT70), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n496), .A2(new_n480), .A3(KEYINPUT4), .A4(new_n492), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n498), .B1(new_n499), .B2(G2105), .ZN(new_n500));
  OAI211_X1 g075(.A(G126), .B(G2105), .C1(new_n491), .C2(new_n490), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n465), .A2(KEYINPUT69), .A3(G126), .A4(G2105), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n500), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n494), .A2(new_n497), .A3(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  AND2_X1   g082(.A1(G75), .A2(G543), .ZN(new_n508));
  OAI21_X1  g083(.A(KEYINPUT5), .B1(KEYINPUT72), .B2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n509), .B1(KEYINPUT73), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT73), .ZN(new_n512));
  NAND4_X1  g087(.A1(new_n512), .A2(KEYINPUT72), .A3(KEYINPUT5), .A4(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n508), .B1(new_n514), .B2(G62), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT74), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  OR3_X1    g092(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n516), .B1(new_n515), .B2(new_n517), .ZN(new_n519));
  AND2_X1   g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n522), .B1(new_n511), .B2(new_n513), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n522), .A2(new_n510), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n523), .A2(G88), .B1(new_n524), .B2(G50), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n518), .A2(new_n519), .A3(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  XOR2_X1   g102(.A(KEYINPUT75), .B(KEYINPUT7), .Z(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n528), .B(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n524), .A2(G51), .ZN(new_n532));
  AND3_X1   g107(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n523), .A2(G89), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  AOI22_X1  g111(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n537), .A2(new_n517), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n523), .A2(G90), .B1(new_n524), .B2(G52), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  AOI22_X1  g116(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(new_n517), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n523), .A2(G81), .B1(new_n524), .B2(G43), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT76), .ZN(G153));
  NAND4_X1  g123(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(G188));
  NAND2_X1  g127(.A1(new_n524), .A2(G53), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(KEYINPUT9), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT9), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n524), .A2(new_n555), .A3(G53), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n554), .A2(new_n556), .B1(G91), .B2(new_n523), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n514), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n517), .B2(new_n558), .ZN(G299));
  NAND2_X1  g134(.A1(new_n523), .A2(G87), .ZN(new_n560));
  OAI21_X1  g135(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n524), .A2(G49), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(G288));
  AOI22_X1  g138(.A1(new_n523), .A2(G86), .B1(new_n524), .B2(G48), .ZN(new_n564));
  INV_X1    g139(.A(G61), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n565), .B1(new_n511), .B2(new_n513), .ZN(new_n566));
  NAND2_X1  g141(.A1(G73), .A2(G543), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT77), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n564), .A2(new_n569), .ZN(G305));
  NAND2_X1  g145(.A1(new_n523), .A2(G85), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n524), .A2(G47), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  XOR2_X1   g148(.A(new_n573), .B(KEYINPUT79), .Z(new_n574));
  AOI22_X1  g149(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n517), .B1(new_n576), .B2(KEYINPUT78), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n577), .B1(KEYINPUT78), .B2(new_n576), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n574), .A2(new_n578), .ZN(G290));
  NAND2_X1  g154(.A1(G301), .A2(G868), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n523), .A2(G92), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n581), .B(KEYINPUT10), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n524), .A2(G54), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n514), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n584), .B2(new_n517), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n580), .B1(new_n586), .B2(G868), .ZN(G284));
  OAI21_X1  g162(.A(new_n580), .B1(new_n586), .B2(G868), .ZN(G321));
  INV_X1    g163(.A(G868), .ZN(new_n589));
  OR3_X1    g164(.A1(G168), .A2(KEYINPUT80), .A3(new_n589), .ZN(new_n590));
  OAI21_X1  g165(.A(KEYINPUT80), .B1(G168), .B2(new_n589), .ZN(new_n591));
  NAND2_X1  g166(.A1(G299), .A2(new_n589), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(G297));
  NAND3_X1  g168(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(G280));
  INV_X1    g169(.A(G559), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n586), .B1(new_n595), .B2(G860), .ZN(G148));
  NAND2_X1  g171(.A1(new_n545), .A2(new_n589), .ZN(new_n597));
  INV_X1    g172(.A(new_n586), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n598), .A2(G559), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n597), .B1(new_n599), .B2(new_n589), .ZN(G323));
  XNOR2_X1  g175(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g176(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n602));
  INV_X1    g177(.A(G111), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(G2105), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n477), .A2(G135), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT82), .ZN(new_n606));
  AOI211_X1 g181(.A(new_n604), .B(new_n606), .C1(G123), .C2(new_n472), .ZN(new_n607));
  INV_X1    g182(.A(G2096), .ZN(new_n608));
  XOR2_X1   g183(.A(KEYINPUT81), .B(G2100), .Z(new_n609));
  AND2_X1   g184(.A1(new_n460), .A2(G2104), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n465), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT12), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT13), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n607), .A2(new_n608), .B1(new_n609), .B2(new_n613), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n613), .A2(new_n609), .ZN(new_n615));
  OAI211_X1 g190(.A(new_n614), .B(new_n615), .C1(new_n608), .C2(new_n607), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT83), .Z(G156));
  XNOR2_X1  g192(.A(G2427), .B(G2438), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(G2430), .ZN(new_n619));
  XNOR2_X1  g194(.A(KEYINPUT15), .B(G2435), .ZN(new_n620));
  OR2_X1    g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n619), .A2(new_n620), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n621), .A2(new_n622), .A3(KEYINPUT14), .ZN(new_n623));
  XOR2_X1   g198(.A(G1341), .B(G1348), .Z(new_n624));
  XNOR2_X1  g199(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n623), .B(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(G2451), .B(G2454), .Z(new_n628));
  XNOR2_X1  g203(.A(G2443), .B(G2446), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n627), .A2(new_n630), .ZN(new_n632));
  AND3_X1   g207(.A1(new_n631), .A2(G14), .A3(new_n632), .ZN(G401));
  INV_X1    g208(.A(KEYINPUT18), .ZN(new_n634));
  XOR2_X1   g209(.A(G2084), .B(G2090), .Z(new_n635));
  XNOR2_X1  g210(.A(G2067), .B(G2678), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(KEYINPUT17), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n635), .A2(new_n636), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n634), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2100), .ZN(new_n641));
  XOR2_X1   g216(.A(G2072), .B(G2078), .Z(new_n642));
  AOI21_X1  g217(.A(new_n642), .B1(new_n637), .B2(KEYINPUT18), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2096), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n641), .B(new_n644), .ZN(G227));
  XOR2_X1   g220(.A(G1971), .B(G1976), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT19), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1956), .B(G2474), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1961), .B(G1966), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AND2_X1   g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  NOR3_X1   g226(.A1(new_n647), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n647), .A2(new_n650), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT20), .Z(new_n654));
  AOI211_X1 g229(.A(new_n652), .B(new_n654), .C1(new_n647), .C2(new_n651), .ZN(new_n655));
  INV_X1    g230(.A(G1981), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G1986), .ZN(new_n658));
  XOR2_X1   g233(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT85), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n658), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1991), .B(G1996), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(G229));
  INV_X1    g238(.A(G29), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(G26), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT28), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n472), .A2(G128), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n477), .A2(G140), .ZN(new_n668));
  OR2_X1    g243(.A1(G104), .A2(G2105), .ZN(new_n669));
  OAI211_X1 g244(.A(new_n669), .B(G2104), .C1(G116), .C2(new_n460), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n667), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n666), .B1(new_n672), .B2(new_n664), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(G2067), .ZN(new_n674));
  XOR2_X1   g249(.A(KEYINPUT31), .B(G11), .Z(new_n675));
  AND2_X1   g250(.A1(new_n607), .A2(G29), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT92), .B(G28), .ZN(new_n677));
  OR2_X1    g252(.A1(new_n677), .A2(KEYINPUT30), .ZN(new_n678));
  AOI21_X1  g253(.A(G29), .B1(new_n677), .B2(KEYINPUT30), .ZN(new_n679));
  AOI211_X1 g254(.A(new_n675), .B(new_n676), .C1(new_n678), .C2(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(G2072), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT25), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n465), .A2(G127), .ZN(new_n684));
  NAND2_X1  g259(.A1(G115), .A2(G2104), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n460), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  AOI211_X1 g261(.A(new_n683), .B(new_n686), .C1(G139), .C2(new_n477), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(G29), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(G29), .B2(G33), .ZN(new_n689));
  INV_X1    g264(.A(G16), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G21), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(G168), .B2(new_n690), .ZN(new_n692));
  OAI221_X1 g267(.A(new_n680), .B1(new_n681), .B2(new_n689), .C1(new_n692), .C2(G1966), .ZN(new_n693));
  AOI211_X1 g268(.A(new_n674), .B(new_n693), .C1(G1966), .C2(new_n692), .ZN(new_n694));
  INV_X1    g269(.A(G34), .ZN(new_n695));
  AOI21_X1  g270(.A(G29), .B1(new_n695), .B2(KEYINPUT24), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(KEYINPUT24), .B2(new_n695), .ZN(new_n697));
  INV_X1    g272(.A(G160), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n697), .B1(new_n698), .B2(new_n664), .ZN(new_n699));
  INV_X1    g274(.A(G2084), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  AND2_X1   g276(.A1(new_n689), .A2(new_n681), .ZN(new_n702));
  INV_X1    g277(.A(G1341), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n546), .A2(G16), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G16), .B2(G19), .ZN(new_n705));
  AOI211_X1 g280(.A(new_n701), .B(new_n702), .C1(new_n703), .C2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n690), .A2(G20), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT95), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT23), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(G299), .B2(G16), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT96), .B(G1956), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  NOR2_X1   g287(.A1(G4), .A2(G16), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT90), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(new_n598), .B2(new_n690), .ZN(new_n715));
  INV_X1    g290(.A(G1348), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g292(.A1(new_n694), .A2(new_n706), .A3(new_n712), .A4(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n664), .A2(G35), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G162), .B2(new_n664), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT29), .Z(new_n721));
  INV_X1    g296(.A(G2090), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n721), .A2(new_n722), .ZN(new_n724));
  NOR2_X1   g299(.A1(G5), .A2(G16), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT93), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G301), .B2(new_n690), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT94), .Z(new_n728));
  INV_X1    g303(.A(G1961), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n723), .A2(new_n724), .A3(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n715), .A2(new_n716), .ZN(new_n732));
  INV_X1    g307(.A(G2078), .ZN(new_n733));
  NAND2_X1  g308(.A1(G164), .A2(G29), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G27), .B2(G29), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n732), .B1(new_n733), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(new_n733), .B2(new_n735), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n664), .A2(G32), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n477), .A2(G141), .B1(G105), .B2(new_n610), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n472), .A2(G129), .ZN(new_n740));
  NAND3_X1  g315(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT26), .Z(new_n742));
  NAND3_X1  g317(.A1(new_n739), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n743), .A2(KEYINPUT91), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(KEYINPUT91), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n738), .B1(new_n747), .B2(new_n664), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT27), .B(G1996), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  OAI221_X1 g325(.A(new_n750), .B1(new_n703), .B2(new_n705), .C1(new_n729), .C2(new_n728), .ZN(new_n751));
  NOR4_X1   g326(.A1(new_n718), .A2(new_n731), .A3(new_n737), .A4(new_n751), .ZN(new_n752));
  MUX2_X1   g327(.A(G6), .B(G305), .S(G16), .Z(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT32), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G1981), .ZN(new_n755));
  NAND2_X1  g330(.A1(G166), .A2(G16), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G16), .B2(G22), .ZN(new_n757));
  INV_X1    g332(.A(G1971), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n757), .A2(new_n758), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n690), .A2(G23), .ZN(new_n761));
  INV_X1    g336(.A(G288), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n761), .B1(new_n762), .B2(new_n690), .ZN(new_n763));
  XOR2_X1   g338(.A(KEYINPUT33), .B(G1976), .Z(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NOR4_X1   g340(.A1(new_n755), .A2(new_n759), .A3(new_n760), .A4(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT34), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n690), .A2(G24), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G290), .B2(G16), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT87), .B(G1986), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n770), .A2(new_n771), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n664), .A2(G25), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n472), .A2(G119), .B1(new_n477), .B2(G131), .ZN(new_n775));
  OR2_X1    g350(.A1(G95), .A2(G2105), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n776), .B(G2104), .C1(G107), .C2(new_n460), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT86), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n774), .B1(new_n779), .B2(new_n664), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT35), .B(G1991), .Z(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n768), .A2(new_n772), .A3(new_n773), .A4(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT88), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n783), .A2(new_n784), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n766), .A2(new_n767), .ZN(new_n787));
  NOR3_X1   g362(.A1(new_n785), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  XOR2_X1   g363(.A(KEYINPUT89), .B(KEYINPUT36), .Z(new_n789));
  OAI21_X1  g364(.A(new_n752), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT36), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n791), .A2(KEYINPUT89), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n788), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n790), .A2(new_n793), .ZN(G311));
  INV_X1    g369(.A(G311), .ZN(G150));
  AOI22_X1  g370(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n796));
  OR3_X1    g371(.A1(new_n796), .A2(KEYINPUT97), .A3(new_n517), .ZN(new_n797));
  OAI21_X1  g372(.A(KEYINPUT97), .B1(new_n796), .B2(new_n517), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT98), .B(G93), .ZN(new_n799));
  AOI22_X1  g374(.A1(new_n523), .A2(new_n799), .B1(new_n524), .B2(G55), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n797), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT99), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n801), .B1(new_n802), .B2(new_n546), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n545), .A2(KEYINPUT99), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n586), .A2(G559), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n807), .B(new_n808), .Z(new_n809));
  AND2_X1   g384(.A1(new_n809), .A2(KEYINPUT39), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n809), .A2(KEYINPUT39), .ZN(new_n811));
  NOR3_X1   g386(.A1(new_n810), .A2(new_n811), .A3(G860), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n801), .A2(G860), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT37), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n812), .A2(new_n814), .ZN(G145));
  XNOR2_X1  g390(.A(new_n746), .B(new_n672), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n816), .A2(new_n506), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n687), .A2(KEYINPUT101), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n816), .A2(new_n506), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n817), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n779), .B(new_n612), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n687), .A2(KEYINPUT101), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n472), .A2(G130), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n460), .A2(G118), .ZN(new_n825));
  OAI21_X1  g400(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(G142), .B2(new_n477), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n823), .B(new_n828), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n822), .B(new_n829), .Z(new_n830));
  XNOR2_X1  g405(.A(G162), .B(new_n698), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(new_n607), .ZN(new_n832));
  AOI21_X1  g407(.A(G37), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(new_n832), .B2(new_n830), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g410(.A1(new_n801), .A2(G868), .ZN(new_n836));
  XNOR2_X1  g411(.A(G290), .B(G288), .ZN(new_n837));
  XNOR2_X1  g412(.A(G303), .B(G305), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT102), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n839), .B1(new_n840), .B2(KEYINPUT42), .ZN(new_n841));
  XNOR2_X1  g416(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n841), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n805), .B(new_n599), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n586), .B(G299), .Z(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(KEYINPUT41), .Z(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n845), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n847), .B1(new_n848), .B2(new_n844), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n843), .B1(KEYINPUT103), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n849), .A2(KEYINPUT103), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n850), .B(new_n851), .Z(new_n852));
  AOI21_X1  g427(.A(new_n836), .B1(new_n852), .B2(G868), .ZN(G295));
  AOI21_X1  g428(.A(new_n836), .B1(new_n852), .B2(G868), .ZN(G331));
  XNOR2_X1  g429(.A(G171), .B(G286), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n805), .B(new_n855), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n856), .A2(new_n846), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n848), .ZN(new_n858));
  AND3_X1   g433(.A1(new_n857), .A2(new_n839), .A3(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT104), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(G37), .B1(new_n859), .B2(new_n860), .ZN(new_n862));
  AND2_X1   g437(.A1(new_n857), .A2(new_n858), .ZN(new_n863));
  OAI211_X1 g438(.A(new_n861), .B(new_n862), .C1(new_n839), .C2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(KEYINPUT43), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT105), .ZN(new_n866));
  AND2_X1   g441(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n858), .A2(new_n866), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n868), .A2(new_n839), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n861), .B(new_n862), .C1(new_n867), .C2(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n865), .B1(new_n870), .B2(KEYINPUT43), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT43), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n864), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n873), .B1(new_n870), .B2(new_n872), .ZN(new_n874));
  MUX2_X1   g449(.A(new_n871), .B(new_n874), .S(KEYINPUT44), .Z(G397));
  INV_X1    g450(.A(G1996), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n747), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(G2067), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n671), .B(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n746), .A2(G1996), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n877), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  OR2_X1    g457(.A1(new_n779), .A2(new_n781), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n779), .A2(new_n781), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(KEYINPUT106), .B(G1384), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n506), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT45), .ZN(new_n888));
  INV_X1    g463(.A(G40), .ZN(new_n889));
  NOR3_X1   g464(.A1(new_n467), .A2(new_n469), .A3(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n887), .A2(new_n888), .A3(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(G290), .A2(G1986), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(G290), .A2(G1986), .ZN(new_n895));
  OR3_X1    g470(.A1(new_n894), .A2(KEYINPUT107), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n891), .B1(new_n894), .B2(KEYINPUT107), .ZN(new_n897));
  AOI22_X1  g472(.A1(new_n885), .A2(new_n892), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT50), .ZN(new_n899));
  INV_X1    g474(.A(G1384), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n506), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n899), .B1(new_n506), .B2(new_n900), .ZN(new_n902));
  INV_X1    g477(.A(new_n890), .ZN(new_n903));
  NOR3_X1   g478(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(new_n722), .ZN(new_n905));
  AOI21_X1  g480(.A(KEYINPUT45), .B1(new_n506), .B2(new_n900), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n506), .A2(KEYINPUT45), .A3(new_n886), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(KEYINPUT108), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT108), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n506), .A2(new_n909), .A3(KEYINPUT45), .A4(new_n886), .ZN(new_n910));
  AOI211_X1 g485(.A(new_n903), .B(new_n906), .C1(new_n908), .C2(new_n910), .ZN(new_n911));
  OAI211_X1 g486(.A(KEYINPUT115), .B(new_n905), .C1(new_n911), .C2(G1971), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT115), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n908), .A2(new_n910), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n506), .A2(new_n900), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n903), .B1(new_n915), .B2(new_n888), .ZN(new_n916));
  AOI21_X1  g491(.A(G1971), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(KEYINPUT50), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n506), .A2(new_n899), .A3(new_n900), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(new_n890), .A3(new_n919), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n920), .A2(G2090), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n913), .B1(new_n917), .B2(new_n921), .ZN(new_n922));
  XOR2_X1   g497(.A(KEYINPUT110), .B(G8), .Z(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n912), .A2(new_n922), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(G303), .A2(G8), .ZN(new_n926));
  XNOR2_X1  g501(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n926), .B(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n925), .A2(new_n930), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n929), .B(G8), .C1(new_n917), .C2(new_n921), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n506), .A2(new_n890), .A3(new_n900), .ZN(new_n934));
  INV_X1    g509(.A(G1976), .ZN(new_n935));
  OAI211_X1 g510(.A(new_n934), .B(new_n924), .C1(new_n935), .C2(G288), .ZN(new_n936));
  NAND2_X1  g511(.A1(KEYINPUT111), .A2(KEYINPUT52), .ZN(new_n937));
  NOR2_X1   g512(.A1(KEYINPUT52), .A2(G1976), .ZN(new_n938));
  AOI22_X1  g513(.A1(new_n936), .A2(new_n937), .B1(G288), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n934), .A2(new_n924), .ZN(new_n940));
  NOR2_X1   g515(.A1(G288), .A2(new_n935), .ZN(new_n941));
  OR3_X1    g516(.A1(new_n940), .A2(new_n941), .A3(new_n937), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n939), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(G305), .A2(KEYINPUT49), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT49), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n564), .A2(new_n569), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n656), .B1(new_n569), .B2(KEYINPUT112), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n944), .A2(new_n948), .A3(new_n946), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(new_n940), .ZN(new_n953));
  AOI21_X1  g528(.A(KEYINPUT113), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  AND4_X1   g529(.A1(KEYINPUT113), .A2(new_n953), .A3(new_n951), .A4(new_n950), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n943), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n933), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(G1966), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT116), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n506), .A2(new_n959), .A3(KEYINPUT45), .A4(new_n900), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n506), .A2(KEYINPUT45), .A3(new_n900), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT116), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n916), .A2(new_n960), .A3(new_n962), .ZN(new_n963));
  AOI22_X1  g538(.A1(new_n958), .A2(new_n963), .B1(new_n904), .B2(new_n700), .ZN(new_n964));
  NOR3_X1   g539(.A1(new_n964), .A2(G286), .A3(new_n923), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n931), .A2(new_n957), .A3(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT63), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT117), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n966), .A2(KEYINPUT117), .A3(new_n967), .ZN(new_n971));
  OAI21_X1  g546(.A(G8), .B1(new_n917), .B2(new_n921), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(new_n930), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n957), .A2(KEYINPUT63), .A3(new_n965), .A4(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n970), .A2(new_n971), .A3(new_n974), .ZN(new_n975));
  XNOR2_X1  g550(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n976), .B(G2072), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n914), .A2(new_n916), .A3(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT118), .ZN(new_n979));
  AND3_X1   g554(.A1(G299), .A2(new_n979), .A3(KEYINPUT57), .ZN(new_n980));
  AOI21_X1  g555(.A(KEYINPUT57), .B1(G299), .B2(new_n979), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G1956), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n920), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n978), .A2(new_n982), .A3(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n902), .A2(new_n903), .ZN(new_n987));
  AOI21_X1  g562(.A(G1348), .B1(new_n987), .B2(new_n919), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n934), .A2(G2067), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n586), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n986), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n982), .B1(new_n978), .B2(new_n984), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n989), .ZN(new_n994));
  OAI211_X1 g569(.A(new_n598), .B(new_n994), .C1(new_n904), .C2(G1348), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n990), .A2(new_n995), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n988), .A2(new_n989), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n598), .A2(KEYINPUT60), .ZN(new_n998));
  AOI22_X1  g573(.A1(new_n996), .A2(KEYINPUT60), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT61), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n1000), .B1(new_n986), .B2(KEYINPUT120), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT59), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n914), .A2(new_n916), .ZN(new_n1003));
  INV_X1    g578(.A(new_n934), .ZN(new_n1004));
  XNOR2_X1  g579(.A(KEYINPUT58), .B(G1341), .ZN(new_n1005));
  OAI22_X1  g580(.A1(new_n1003), .A2(G1996), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1002), .B1(new_n1006), .B2(new_n546), .ZN(new_n1007));
  AND3_X1   g582(.A1(new_n1006), .A2(new_n1002), .A3(new_n546), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n999), .B(new_n1001), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n992), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1010), .A2(KEYINPUT121), .A3(KEYINPUT61), .A4(new_n985), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT121), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n985), .A2(KEYINPUT61), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1012), .B1(new_n1013), .B2(new_n992), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1011), .A2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n993), .B1(new_n1009), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G8), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n963), .A2(new_n958), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n904), .A2(new_n700), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1017), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(G168), .A2(new_n923), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT51), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT122), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n923), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1021), .A2(KEYINPUT51), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1023), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  OAI211_X1 g602(.A(KEYINPUT122), .B(new_n1025), .C1(new_n964), .C2(new_n923), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1022), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  OR3_X1    g604(.A1(new_n964), .A2(G168), .A3(new_n923), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT123), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1032), .B1(new_n904), .B2(G1961), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n920), .A2(KEYINPUT123), .A3(new_n729), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n733), .A2(KEYINPUT53), .ZN(new_n1035));
  AOI211_X1 g610(.A(new_n1035), .B(new_n903), .C1(new_n887), .C2(new_n888), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(new_n914), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1033), .A2(new_n1034), .A3(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n914), .A2(new_n733), .A3(new_n916), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n1040));
  AND2_X1   g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(G171), .B1(new_n1038), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT124), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n1044));
  OAI22_X1  g619(.A1(new_n963), .A2(new_n1035), .B1(new_n904), .B2(G1961), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1045), .B1(new_n1040), .B2(new_n1039), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1044), .B1(new_n1046), .B2(G301), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT124), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1048), .B(G171), .C1(new_n1038), .C2(new_n1041), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1043), .A2(new_n1047), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n931), .A2(new_n957), .ZN(new_n1051));
  OAI21_X1  g626(.A(G171), .B1(new_n1041), .B2(new_n1045), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n920), .A2(new_n729), .ZN(new_n1053));
  AOI22_X1  g628(.A1(new_n1053), .A2(new_n1032), .B1(new_n914), .B2(new_n1036), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1054), .A2(new_n1055), .A3(G301), .A4(new_n1034), .ZN(new_n1056));
  AOI21_X1  g631(.A(KEYINPUT54), .B1(new_n1052), .B2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1051), .A2(new_n1057), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1016), .A2(new_n1031), .A3(new_n1050), .A4(new_n1058), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n956), .A2(new_n932), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n935), .B(new_n762), .C1(new_n954), .C2(new_n955), .ZN(new_n1061));
  NOR2_X1   g636(.A1(G305), .A2(G1981), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT114), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n940), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1061), .A2(KEYINPUT114), .A3(new_n1063), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1060), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n975), .A2(new_n1059), .A3(KEYINPUT125), .A4(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1031), .A2(KEYINPUT62), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT62), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1029), .A2(new_n1071), .A3(new_n1030), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1052), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n931), .A2(new_n957), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  AND4_X1   g650(.A1(KEYINPUT126), .A2(new_n1070), .A3(new_n1072), .A4(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1074), .B1(new_n1031), .B2(KEYINPUT62), .ZN(new_n1077));
  AOI21_X1  g652(.A(KEYINPUT126), .B1(new_n1077), .B2(new_n1072), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1069), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1068), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1051), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1057), .ZN(new_n1083));
  AND4_X1   g658(.A1(new_n1082), .A2(new_n1031), .A3(new_n1050), .A4(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1081), .B1(new_n1084), .B2(new_n1016), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT125), .B1(new_n1085), .B2(new_n975), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n898), .B1(new_n1080), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n879), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n892), .B1(new_n746), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT46), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1090), .B1(new_n892), .B2(new_n876), .ZN(new_n1091));
  NOR3_X1   g666(.A1(new_n891), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1089), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  XOR2_X1   g668(.A(new_n1093), .B(KEYINPUT47), .Z(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT48), .B1(new_n895), .B2(new_n892), .ZN(new_n1095));
  INV_X1    g670(.A(new_n895), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT48), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n1096), .A2(new_n1097), .A3(new_n891), .ZN(new_n1098));
  AOI211_X1 g673(.A(new_n1095), .B(new_n1098), .C1(new_n885), .C2(new_n892), .ZN(new_n1099));
  OAI22_X1  g674(.A1(new_n881), .A2(new_n884), .B1(G2067), .B2(new_n671), .ZN(new_n1100));
  AOI211_X1 g675(.A(new_n1094), .B(new_n1099), .C1(new_n892), .C2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1087), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(KEYINPUT127), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT127), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1087), .A2(new_n1104), .A3(new_n1101), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1103), .A2(new_n1105), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g681(.A1(G229), .A2(new_n458), .A3(G401), .A4(G227), .ZN(new_n1108));
  NAND3_X1  g682(.A1(new_n1108), .A2(new_n871), .A3(new_n834), .ZN(G225));
  INV_X1    g683(.A(G225), .ZN(G308));
endmodule


