

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X1 U551 ( .A(n661), .Z(n675) );
  INV_X2 U552 ( .A(KEYINPUT66), .ZN(n528) );
  NOR2_X2 U553 ( .A1(n778), .A2(G1384), .ZN(n603) );
  XNOR2_X1 U554 ( .A(n649), .B(n648), .ZN(n650) );
  BUF_X1 U555 ( .A(n700), .Z(n701) );
  XNOR2_X1 U556 ( .A(n622), .B(KEYINPUT100), .ZN(n639) );
  INV_X1 U557 ( .A(n639), .ZN(n640) );
  XNOR2_X1 U558 ( .A(n607), .B(KEYINPUT27), .ZN(n608) );
  INV_X1 U559 ( .A(n742), .ZN(n694) );
  NAND2_X1 U560 ( .A1(G8), .A2(n661), .ZN(n742) );
  INV_X1 U561 ( .A(KEYINPUT23), .ZN(n520) );
  NOR2_X1 U562 ( .A1(n644), .A2(n643), .ZN(n646) );
  NOR2_X1 U563 ( .A1(n647), .A2(G299), .ZN(n644) );
  INV_X1 U564 ( .A(KEYINPUT101), .ZN(n645) );
  INV_X1 U565 ( .A(KEYINPUT28), .ZN(n648) );
  AND2_X2 U566 ( .A1(n696), .A2(n604), .ZN(n653) );
  XNOR2_X1 U567 ( .A(n530), .B(n529), .ZN(n593) );
  XNOR2_X1 U568 ( .A(n528), .B(KEYINPUT17), .ZN(n530) );
  NAND2_X1 U569 ( .A1(n731), .A2(n517), .ZN(n732) );
  XNOR2_X1 U570 ( .A(n521), .B(n520), .ZN(n524) );
  NOR2_X1 U571 ( .A1(n684), .A2(n663), .ZN(n516) );
  OR2_X1 U572 ( .A1(n730), .A2(n742), .ZN(n517) );
  AND2_X1 U573 ( .A1(n695), .A2(n694), .ZN(n518) );
  INV_X1 U574 ( .A(G8), .ZN(n663) );
  BUF_X1 U575 ( .A(n653), .Z(n655) );
  AND2_X1 U576 ( .A1(n685), .A2(n516), .ZN(n664) );
  INV_X1 U577 ( .A(G168), .ZN(n665) );
  AND2_X1 U578 ( .A1(n666), .A2(n665), .ZN(n669) );
  INV_X1 U579 ( .A(KEYINPUT31), .ZN(n670) );
  NOR2_X1 U580 ( .A1(n742), .A2(G1966), .ZN(n662) );
  XNOR2_X1 U581 ( .A(n662), .B(KEYINPUT95), .ZN(n685) );
  XNOR2_X1 U582 ( .A(n603), .B(KEYINPUT64), .ZN(n696) );
  INV_X1 U583 ( .A(G2105), .ZN(n519) );
  INV_X1 U584 ( .A(G2104), .ZN(n522) );
  AND2_X2 U585 ( .A1(n522), .A2(G2105), .ZN(n894) );
  BUF_X1 U586 ( .A(n593), .Z(n700) );
  XNOR2_X1 U587 ( .A(n618), .B(KEYINPUT15), .ZN(n975) );
  AND2_X4 U588 ( .A1(n519), .A2(G2104), .ZN(n594) );
  NAND2_X1 U589 ( .A1(n594), .A2(G101), .ZN(n521) );
  NAND2_X1 U590 ( .A1(n894), .A2(G125), .ZN(n523) );
  NAND2_X1 U591 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U592 ( .A(n525), .B(KEYINPUT65), .ZN(n527) );
  AND2_X1 U593 ( .A1(G2104), .A2(G2105), .ZN(n891) );
  NAND2_X1 U594 ( .A1(G113), .A2(n891), .ZN(n526) );
  NAND2_X1 U595 ( .A1(n527), .A2(n526), .ZN(n533) );
  NOR2_X1 U596 ( .A1(G2104), .A2(G2105), .ZN(n529) );
  NAND2_X1 U597 ( .A1(G137), .A2(n700), .ZN(n531) );
  XNOR2_X2 U598 ( .A(n531), .B(KEYINPUT67), .ZN(n532) );
  NOR2_X4 U599 ( .A1(n533), .A2(n532), .ZN(G160) );
  XOR2_X1 U600 ( .A(KEYINPUT0), .B(G543), .Z(n575) );
  INV_X1 U601 ( .A(G651), .ZN(n535) );
  NOR2_X1 U602 ( .A1(n575), .A2(n535), .ZN(n798) );
  NAND2_X1 U603 ( .A1(G78), .A2(n798), .ZN(n534) );
  XNOR2_X1 U604 ( .A(n534), .B(KEYINPUT70), .ZN(n543) );
  NOR2_X1 U605 ( .A1(G543), .A2(n535), .ZN(n536) );
  XOR2_X1 U606 ( .A(KEYINPUT1), .B(n536), .Z(n794) );
  NAND2_X1 U607 ( .A1(G65), .A2(n794), .ZN(n538) );
  NOR2_X4 U608 ( .A1(G651), .A2(n575), .ZN(n799) );
  NAND2_X1 U609 ( .A1(G53), .A2(n799), .ZN(n537) );
  NAND2_X1 U610 ( .A1(n538), .A2(n537), .ZN(n541) );
  NOR2_X1 U611 ( .A1(G651), .A2(G543), .ZN(n795) );
  NAND2_X1 U612 ( .A1(G91), .A2(n795), .ZN(n539) );
  XNOR2_X1 U613 ( .A(KEYINPUT69), .B(n539), .ZN(n540) );
  NOR2_X1 U614 ( .A1(n541), .A2(n540), .ZN(n542) );
  NAND2_X1 U615 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U616 ( .A(KEYINPUT71), .B(n544), .Z(G299) );
  NAND2_X1 U617 ( .A1(n795), .A2(G89), .ZN(n545) );
  XNOR2_X1 U618 ( .A(n545), .B(KEYINPUT4), .ZN(n547) );
  NAND2_X1 U619 ( .A1(G76), .A2(n798), .ZN(n546) );
  NAND2_X1 U620 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U621 ( .A(n548), .B(KEYINPUT5), .ZN(n553) );
  NAND2_X1 U622 ( .A1(G63), .A2(n794), .ZN(n550) );
  NAND2_X1 U623 ( .A1(G51), .A2(n799), .ZN(n549) );
  NAND2_X1 U624 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U625 ( .A(KEYINPUT6), .B(n551), .Z(n552) );
  NAND2_X1 U626 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U627 ( .A(n554), .B(KEYINPUT7), .ZN(G168) );
  XNOR2_X1 U628 ( .A(G168), .B(KEYINPUT8), .ZN(n555) );
  XNOR2_X1 U629 ( .A(n555), .B(KEYINPUT75), .ZN(G286) );
  NAND2_X1 U630 ( .A1(G52), .A2(n799), .ZN(n556) );
  XOR2_X1 U631 ( .A(KEYINPUT68), .B(n556), .Z(n563) );
  NAND2_X1 U632 ( .A1(G90), .A2(n795), .ZN(n558) );
  NAND2_X1 U633 ( .A1(G77), .A2(n798), .ZN(n557) );
  NAND2_X1 U634 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U635 ( .A(n559), .B(KEYINPUT9), .ZN(n561) );
  NAND2_X1 U636 ( .A1(G64), .A2(n794), .ZN(n560) );
  NAND2_X1 U637 ( .A1(n561), .A2(n560), .ZN(n562) );
  NOR2_X1 U638 ( .A1(n563), .A2(n562), .ZN(G171) );
  NAND2_X1 U639 ( .A1(n794), .A2(G62), .ZN(n564) );
  XOR2_X1 U640 ( .A(KEYINPUT81), .B(n564), .Z(n566) );
  NAND2_X1 U641 ( .A1(n799), .A2(G50), .ZN(n565) );
  NAND2_X1 U642 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U643 ( .A(KEYINPUT82), .B(n567), .Z(n571) );
  NAND2_X1 U644 ( .A1(G88), .A2(n795), .ZN(n569) );
  NAND2_X1 U645 ( .A1(G75), .A2(n798), .ZN(n568) );
  AND2_X1 U646 ( .A1(n569), .A2(n568), .ZN(n570) );
  NAND2_X1 U647 ( .A1(n571), .A2(n570), .ZN(G303) );
  NAND2_X1 U648 ( .A1(G49), .A2(n799), .ZN(n573) );
  NAND2_X1 U649 ( .A1(G74), .A2(G651), .ZN(n572) );
  NAND2_X1 U650 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X1 U651 ( .A1(n794), .A2(n574), .ZN(n577) );
  NAND2_X1 U652 ( .A1(n575), .A2(G87), .ZN(n576) );
  NAND2_X1 U653 ( .A1(n577), .A2(n576), .ZN(G288) );
  NAND2_X1 U654 ( .A1(G73), .A2(n798), .ZN(n578) );
  XNOR2_X1 U655 ( .A(n578), .B(KEYINPUT2), .ZN(n585) );
  NAND2_X1 U656 ( .A1(G61), .A2(n794), .ZN(n580) );
  NAND2_X1 U657 ( .A1(G86), .A2(n795), .ZN(n579) );
  NAND2_X1 U658 ( .A1(n580), .A2(n579), .ZN(n583) );
  NAND2_X1 U659 ( .A1(G48), .A2(n799), .ZN(n581) );
  XNOR2_X1 U660 ( .A(KEYINPUT79), .B(n581), .ZN(n582) );
  NOR2_X1 U661 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U662 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U663 ( .A(KEYINPUT80), .B(n586), .ZN(G305) );
  NAND2_X1 U664 ( .A1(G85), .A2(n795), .ZN(n588) );
  NAND2_X1 U665 ( .A1(G72), .A2(n798), .ZN(n587) );
  NAND2_X1 U666 ( .A1(n588), .A2(n587), .ZN(n592) );
  NAND2_X1 U667 ( .A1(G60), .A2(n794), .ZN(n590) );
  NAND2_X1 U668 ( .A1(G47), .A2(n799), .ZN(n589) );
  NAND2_X1 U669 ( .A1(n590), .A2(n589), .ZN(n591) );
  OR2_X1 U670 ( .A1(n592), .A2(n591), .ZN(G290) );
  NAND2_X1 U671 ( .A1(n593), .A2(G138), .ZN(n596) );
  NAND2_X1 U672 ( .A1(G102), .A2(n594), .ZN(n595) );
  NAND2_X1 U673 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U674 ( .A(n597), .B(KEYINPUT90), .ZN(n602) );
  NAND2_X1 U675 ( .A1(G126), .A2(n894), .ZN(n599) );
  NAND2_X1 U676 ( .A1(G114), .A2(n891), .ZN(n598) );
  NAND2_X1 U677 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U678 ( .A(KEYINPUT89), .B(n600), .Z(n601) );
  NOR2_X1 U679 ( .A1(n602), .A2(n601), .ZN(n778) );
  NAND2_X1 U680 ( .A1(G160), .A2(G40), .ZN(n697) );
  INV_X1 U681 ( .A(n697), .ZN(n604) );
  INV_X2 U682 ( .A(n653), .ZN(n661) );
  NAND2_X1 U683 ( .A1(G1956), .A2(n661), .ZN(n606) );
  INV_X1 U684 ( .A(KEYINPUT98), .ZN(n605) );
  XNOR2_X1 U685 ( .A(n606), .B(n605), .ZN(n609) );
  NAND2_X1 U686 ( .A1(n653), .A2(G2072), .ZN(n607) );
  NOR2_X2 U687 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X2 U688 ( .A(n610), .B(KEYINPUT99), .ZN(n647) );
  NAND2_X1 U689 ( .A1(G79), .A2(n798), .ZN(n617) );
  NAND2_X1 U690 ( .A1(G66), .A2(n794), .ZN(n612) );
  NAND2_X1 U691 ( .A1(G92), .A2(n795), .ZN(n611) );
  NAND2_X1 U692 ( .A1(n612), .A2(n611), .ZN(n615) );
  NAND2_X1 U693 ( .A1(n799), .A2(G54), .ZN(n613) );
  XOR2_X1 U694 ( .A(KEYINPUT74), .B(n613), .Z(n614) );
  NOR2_X1 U695 ( .A1(n615), .A2(n614), .ZN(n616) );
  NAND2_X1 U696 ( .A1(n617), .A2(n616), .ZN(n618) );
  INV_X1 U697 ( .A(n975), .ZN(n623) );
  INV_X1 U698 ( .A(G1348), .ZN(n619) );
  OR2_X1 U699 ( .A1(n653), .A2(n619), .ZN(n621) );
  NAND2_X1 U700 ( .A1(G2067), .A2(n653), .ZN(n620) );
  NAND2_X1 U701 ( .A1(n621), .A2(n620), .ZN(n622) );
  NAND2_X1 U702 ( .A1(n623), .A2(n639), .ZN(n638) );
  INV_X1 U703 ( .A(G1996), .ZN(n957) );
  NOR2_X1 U704 ( .A1(n661), .A2(n957), .ZN(n624) );
  XOR2_X1 U705 ( .A(n624), .B(KEYINPUT26), .Z(n636) );
  AND2_X1 U706 ( .A1(n675), .A2(G1341), .ZN(n634) );
  NAND2_X1 U707 ( .A1(G56), .A2(n794), .ZN(n625) );
  XOR2_X1 U708 ( .A(KEYINPUT14), .B(n625), .Z(n631) );
  NAND2_X1 U709 ( .A1(n795), .A2(G81), .ZN(n626) );
  XNOR2_X1 U710 ( .A(n626), .B(KEYINPUT12), .ZN(n628) );
  NAND2_X1 U711 ( .A1(G68), .A2(n798), .ZN(n627) );
  NAND2_X1 U712 ( .A1(n628), .A2(n627), .ZN(n629) );
  XOR2_X1 U713 ( .A(KEYINPUT13), .B(n629), .Z(n630) );
  NOR2_X1 U714 ( .A1(n631), .A2(n630), .ZN(n633) );
  NAND2_X1 U715 ( .A1(n799), .A2(G43), .ZN(n632) );
  NAND2_X1 U716 ( .A1(n633), .A2(n632), .ZN(n988) );
  NOR2_X1 U717 ( .A1(n634), .A2(n988), .ZN(n635) );
  AND2_X1 U718 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U719 ( .A1(n638), .A2(n637), .ZN(n642) );
  NAND2_X1 U720 ( .A1(n640), .A2(n975), .ZN(n641) );
  NAND2_X1 U721 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U722 ( .A(n646), .B(n645), .ZN(n651) );
  NAND2_X1 U723 ( .A1(n647), .A2(G299), .ZN(n649) );
  NOR2_X2 U724 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U725 ( .A(n652), .B(KEYINPUT29), .ZN(n660) );
  XNOR2_X1 U726 ( .A(G2078), .B(KEYINPUT25), .ZN(n956) );
  NAND2_X1 U727 ( .A1(n655), .A2(n956), .ZN(n654) );
  XOR2_X1 U728 ( .A(KEYINPUT96), .B(n654), .Z(n657) );
  NOR2_X1 U729 ( .A1(n655), .A2(G1961), .ZN(n656) );
  NOR2_X1 U730 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U731 ( .A(KEYINPUT97), .B(n658), .ZN(n667) );
  NAND2_X1 U732 ( .A1(n667), .A2(G171), .ZN(n659) );
  NAND2_X1 U733 ( .A1(n660), .A2(n659), .ZN(n673) );
  NOR2_X1 U734 ( .A1(G2084), .A2(n675), .ZN(n684) );
  XNOR2_X1 U735 ( .A(n664), .B(KEYINPUT30), .ZN(n666) );
  NOR2_X1 U736 ( .A1(G171), .A2(n667), .ZN(n668) );
  NOR2_X1 U737 ( .A1(n669), .A2(n668), .ZN(n671) );
  XNOR2_X1 U738 ( .A(n671), .B(n670), .ZN(n672) );
  NAND2_X1 U739 ( .A1(n673), .A2(n672), .ZN(n686) );
  NAND2_X1 U740 ( .A1(n686), .A2(G286), .ZN(n674) );
  XNOR2_X1 U741 ( .A(n674), .B(KEYINPUT102), .ZN(n680) );
  NOR2_X1 U742 ( .A1(G1971), .A2(n742), .ZN(n677) );
  NOR2_X1 U743 ( .A1(G2090), .A2(n675), .ZN(n676) );
  NOR2_X1 U744 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U745 ( .A1(n678), .A2(G303), .ZN(n679) );
  NAND2_X1 U746 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U747 ( .A1(n681), .A2(G8), .ZN(n683) );
  XOR2_X1 U748 ( .A(KEYINPUT32), .B(KEYINPUT103), .Z(n682) );
  XNOR2_X1 U749 ( .A(n683), .B(n682), .ZN(n734) );
  NAND2_X1 U750 ( .A1(G8), .A2(n684), .ZN(n688) );
  AND2_X1 U751 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U752 ( .A1(n688), .A2(n687), .ZN(n735) );
  NAND2_X1 U753 ( .A1(G1976), .A2(G288), .ZN(n979) );
  AND2_X1 U754 ( .A1(n735), .A2(n979), .ZN(n689) );
  NAND2_X1 U755 ( .A1(n734), .A2(n689), .ZN(n693) );
  INV_X1 U756 ( .A(n979), .ZN(n691) );
  NOR2_X1 U757 ( .A1(G1976), .A2(G288), .ZN(n978) );
  NOR2_X1 U758 ( .A1(G1971), .A2(G303), .ZN(n985) );
  NOR2_X1 U759 ( .A1(n978), .A2(n985), .ZN(n690) );
  OR2_X1 U760 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U761 ( .A1(n693), .A2(n692), .ZN(n695) );
  NOR2_X1 U762 ( .A1(KEYINPUT33), .A2(n518), .ZN(n733) );
  XOR2_X1 U763 ( .A(G1981), .B(G305), .Z(n972) );
  NOR2_X1 U764 ( .A1(n696), .A2(n697), .ZN(n698) );
  XOR2_X1 U765 ( .A(KEYINPUT91), .B(n698), .Z(n764) );
  NAND2_X1 U766 ( .A1(n594), .A2(G104), .ZN(n699) );
  XNOR2_X1 U767 ( .A(n699), .B(KEYINPUT92), .ZN(n703) );
  NAND2_X1 U768 ( .A1(G140), .A2(n701), .ZN(n702) );
  NAND2_X1 U769 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U770 ( .A(KEYINPUT34), .B(n704), .ZN(n709) );
  NAND2_X1 U771 ( .A1(G128), .A2(n894), .ZN(n706) );
  NAND2_X1 U772 ( .A1(G116), .A2(n891), .ZN(n705) );
  NAND2_X1 U773 ( .A1(n706), .A2(n705), .ZN(n707) );
  XOR2_X1 U774 ( .A(KEYINPUT35), .B(n707), .Z(n708) );
  NOR2_X1 U775 ( .A1(n709), .A2(n708), .ZN(n710) );
  XOR2_X1 U776 ( .A(KEYINPUT36), .B(n710), .Z(n899) );
  XOR2_X1 U777 ( .A(G2067), .B(KEYINPUT37), .Z(n754) );
  NAND2_X1 U778 ( .A1(n899), .A2(n754), .ZN(n711) );
  XNOR2_X1 U779 ( .A(KEYINPUT93), .B(n711), .ZN(n948) );
  NAND2_X1 U780 ( .A1(n764), .A2(n948), .ZN(n761) );
  AND2_X1 U781 ( .A1(n972), .A2(n761), .ZN(n729) );
  NAND2_X1 U782 ( .A1(n701), .A2(G131), .ZN(n712) );
  XNOR2_X1 U783 ( .A(n712), .B(KEYINPUT94), .ZN(n714) );
  NAND2_X1 U784 ( .A1(n894), .A2(G119), .ZN(n713) );
  NAND2_X1 U785 ( .A1(n714), .A2(n713), .ZN(n718) );
  NAND2_X1 U786 ( .A1(G107), .A2(n891), .ZN(n716) );
  NAND2_X1 U787 ( .A1(G95), .A2(n594), .ZN(n715) );
  NAND2_X1 U788 ( .A1(n716), .A2(n715), .ZN(n717) );
  NOR2_X1 U789 ( .A1(n718), .A2(n717), .ZN(n881) );
  INV_X1 U790 ( .A(G1991), .ZN(n952) );
  NOR2_X1 U791 ( .A1(n881), .A2(n952), .ZN(n727) );
  NAND2_X1 U792 ( .A1(G129), .A2(n894), .ZN(n720) );
  NAND2_X1 U793 ( .A1(G117), .A2(n891), .ZN(n719) );
  NAND2_X1 U794 ( .A1(n720), .A2(n719), .ZN(n723) );
  NAND2_X1 U795 ( .A1(n594), .A2(G105), .ZN(n721) );
  XOR2_X1 U796 ( .A(KEYINPUT38), .B(n721), .Z(n722) );
  NOR2_X1 U797 ( .A1(n723), .A2(n722), .ZN(n725) );
  NAND2_X1 U798 ( .A1(G141), .A2(n701), .ZN(n724) );
  NAND2_X1 U799 ( .A1(n725), .A2(n724), .ZN(n869) );
  AND2_X1 U800 ( .A1(n869), .A2(G1996), .ZN(n726) );
  NOR2_X1 U801 ( .A1(n727), .A2(n726), .ZN(n942) );
  INV_X1 U802 ( .A(n764), .ZN(n750) );
  NOR2_X1 U803 ( .A1(n942), .A2(n750), .ZN(n758) );
  INV_X1 U804 ( .A(n758), .ZN(n728) );
  AND2_X1 U805 ( .A1(n729), .A2(n728), .ZN(n731) );
  NAND2_X1 U806 ( .A1(n978), .A2(KEYINPUT33), .ZN(n730) );
  NOR2_X1 U807 ( .A1(n733), .A2(n732), .ZN(n748) );
  NAND2_X1 U808 ( .A1(n735), .A2(n734), .ZN(n738) );
  NOR2_X1 U809 ( .A1(G2090), .A2(G303), .ZN(n736) );
  NAND2_X1 U810 ( .A1(G8), .A2(n736), .ZN(n737) );
  NAND2_X1 U811 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U812 ( .A1(n739), .A2(n742), .ZN(n744) );
  NOR2_X1 U813 ( .A1(G1981), .A2(G305), .ZN(n740) );
  XOR2_X1 U814 ( .A(n740), .B(KEYINPUT24), .Z(n741) );
  OR2_X1 U815 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U816 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U817 ( .A1(n745), .A2(n761), .ZN(n746) );
  NOR2_X1 U818 ( .A1(n746), .A2(n758), .ZN(n747) );
  NOR2_X1 U819 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U820 ( .A(n749), .B(KEYINPUT104), .ZN(n752) );
  XOR2_X1 U821 ( .A(G1986), .B(G290), .Z(n982) );
  NOR2_X1 U822 ( .A1(n750), .A2(n982), .ZN(n751) );
  NOR2_X2 U823 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U824 ( .A(n753), .B(KEYINPUT105), .ZN(n767) );
  OR2_X1 U825 ( .A1(n899), .A2(n754), .ZN(n935) );
  NOR2_X1 U826 ( .A1(G1996), .A2(n869), .ZN(n932) );
  AND2_X1 U827 ( .A1(n952), .A2(n881), .ZN(n940) );
  NOR2_X1 U828 ( .A1(G1986), .A2(G290), .ZN(n755) );
  XNOR2_X1 U829 ( .A(KEYINPUT106), .B(n755), .ZN(n756) );
  NOR2_X1 U830 ( .A1(n940), .A2(n756), .ZN(n757) );
  NOR2_X1 U831 ( .A1(n758), .A2(n757), .ZN(n759) );
  NOR2_X1 U832 ( .A1(n932), .A2(n759), .ZN(n760) );
  XNOR2_X1 U833 ( .A(n760), .B(KEYINPUT39), .ZN(n762) );
  NAND2_X1 U834 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U835 ( .A1(n935), .A2(n763), .ZN(n765) );
  NAND2_X1 U836 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U837 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U838 ( .A(n768), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U839 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U840 ( .A1(G123), .A2(n894), .ZN(n769) );
  XNOR2_X1 U841 ( .A(n769), .B(KEYINPUT18), .ZN(n776) );
  NAND2_X1 U842 ( .A1(G99), .A2(n594), .ZN(n771) );
  NAND2_X1 U843 ( .A1(G135), .A2(n701), .ZN(n770) );
  NAND2_X1 U844 ( .A1(n771), .A2(n770), .ZN(n774) );
  NAND2_X1 U845 ( .A1(G111), .A2(n891), .ZN(n772) );
  XNOR2_X1 U846 ( .A(KEYINPUT77), .B(n772), .ZN(n773) );
  NOR2_X1 U847 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U848 ( .A1(n776), .A2(n775), .ZN(n937) );
  XNOR2_X1 U849 ( .A(G2096), .B(n937), .ZN(n777) );
  OR2_X1 U850 ( .A1(G2100), .A2(n777), .ZN(G156) );
  BUF_X1 U851 ( .A(n778), .Z(G164) );
  INV_X1 U852 ( .A(G120), .ZN(G236) );
  INV_X1 U853 ( .A(G69), .ZN(G235) );
  INV_X1 U854 ( .A(G57), .ZN(G237) );
  NAND2_X1 U855 ( .A1(G7), .A2(G661), .ZN(n779) );
  XNOR2_X1 U856 ( .A(n779), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U857 ( .A(G223), .ZN(n834) );
  NAND2_X1 U858 ( .A1(n834), .A2(G567), .ZN(n780) );
  XOR2_X1 U859 ( .A(KEYINPUT11), .B(n780), .Z(G234) );
  INV_X1 U860 ( .A(G860), .ZN(n785) );
  OR2_X1 U861 ( .A1(n988), .A2(n785), .ZN(G153) );
  INV_X1 U862 ( .A(G171), .ZN(G301) );
  NAND2_X1 U863 ( .A1(G868), .A2(G301), .ZN(n782) );
  OR2_X1 U864 ( .A1(n975), .A2(G868), .ZN(n781) );
  NAND2_X1 U865 ( .A1(n782), .A2(n781), .ZN(G284) );
  NAND2_X1 U866 ( .A1(G286), .A2(G868), .ZN(n784) );
  INV_X1 U867 ( .A(G868), .ZN(n814) );
  NAND2_X1 U868 ( .A1(G299), .A2(n814), .ZN(n783) );
  NAND2_X1 U869 ( .A1(n784), .A2(n783), .ZN(G297) );
  NAND2_X1 U870 ( .A1(n785), .A2(G559), .ZN(n786) );
  NAND2_X1 U871 ( .A1(n786), .A2(n975), .ZN(n787) );
  XNOR2_X1 U872 ( .A(n787), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U873 ( .A1(G868), .A2(n988), .ZN(n788) );
  XNOR2_X1 U874 ( .A(KEYINPUT76), .B(n788), .ZN(n791) );
  NAND2_X1 U875 ( .A1(G868), .A2(n975), .ZN(n789) );
  NOR2_X1 U876 ( .A1(G559), .A2(n789), .ZN(n790) );
  NOR2_X1 U877 ( .A1(n791), .A2(n790), .ZN(G282) );
  XNOR2_X1 U878 ( .A(n988), .B(KEYINPUT78), .ZN(n793) );
  NAND2_X1 U879 ( .A1(n975), .A2(G559), .ZN(n792) );
  XNOR2_X1 U880 ( .A(n793), .B(n792), .ZN(n811) );
  NOR2_X1 U881 ( .A1(G860), .A2(n811), .ZN(n804) );
  NAND2_X1 U882 ( .A1(G67), .A2(n794), .ZN(n797) );
  NAND2_X1 U883 ( .A1(G93), .A2(n795), .ZN(n796) );
  NAND2_X1 U884 ( .A1(n797), .A2(n796), .ZN(n803) );
  NAND2_X1 U885 ( .A1(G80), .A2(n798), .ZN(n801) );
  NAND2_X1 U886 ( .A1(G55), .A2(n799), .ZN(n800) );
  NAND2_X1 U887 ( .A1(n801), .A2(n800), .ZN(n802) );
  OR2_X1 U888 ( .A1(n803), .A2(n802), .ZN(n813) );
  XOR2_X1 U889 ( .A(n804), .B(n813), .Z(G145) );
  XOR2_X1 U890 ( .A(KEYINPUT83), .B(KEYINPUT19), .Z(n805) );
  XNOR2_X1 U891 ( .A(G288), .B(n805), .ZN(n808) );
  XNOR2_X1 U892 ( .A(G305), .B(G299), .ZN(n806) );
  XNOR2_X1 U893 ( .A(n806), .B(G303), .ZN(n807) );
  XNOR2_X1 U894 ( .A(n808), .B(n807), .ZN(n810) );
  XOR2_X1 U895 ( .A(G290), .B(n813), .Z(n809) );
  XNOR2_X1 U896 ( .A(n810), .B(n809), .ZN(n903) );
  XNOR2_X1 U897 ( .A(n811), .B(n903), .ZN(n812) );
  NAND2_X1 U898 ( .A1(n812), .A2(G868), .ZN(n816) );
  NAND2_X1 U899 ( .A1(n814), .A2(n813), .ZN(n815) );
  NAND2_X1 U900 ( .A1(n816), .A2(n815), .ZN(G295) );
  NAND2_X1 U901 ( .A1(G2078), .A2(G2084), .ZN(n817) );
  XOR2_X1 U902 ( .A(KEYINPUT20), .B(n817), .Z(n818) );
  NAND2_X1 U903 ( .A1(G2090), .A2(n818), .ZN(n819) );
  XNOR2_X1 U904 ( .A(KEYINPUT21), .B(n819), .ZN(n820) );
  NAND2_X1 U905 ( .A1(n820), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U906 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U907 ( .A(KEYINPUT72), .B(G132), .Z(G219) );
  XNOR2_X1 U908 ( .A(KEYINPUT73), .B(G82), .ZN(G220) );
  NOR2_X1 U909 ( .A1(G235), .A2(G236), .ZN(n821) );
  XNOR2_X1 U910 ( .A(n821), .B(KEYINPUT85), .ZN(n822) );
  NOR2_X1 U911 ( .A1(G237), .A2(n822), .ZN(n823) );
  XNOR2_X1 U912 ( .A(KEYINPUT86), .B(n823), .ZN(n824) );
  NAND2_X1 U913 ( .A1(n824), .A2(G108), .ZN(n839) );
  AND2_X1 U914 ( .A1(G567), .A2(n839), .ZN(n830) );
  NOR2_X1 U915 ( .A1(G219), .A2(G220), .ZN(n825) );
  XOR2_X1 U916 ( .A(KEYINPUT22), .B(n825), .Z(n826) );
  NOR2_X1 U917 ( .A1(G218), .A2(n826), .ZN(n827) );
  NAND2_X1 U918 ( .A1(G96), .A2(n827), .ZN(n838) );
  NAND2_X1 U919 ( .A1(G2106), .A2(n838), .ZN(n828) );
  XOR2_X1 U920 ( .A(KEYINPUT84), .B(n828), .Z(n829) );
  NOR2_X1 U921 ( .A1(n830), .A2(n829), .ZN(G319) );
  NAND2_X1 U922 ( .A1(G661), .A2(G483), .ZN(n831) );
  XNOR2_X1 U923 ( .A(KEYINPUT87), .B(n831), .ZN(n832) );
  NAND2_X1 U924 ( .A1(n832), .A2(G319), .ZN(n833) );
  XOR2_X1 U925 ( .A(KEYINPUT88), .B(n833), .Z(n837) );
  NAND2_X1 U926 ( .A1(G36), .A2(n837), .ZN(G176) );
  NAND2_X1 U927 ( .A1(G2106), .A2(n834), .ZN(G217) );
  AND2_X1 U928 ( .A1(G15), .A2(G2), .ZN(n835) );
  NAND2_X1 U929 ( .A1(G661), .A2(n835), .ZN(G259) );
  NAND2_X1 U930 ( .A1(G3), .A2(G1), .ZN(n836) );
  NAND2_X1 U931 ( .A1(n837), .A2(n836), .ZN(G188) );
  INV_X1 U933 ( .A(G108), .ZN(G238) );
  INV_X1 U934 ( .A(G96), .ZN(G221) );
  NOR2_X1 U935 ( .A1(n839), .A2(n838), .ZN(G325) );
  INV_X1 U936 ( .A(G325), .ZN(G261) );
  XOR2_X1 U937 ( .A(G1981), .B(G1966), .Z(n841) );
  XNOR2_X1 U938 ( .A(G1996), .B(G1991), .ZN(n840) );
  XNOR2_X1 U939 ( .A(n841), .B(n840), .ZN(n851) );
  XOR2_X1 U940 ( .A(KEYINPUT112), .B(KEYINPUT41), .Z(n843) );
  XNOR2_X1 U941 ( .A(G1986), .B(KEYINPUT113), .ZN(n842) );
  XNOR2_X1 U942 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U943 ( .A(G1976), .B(G1971), .Z(n845) );
  XNOR2_X1 U944 ( .A(G1961), .B(G1956), .ZN(n844) );
  XNOR2_X1 U945 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U946 ( .A(n847), .B(n846), .Z(n849) );
  XNOR2_X1 U947 ( .A(KEYINPUT111), .B(G2474), .ZN(n848) );
  XNOR2_X1 U948 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U949 ( .A(n851), .B(n850), .Z(G229) );
  XOR2_X1 U950 ( .A(G2096), .B(KEYINPUT43), .Z(n853) );
  XNOR2_X1 U951 ( .A(G2090), .B(G2678), .ZN(n852) );
  XNOR2_X1 U952 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U953 ( .A(n854), .B(KEYINPUT110), .Z(n856) );
  XNOR2_X1 U954 ( .A(G2067), .B(G2072), .ZN(n855) );
  XNOR2_X1 U955 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U956 ( .A(KEYINPUT42), .B(G2100), .Z(n858) );
  XNOR2_X1 U957 ( .A(G2078), .B(G2084), .ZN(n857) );
  XNOR2_X1 U958 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U959 ( .A(n860), .B(n859), .ZN(G227) );
  NAND2_X1 U960 ( .A1(G112), .A2(n891), .ZN(n862) );
  NAND2_X1 U961 ( .A1(G100), .A2(n594), .ZN(n861) );
  NAND2_X1 U962 ( .A1(n862), .A2(n861), .ZN(n863) );
  XNOR2_X1 U963 ( .A(KEYINPUT114), .B(n863), .ZN(n868) );
  NAND2_X1 U964 ( .A1(n894), .A2(G124), .ZN(n864) );
  XNOR2_X1 U965 ( .A(n864), .B(KEYINPUT44), .ZN(n866) );
  NAND2_X1 U966 ( .A1(G136), .A2(n701), .ZN(n865) );
  NAND2_X1 U967 ( .A1(n866), .A2(n865), .ZN(n867) );
  NOR2_X1 U968 ( .A1(n868), .A2(n867), .ZN(G162) );
  XOR2_X1 U969 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n871) );
  XOR2_X1 U970 ( .A(n869), .B(KEYINPUT118), .Z(n870) );
  XNOR2_X1 U971 ( .A(n871), .B(n870), .ZN(n880) );
  NAND2_X1 U972 ( .A1(G127), .A2(n894), .ZN(n873) );
  NAND2_X1 U973 ( .A1(G115), .A2(n891), .ZN(n872) );
  NAND2_X1 U974 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U975 ( .A(n874), .B(KEYINPUT47), .ZN(n876) );
  NAND2_X1 U976 ( .A1(G103), .A2(n594), .ZN(n875) );
  NAND2_X1 U977 ( .A1(n876), .A2(n875), .ZN(n879) );
  NAND2_X1 U978 ( .A1(G139), .A2(n701), .ZN(n877) );
  XNOR2_X1 U979 ( .A(KEYINPUT117), .B(n877), .ZN(n878) );
  NOR2_X1 U980 ( .A1(n879), .A2(n878), .ZN(n927) );
  XOR2_X1 U981 ( .A(n880), .B(n927), .Z(n883) );
  XNOR2_X1 U982 ( .A(G160), .B(n881), .ZN(n882) );
  XNOR2_X1 U983 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U984 ( .A(n937), .B(n884), .ZN(n886) );
  XNOR2_X1 U985 ( .A(G164), .B(G162), .ZN(n885) );
  XNOR2_X1 U986 ( .A(n886), .B(n885), .ZN(n901) );
  NAND2_X1 U987 ( .A1(G142), .A2(n701), .ZN(n887) );
  XNOR2_X1 U988 ( .A(n887), .B(KEYINPUT116), .ZN(n889) );
  NAND2_X1 U989 ( .A1(G106), .A2(n594), .ZN(n888) );
  NAND2_X1 U990 ( .A1(n889), .A2(n888), .ZN(n890) );
  XNOR2_X1 U991 ( .A(n890), .B(KEYINPUT45), .ZN(n893) );
  NAND2_X1 U992 ( .A1(G118), .A2(n891), .ZN(n892) );
  NAND2_X1 U993 ( .A1(n893), .A2(n892), .ZN(n897) );
  NAND2_X1 U994 ( .A1(G130), .A2(n894), .ZN(n895) );
  XNOR2_X1 U995 ( .A(KEYINPUT115), .B(n895), .ZN(n896) );
  NOR2_X1 U996 ( .A1(n897), .A2(n896), .ZN(n898) );
  XNOR2_X1 U997 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U998 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U999 ( .A1(G37), .A2(n902), .ZN(G395) );
  XOR2_X1 U1000 ( .A(KEYINPUT119), .B(n903), .Z(n905) );
  XNOR2_X1 U1001 ( .A(G171), .B(G286), .ZN(n904) );
  XNOR2_X1 U1002 ( .A(n905), .B(n904), .ZN(n907) );
  XOR2_X1 U1003 ( .A(n988), .B(n975), .Z(n906) );
  XNOR2_X1 U1004 ( .A(n907), .B(n906), .ZN(n908) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n908), .ZN(G397) );
  XOR2_X1 U1006 ( .A(G2443), .B(G2451), .Z(n910) );
  XNOR2_X1 U1007 ( .A(G2454), .B(G2427), .ZN(n909) );
  XNOR2_X1 U1008 ( .A(n910), .B(n909), .ZN(n911) );
  XOR2_X1 U1009 ( .A(n911), .B(G2430), .Z(n913) );
  XNOR2_X1 U1010 ( .A(G1341), .B(G1348), .ZN(n912) );
  XNOR2_X1 U1011 ( .A(n913), .B(n912), .ZN(n917) );
  XOR2_X1 U1012 ( .A(KEYINPUT108), .B(G2435), .Z(n915) );
  XNOR2_X1 U1013 ( .A(KEYINPUT109), .B(G2438), .ZN(n914) );
  XNOR2_X1 U1014 ( .A(n915), .B(n914), .ZN(n916) );
  XOR2_X1 U1015 ( .A(n917), .B(n916), .Z(n919) );
  XNOR2_X1 U1016 ( .A(G2446), .B(KEYINPUT107), .ZN(n918) );
  XNOR2_X1 U1017 ( .A(n919), .B(n918), .ZN(n920) );
  NAND2_X1 U1018 ( .A1(n920), .A2(G14), .ZN(n926) );
  NAND2_X1 U1019 ( .A1(G319), .A2(n926), .ZN(n923) );
  NOR2_X1 U1020 ( .A1(G229), .A2(G227), .ZN(n921) );
  XNOR2_X1 U1021 ( .A(KEYINPUT49), .B(n921), .ZN(n922) );
  NOR2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(n925) );
  NOR2_X1 U1023 ( .A1(G395), .A2(G397), .ZN(n924) );
  NAND2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(G225) );
  INV_X1 U1025 ( .A(G225), .ZN(G308) );
  INV_X1 U1026 ( .A(G303), .ZN(G166) );
  INV_X1 U1027 ( .A(n926), .ZN(G401) );
  XOR2_X1 U1028 ( .A(G2072), .B(n927), .Z(n929) );
  XOR2_X1 U1029 ( .A(G164), .B(G2078), .Z(n928) );
  NOR2_X1 U1030 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1031 ( .A(KEYINPUT50), .B(n930), .ZN(n946) );
  XOR2_X1 U1032 ( .A(G2090), .B(G162), .Z(n931) );
  NOR2_X1 U1033 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1034 ( .A(KEYINPUT120), .B(n933), .Z(n934) );
  XNOR2_X1 U1035 ( .A(n934), .B(KEYINPUT51), .ZN(n936) );
  NAND2_X1 U1036 ( .A1(n936), .A2(n935), .ZN(n944) );
  XNOR2_X1 U1037 ( .A(G160), .B(G2084), .ZN(n938) );
  NAND2_X1 U1038 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1040 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1041 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1042 ( .A1(n946), .A2(n945), .ZN(n947) );
  NOR2_X1 U1043 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1044 ( .A(KEYINPUT52), .B(n949), .ZN(n950) );
  INV_X1 U1045 ( .A(KEYINPUT55), .ZN(n1029) );
  NAND2_X1 U1046 ( .A1(n950), .A2(n1029), .ZN(n951) );
  NAND2_X1 U1047 ( .A1(n951), .A2(G29), .ZN(n1036) );
  XNOR2_X1 U1048 ( .A(G2090), .B(G35), .ZN(n966) );
  XNOR2_X1 U1049 ( .A(G25), .B(n952), .ZN(n953) );
  NAND2_X1 U1050 ( .A1(n953), .A2(G28), .ZN(n963) );
  XNOR2_X1 U1051 ( .A(G2067), .B(G26), .ZN(n955) );
  XNOR2_X1 U1052 ( .A(G33), .B(G2072), .ZN(n954) );
  NOR2_X1 U1053 ( .A1(n955), .A2(n954), .ZN(n961) );
  XOR2_X1 U1054 ( .A(n956), .B(G27), .Z(n959) );
  XOR2_X1 U1055 ( .A(n957), .B(G32), .Z(n958) );
  NOR2_X1 U1056 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1057 ( .A1(n961), .A2(n960), .ZN(n962) );
  NOR2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1059 ( .A(KEYINPUT53), .B(n964), .ZN(n965) );
  NOR2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n969) );
  XOR2_X1 U1061 ( .A(G2084), .B(G34), .Z(n967) );
  XNOR2_X1 U1062 ( .A(KEYINPUT54), .B(n967), .ZN(n968) );
  NAND2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n1030) );
  NOR2_X1 U1064 ( .A1(G29), .A2(KEYINPUT55), .ZN(n970) );
  NAND2_X1 U1065 ( .A1(n1030), .A2(n970), .ZN(n971) );
  NAND2_X1 U1066 ( .A1(G11), .A2(n971), .ZN(n1034) );
  XNOR2_X1 U1067 ( .A(G16), .B(KEYINPUT56), .ZN(n998) );
  XNOR2_X1 U1068 ( .A(G1966), .B(G168), .ZN(n973) );
  NAND2_X1 U1069 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1070 ( .A(n974), .B(KEYINPUT57), .ZN(n996) );
  XOR2_X1 U1071 ( .A(G299), .B(G1956), .Z(n977) );
  XNOR2_X1 U1072 ( .A(n975), .B(G1348), .ZN(n976) );
  NAND2_X1 U1073 ( .A1(n977), .A2(n976), .ZN(n994) );
  INV_X1 U1074 ( .A(n978), .ZN(n980) );
  NAND2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1076 ( .A(n981), .B(KEYINPUT121), .ZN(n983) );
  NAND2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n984) );
  NOR2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n992) );
  XNOR2_X1 U1079 ( .A(G171), .B(G1961), .ZN(n987) );
  NAND2_X1 U1080 ( .A1(G1971), .A2(G303), .ZN(n986) );
  NAND2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n990) );
  XNOR2_X1 U1082 ( .A(G1341), .B(n988), .ZN(n989) );
  NOR2_X1 U1083 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n993) );
  NOR2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n1027) );
  INV_X1 U1088 ( .A(G16), .ZN(n1025) );
  XNOR2_X1 U1089 ( .A(G1986), .B(G24), .ZN(n1003) );
  XNOR2_X1 U1090 ( .A(G1971), .B(G22), .ZN(n1000) );
  XNOR2_X1 U1091 ( .A(G1976), .B(G23), .ZN(n999) );
  NOR2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1093 ( .A(KEYINPUT125), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1095 ( .A(KEYINPUT126), .B(n1004), .ZN(n1005) );
  XNOR2_X1 U1096 ( .A(n1005), .B(KEYINPUT58), .ZN(n1020) );
  XNOR2_X1 U1097 ( .A(G1966), .B(G21), .ZN(n1018) );
  XOR2_X1 U1098 ( .A(G1341), .B(G19), .Z(n1007) );
  XOR2_X1 U1099 ( .A(G1981), .B(G6), .Z(n1006) );
  NAND2_X1 U1100 ( .A1(n1007), .A2(n1006), .ZN(n1009) );
  XNOR2_X1 U1101 ( .A(G20), .B(G1956), .ZN(n1008) );
  NOR2_X1 U1102 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1103 ( .A(KEYINPUT122), .B(n1010), .ZN(n1014) );
  XOR2_X1 U1104 ( .A(KEYINPUT123), .B(G4), .Z(n1012) );
  XNOR2_X1 U1105 ( .A(G1348), .B(KEYINPUT59), .ZN(n1011) );
  XNOR2_X1 U1106 ( .A(n1012), .B(n1011), .ZN(n1013) );
  NAND2_X1 U1107 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1108 ( .A(n1015), .B(KEYINPUT124), .ZN(n1016) );
  XNOR2_X1 U1109 ( .A(n1016), .B(KEYINPUT60), .ZN(n1017) );
  NOR2_X1 U1110 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1111 ( .A1(n1020), .A2(n1019), .ZN(n1022) );
  XNOR2_X1 U1112 ( .A(G5), .B(G1961), .ZN(n1021) );
  NOR2_X1 U1113 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1114 ( .A(KEYINPUT61), .B(n1023), .ZN(n1024) );
  NAND2_X1 U1115 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1116 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1117 ( .A(n1028), .B(KEYINPUT127), .ZN(n1032) );
  OR2_X1 U1118 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1119 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NOR2_X1 U1120 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NAND2_X1 U1121 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  XOR2_X1 U1122 ( .A(KEYINPUT62), .B(n1037), .Z(G311) );
  INV_X1 U1123 ( .A(G311), .ZN(G150) );
endmodule

