//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 0 0 0 1 1 1 1 1 1 0 0 1 1 0 0 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 1 1 0 1 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 0 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:50 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT77), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n190), .B(KEYINPUT22), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n191), .B(G137), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G140), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G125), .ZN(new_n195));
  INV_X1    g009(.A(G125), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G140), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n195), .A2(new_n197), .A3(KEYINPUT16), .ZN(new_n198));
  OR3_X1    g012(.A1(new_n196), .A2(KEYINPUT16), .A3(G140), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n198), .A2(new_n199), .A3(G146), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  AOI21_X1  g015(.A(G146), .B1(new_n198), .B2(new_n199), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G128), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(G119), .ZN(new_n205));
  XNOR2_X1  g019(.A(KEYINPUT67), .B(G128), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n205), .B1(new_n207), .B2(G119), .ZN(new_n208));
  XOR2_X1   g022(.A(KEYINPUT24), .B(G110), .Z(new_n209));
  AOI21_X1  g023(.A(new_n203), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n207), .A2(KEYINPUT23), .A3(G119), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT73), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n212), .B(KEYINPUT23), .C1(new_n204), .C2(G119), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT23), .ZN(new_n215));
  INV_X1    g029(.A(G119), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n215), .B1(new_n216), .B2(G128), .ZN(new_n217));
  OAI22_X1  g031(.A1(new_n217), .A2(new_n212), .B1(new_n216), .B2(G128), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n211), .B1(new_n214), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G110), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n210), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT74), .B(G110), .ZN(new_n222));
  OAI22_X1  g036(.A1(new_n219), .A2(new_n222), .B1(new_n208), .B2(new_n209), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n195), .A2(new_n197), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT75), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT75), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n195), .A2(new_n197), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G146), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n225), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  XNOR2_X1  g043(.A(new_n229), .B(KEYINPUT76), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n223), .A2(new_n230), .A3(new_n200), .ZN(new_n231));
  AOI211_X1 g045(.A(new_n188), .B(new_n193), .C1(new_n221), .C2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n192), .A2(KEYINPUT77), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n193), .A2(new_n188), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n221), .A2(new_n231), .A3(new_n233), .A4(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n187), .B1(new_n232), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(KEYINPUT25), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n221), .A2(new_n231), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n239), .A2(KEYINPUT77), .A3(new_n192), .ZN(new_n240));
  AOI21_X1  g054(.A(G902), .B1(new_n240), .B2(new_n235), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT25), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G217), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n244), .B1(G234), .B2(new_n187), .ZN(new_n245));
  AND3_X1   g059(.A1(new_n238), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n245), .A2(G902), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n247), .B1(new_n232), .B2(new_n236), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT78), .ZN(new_n249));
  XNOR2_X1  g063(.A(new_n248), .B(new_n249), .ZN(new_n250));
  OR2_X1    g064(.A1(new_n246), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G472), .ZN(new_n252));
  INV_X1    g066(.A(G134), .ZN(new_n253));
  OAI21_X1  g067(.A(KEYINPUT66), .B1(new_n253), .B2(G137), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT66), .ZN(new_n255));
  INV_X1    g069(.A(G137), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n255), .A2(new_n256), .A3(G134), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n253), .A2(G137), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n254), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G131), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT11), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n261), .B1(new_n253), .B2(G137), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n256), .A2(KEYINPUT11), .A3(G134), .ZN(new_n263));
  INV_X1    g077(.A(G131), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n262), .A2(new_n263), .A3(new_n264), .A4(new_n258), .ZN(new_n265));
  INV_X1    g079(.A(G143), .ZN(new_n266));
  OAI21_X1  g080(.A(KEYINPUT1), .B1(new_n266), .B2(G146), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n228), .A2(G143), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(G146), .ZN(new_n269));
  AOI22_X1  g083(.A1(new_n206), .A2(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT1), .ZN(new_n271));
  AND4_X1   g085(.A1(new_n271), .A2(new_n268), .A3(new_n269), .A4(G128), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n260), .B(new_n265), .C1(new_n270), .C2(new_n272), .ZN(new_n273));
  XNOR2_X1  g087(.A(G116), .B(G119), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  XNOR2_X1  g089(.A(KEYINPUT2), .B(G113), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n276), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(new_n274), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n262), .A2(new_n258), .A3(new_n263), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G131), .ZN(new_n282));
  AND2_X1   g096(.A1(new_n282), .A2(new_n265), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT65), .ZN(new_n284));
  XNOR2_X1  g098(.A(G143), .B(G146), .ZN(new_n285));
  XNOR2_X1  g099(.A(KEYINPUT0), .B(G128), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n268), .A2(new_n269), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n204), .A2(KEYINPUT0), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT0), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G128), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n288), .A2(new_n292), .A3(KEYINPUT65), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n285), .A2(KEYINPUT0), .A3(G128), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n287), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n273), .B(new_n280), .C1(new_n283), .C2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT68), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT27), .ZN(new_n298));
  INV_X1    g112(.A(G237), .ZN(new_n299));
  AND4_X1   g113(.A1(new_n298), .A2(new_n299), .A3(new_n189), .A4(G210), .ZN(new_n300));
  NOR2_X1   g114(.A1(G237), .A2(G953), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n298), .B1(new_n301), .B2(G210), .ZN(new_n302));
  OAI21_X1  g116(.A(KEYINPUT26), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n299), .A2(new_n189), .A3(G210), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT27), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT26), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n301), .A2(new_n298), .A3(G210), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  AND3_X1   g122(.A1(new_n303), .A2(G101), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(G101), .B1(new_n303), .B2(new_n308), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AND3_X1   g125(.A1(new_n296), .A2(new_n297), .A3(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n297), .B1(new_n296), .B2(new_n311), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n277), .A2(new_n279), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT64), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT30), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n288), .A2(new_n292), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n268), .A2(new_n269), .A3(G128), .ZN(new_n319));
  AOI22_X1  g133(.A1(new_n318), .A2(new_n284), .B1(new_n319), .B2(KEYINPUT0), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n282), .A2(new_n265), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n321), .A3(new_n293), .ZN(new_n322));
  AOI211_X1 g136(.A(new_n316), .B(new_n317), .C1(new_n322), .C2(new_n273), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n273), .B1(new_n283), .B2(new_n295), .ZN(new_n324));
  AOI21_X1  g138(.A(KEYINPUT30), .B1(new_n324), .B2(KEYINPUT64), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n315), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT31), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n314), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n311), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n315), .B1(new_n324), .B2(KEYINPUT69), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT69), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n322), .A2(new_n331), .A3(new_n273), .ZN(new_n332));
  AOI21_X1  g146(.A(KEYINPUT28), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT28), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n324), .A2(new_n315), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n334), .B1(new_n335), .B2(new_n296), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n329), .B1(new_n333), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n328), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n327), .B1(new_n314), .B2(new_n326), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n252), .B(new_n187), .C1(new_n338), .C2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT70), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT32), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n324), .A2(KEYINPUT64), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n317), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n324), .A2(KEYINPUT64), .A3(KEYINPUT30), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n280), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n296), .A2(new_n311), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT68), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n296), .A2(new_n311), .A3(new_n297), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(KEYINPUT31), .B1(new_n346), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n351), .A2(new_n337), .A3(new_n328), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT70), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n352), .A2(new_n353), .A3(new_n252), .A4(new_n187), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n341), .A2(new_n342), .A3(new_n354), .ZN(new_n355));
  OR2_X1    g169(.A1(new_n340), .A2(new_n342), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT72), .ZN(new_n358));
  NOR3_X1   g172(.A1(new_n333), .A2(new_n336), .A3(new_n329), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(KEYINPUT29), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n187), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT71), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n326), .A2(new_n296), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n362), .B1(new_n363), .B2(new_n329), .ZN(new_n364));
  AOI211_X1 g178(.A(KEYINPUT71), .B(new_n311), .C1(new_n326), .C2(new_n296), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n359), .A2(KEYINPUT29), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n361), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n358), .B1(new_n368), .B2(new_n252), .ZN(new_n369));
  INV_X1    g183(.A(new_n296), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n346), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(KEYINPUT71), .B1(new_n371), .B2(new_n311), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n363), .A2(new_n362), .A3(new_n329), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n372), .A2(new_n367), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(G902), .B1(new_n359), .B2(KEYINPUT29), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(KEYINPUT72), .A3(G472), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n369), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n251), .B1(new_n357), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g193(.A(G210), .B1(G237), .B2(G902), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT5), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n381), .A2(new_n216), .A3(G116), .ZN(new_n382));
  OAI211_X1 g196(.A(G113), .B(new_n382), .C1(new_n275), .C2(new_n381), .ZN(new_n383));
  AND2_X1   g197(.A1(new_n383), .A2(new_n279), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT79), .ZN(new_n385));
  INV_X1    g199(.A(G104), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n385), .B1(new_n386), .B2(G107), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(G107), .ZN(new_n388));
  INV_X1    g202(.A(G107), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(KEYINPUT79), .A3(G104), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n387), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(G101), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT80), .ZN(new_n393));
  OAI21_X1  g207(.A(KEYINPUT3), .B1(new_n386), .B2(G107), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT3), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n395), .A2(new_n389), .A3(G104), .ZN(new_n396));
  INV_X1    g210(.A(G101), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n394), .A2(new_n396), .A3(new_n397), .A4(new_n388), .ZN(new_n398));
  AND3_X1   g212(.A1(new_n392), .A2(new_n393), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n393), .B1(new_n392), .B2(new_n398), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n384), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n394), .A2(new_n396), .A3(new_n388), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G101), .ZN(new_n403));
  OR2_X1    g217(.A1(new_n403), .A2(KEYINPUT4), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n403), .A2(KEYINPUT4), .A3(new_n398), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n404), .A2(new_n315), .A3(new_n405), .ZN(new_n406));
  XNOR2_X1  g220(.A(G110), .B(G122), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n401), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n295), .A2(G125), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n270), .A2(new_n272), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n196), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n189), .A2(G224), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n409), .A2(new_n411), .A3(KEYINPUT7), .A4(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n409), .A2(new_n411), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT7), .ZN(new_n415));
  INV_X1    g229(.A(new_n412), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n414), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  AND3_X1   g231(.A1(new_n408), .A2(new_n413), .A3(new_n417), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n392), .A2(new_n398), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n401), .B1(new_n419), .B2(new_n384), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n407), .B(KEYINPUT8), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(G902), .B1(new_n418), .B2(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n414), .B(new_n416), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n401), .A2(new_n406), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT82), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n407), .A2(new_n426), .ZN(new_n427));
  AOI22_X1  g241(.A1(new_n408), .A2(KEYINPUT6), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  AND3_X1   g242(.A1(new_n425), .A2(KEYINPUT6), .A3(new_n427), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n424), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n380), .B1(new_n423), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n423), .A2(new_n430), .A3(new_n380), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(KEYINPUT83), .A3(new_n433), .ZN(new_n434));
  OR2_X1    g248(.A1(new_n433), .A2(KEYINPUT83), .ZN(new_n435));
  AND2_X1   g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(KEYINPUT9), .B(G234), .ZN(new_n437));
  OAI21_X1  g251(.A(G221), .B1(new_n437), .B2(G902), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(G214), .B1(G237), .B2(G902), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(G469), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n444), .A2(new_n187), .ZN(new_n445));
  OAI221_X1 g259(.A(KEYINPUT10), .B1(new_n270), .B2(new_n272), .C1(new_n399), .C2(new_n400), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n204), .B1(new_n268), .B2(KEYINPUT1), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n447), .A2(new_n285), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n419), .B1(new_n272), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT10), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n404), .A2(new_n293), .A3(new_n320), .A4(new_n405), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n446), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n321), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n446), .A2(new_n451), .A3(new_n283), .A4(new_n452), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g270(.A(G110), .B(G140), .ZN(new_n457));
  AND2_X1   g271(.A1(new_n189), .A2(G227), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n457), .B(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n459), .ZN(new_n461));
  INV_X1    g275(.A(new_n399), .ZN(new_n462));
  INV_X1    g276(.A(new_n400), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n462), .A2(new_n410), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n449), .ZN(new_n465));
  AOI21_X1  g279(.A(KEYINPUT12), .B1(new_n465), .B2(new_n321), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT12), .ZN(new_n467));
  AOI211_X1 g281(.A(new_n467), .B(new_n283), .C1(new_n464), .C2(new_n449), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n461), .B(new_n455), .C1(new_n466), .C2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(G902), .B1(new_n460), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n445), .B1(new_n470), .B2(new_n444), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n455), .B1(new_n466), .B2(new_n468), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n459), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n455), .A2(new_n461), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT81), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n455), .A2(KEYINPUT81), .A3(new_n461), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n476), .A2(new_n454), .A3(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n473), .A2(new_n478), .A3(G469), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n443), .B1(new_n471), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n436), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(G475), .ZN(new_n483));
  XNOR2_X1  g297(.A(G113), .B(G122), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n484), .B(new_n386), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n224), .A2(G146), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(KEYINPUT86), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n229), .A2(KEYINPUT76), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n229), .A2(KEYINPUT76), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT84), .ZN(new_n491));
  INV_X1    g305(.A(G214), .ZN(new_n492));
  NOR3_X1   g306(.A1(new_n492), .A2(G237), .A3(G953), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n491), .B1(new_n493), .B2(G143), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n299), .A2(new_n189), .A3(G214), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n495), .A2(KEYINPUT84), .A3(new_n266), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n299), .A2(new_n189), .A3(G143), .A4(G214), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT85), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n301), .A2(KEYINPUT85), .A3(G143), .A4(G214), .ZN(new_n500));
  AOI22_X1  g314(.A1(new_n494), .A2(new_n496), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  AND2_X1   g315(.A1(KEYINPUT18), .A2(G131), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n501), .B(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n490), .A2(new_n503), .ZN(new_n504));
  AOI211_X1 g318(.A(G143), .B(new_n491), .C1(new_n301), .C2(G214), .ZN(new_n505));
  AOI21_X1  g319(.A(KEYINPUT84), .B1(new_n495), .B2(new_n266), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AND2_X1   g321(.A1(new_n499), .A2(new_n500), .ZN(new_n508));
  OAI211_X1 g322(.A(KEYINPUT17), .B(G131), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(KEYINPUT87), .A3(new_n203), .ZN(new_n510));
  OAI21_X1  g324(.A(G131), .B1(new_n507), .B2(new_n508), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n501), .A2(new_n264), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT17), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(KEYINPUT87), .B1(new_n509), .B2(new_n203), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n485), .B(new_n504), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(KEYINPUT88), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n509), .A2(new_n203), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT87), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n521), .A2(new_n514), .A3(new_n510), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT88), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n522), .A2(new_n523), .A3(new_n485), .A4(new_n504), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n518), .A2(new_n524), .ZN(new_n525));
  AND2_X1   g339(.A1(new_n522), .A2(new_n504), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n525), .B1(new_n485), .B2(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n483), .B1(new_n527), .B2(new_n187), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n511), .A2(new_n512), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n224), .A2(KEYINPUT19), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n225), .A2(new_n227), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n530), .B1(new_n531), .B2(KEYINPUT19), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n529), .B(new_n200), .C1(G146), .C2(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n485), .B1(new_n533), .B2(new_n504), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n525), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT89), .ZN(new_n537));
  NOR2_X1   g351(.A1(G475), .A2(G902), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT89), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n525), .A2(new_n539), .A3(new_n535), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n537), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(KEYINPUT20), .ZN(new_n542));
  INV_X1    g356(.A(new_n538), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n543), .A2(KEYINPUT20), .ZN(new_n544));
  MUX2_X1   g358(.A(new_n543), .B(new_n544), .S(KEYINPUT90), .Z(new_n545));
  NAND2_X1  g359(.A1(new_n536), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n528), .B1(new_n542), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(G478), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n548), .A2(KEYINPUT15), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT92), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT91), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n207), .A2(G143), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n204), .A2(G143), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n551), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n206), .A2(new_n266), .ZN(new_n556));
  NOR3_X1   g370(.A1(new_n556), .A2(KEYINPUT91), .A3(new_n553), .ZN(new_n557));
  OR3_X1    g371(.A1(new_n555), .A2(new_n557), .A3(new_n253), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n253), .B1(new_n555), .B2(new_n557), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(G116), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n561), .A2(KEYINPUT14), .A3(G122), .ZN(new_n562));
  XNOR2_X1  g376(.A(G116), .B(G122), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n562), .B(G107), .C1(new_n564), .C2(KEYINPUT14), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n563), .A2(new_n389), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n560), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n553), .B(KEYINPUT13), .ZN(new_n570));
  OAI21_X1  g384(.A(G134), .B1(new_n570), .B2(new_n556), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n563), .B(new_n389), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n559), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NOR3_X1   g387(.A1(new_n437), .A2(new_n244), .A3(G953), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n569), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n574), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n567), .B1(new_n558), .B2(new_n559), .ZN(new_n577));
  AND3_X1   g391(.A1(new_n559), .A2(new_n571), .A3(new_n572), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n550), .B1(new_n580), .B2(new_n187), .ZN(new_n581));
  AOI211_X1 g395(.A(KEYINPUT92), .B(G902), .C1(new_n575), .C2(new_n579), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n549), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n580), .A2(new_n187), .ZN(new_n584));
  OR2_X1    g398(.A1(new_n584), .A2(new_n549), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n189), .A2(G952), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n586), .B1(G234), .B2(G237), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  XOR2_X1   g402(.A(KEYINPUT21), .B(G898), .Z(new_n589));
  NAND2_X1  g403(.A1(G234), .A2(G237), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n590), .A2(G902), .A3(G953), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n588), .B1(new_n589), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n583), .A2(new_n585), .A3(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(KEYINPUT93), .B1(new_n547), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n546), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n597), .B1(new_n541), .B2(KEYINPUT20), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT93), .ZN(new_n599));
  NOR4_X1   g413(.A1(new_n598), .A2(new_n599), .A3(new_n594), .A4(new_n528), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n379), .B(new_n482), .C1(new_n596), .C2(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(G101), .ZN(G3));
  OAI21_X1  g416(.A(KEYINPUT33), .B1(new_n574), .B2(KEYINPUT95), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n580), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n603), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n605), .B1(new_n575), .B2(new_n579), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n187), .A2(G478), .ZN(new_n607));
  NOR3_X1   g421(.A1(new_n604), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n584), .A2(KEYINPUT92), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n580), .A2(new_n550), .A3(new_n187), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n608), .B1(new_n548), .B2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n433), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n593), .B(new_n440), .C1(new_n613), .C2(new_n431), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n539), .B1(new_n525), .B2(new_n535), .ZN(new_n615));
  AOI211_X1 g429(.A(KEYINPUT89), .B(new_n534), .C1(new_n518), .C2(new_n524), .ZN(new_n616));
  NOR3_X1   g430(.A1(new_n615), .A2(new_n616), .A3(new_n543), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT20), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n546), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n528), .ZN(new_n620));
  AOI211_X1 g434(.A(new_n612), .B(new_n614), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n352), .A2(new_n187), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n252), .B1(new_n623), .B2(KEYINPUT94), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n624), .B1(KEYINPUT94), .B2(new_n623), .ZN(new_n625));
  AND2_X1   g439(.A1(new_n341), .A2(new_n354), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n246), .A2(new_n250), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n470), .A2(new_n444), .ZN(new_n629));
  INV_X1    g443(.A(new_n445), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n629), .A2(new_n479), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n438), .ZN(new_n632));
  OR2_X1    g446(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n622), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT34), .B(G104), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G6));
  NOR2_X1   g450(.A1(new_n615), .A2(new_n616), .ZN(new_n637));
  AOI22_X1  g451(.A1(new_n541), .A2(KEYINPUT20), .B1(new_n637), .B2(new_n544), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n583), .A2(new_n585), .ZN(new_n639));
  NOR4_X1   g453(.A1(new_n638), .A2(new_n639), .A3(new_n528), .A4(new_n614), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n641), .A2(new_n633), .ZN(new_n642));
  XNOR2_X1  g456(.A(KEYINPUT35), .B(G107), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G9));
  NAND3_X1  g458(.A1(new_n619), .A2(new_n620), .A3(new_n595), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n599), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n547), .A2(KEYINPUT93), .A3(new_n595), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n238), .A2(new_n243), .A3(new_n245), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n193), .A2(KEYINPUT36), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n239), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n247), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(KEYINPUT96), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT96), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n649), .A2(new_n655), .A3(new_n652), .ZN(new_n656));
  AND2_X1   g470(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  AND3_X1   g471(.A1(new_n657), .A2(new_n626), .A3(new_n625), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n648), .A2(new_n658), .A3(new_n482), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT37), .B(G110), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G12));
  NAND2_X1  g475(.A1(new_n654), .A2(new_n656), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n662), .B1(new_n357), .B2(new_n378), .ZN(new_n663));
  INV_X1    g477(.A(G900), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n587), .B1(new_n591), .B2(new_n664), .ZN(new_n665));
  NOR4_X1   g479(.A1(new_n638), .A2(new_n639), .A3(new_n528), .A4(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n441), .B1(new_n432), .B2(new_n433), .ZN(new_n667));
  INV_X1    g481(.A(new_n632), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n663), .A2(new_n666), .A3(new_n667), .A4(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G128), .ZN(G30));
  INV_X1    g484(.A(KEYINPUT40), .ZN(new_n671));
  XOR2_X1   g485(.A(new_n665), .B(KEYINPUT39), .Z(new_n672));
  NAND3_X1  g486(.A1(new_n631), .A2(new_n438), .A3(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT98), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n673), .A2(new_n674), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n671), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n677), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n679), .A2(KEYINPUT40), .A3(new_n675), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n434), .A2(new_n435), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT38), .ZN(new_n683));
  NOR4_X1   g497(.A1(new_n683), .A2(new_n547), .A3(new_n639), .A4(new_n441), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n314), .A2(new_n326), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n335), .A2(new_n296), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n252), .B1(new_n686), .B2(new_n329), .ZN(new_n687));
  AOI22_X1  g501(.A1(new_n685), .A2(new_n687), .B1(G472), .B2(G902), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(KEYINPUT97), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n653), .B1(new_n357), .B2(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n681), .A2(new_n684), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G143), .ZN(G45));
  AOI211_X1 g506(.A(new_n612), .B(new_n665), .C1(new_n619), .C2(new_n620), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n663), .A2(new_n693), .A3(new_n667), .A4(new_n668), .ZN(new_n694));
  XOR2_X1   g508(.A(KEYINPUT99), .B(G146), .Z(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G48));
  OR2_X1    g510(.A1(new_n470), .A2(new_n444), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n697), .A2(new_n629), .A3(new_n438), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(KEYINPUT100), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n379), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n700), .A2(new_n622), .ZN(new_n701));
  XOR2_X1   g515(.A(KEYINPUT41), .B(G113), .Z(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G15));
  NOR2_X1   g517(.A1(new_n700), .A2(new_n641), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(new_n561), .ZN(G18));
  NOR2_X1   g519(.A1(new_n596), .A2(new_n600), .ZN(new_n706));
  INV_X1    g520(.A(new_n667), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n707), .A2(new_n698), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n663), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g523(.A(KEYINPUT101), .B1(new_n706), .B2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT101), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n648), .A2(new_n711), .A3(new_n663), .A4(new_n708), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G119), .ZN(G21));
  NAND2_X1  g528(.A1(new_n583), .A2(new_n585), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n715), .B(new_n667), .C1(new_n598), .C2(new_n528), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT102), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n619), .A2(new_n620), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n719), .A2(KEYINPUT102), .A3(new_n715), .A4(new_n667), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n623), .A2(G472), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n340), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n251), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n593), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT100), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n698), .B(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n721), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G122), .ZN(G24));
  OR2_X1    g544(.A1(new_n604), .A2(new_n606), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n581), .A2(new_n582), .ZN(new_n732));
  OAI22_X1  g546(.A1(new_n731), .A2(new_n607), .B1(new_n732), .B2(G478), .ZN(new_n733));
  INV_X1    g547(.A(new_n665), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n719), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(new_n653), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n736), .A2(new_n723), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n708), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(new_n196), .ZN(G27));
  INV_X1    g554(.A(KEYINPUT42), .ZN(new_n741));
  AOI21_X1  g555(.A(KEYINPUT72), .B1(new_n376), .B2(G472), .ZN(new_n742));
  AOI211_X1 g556(.A(new_n358), .B(new_n252), .C1(new_n374), .C2(new_n375), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n355), .B(new_n356), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n436), .A2(new_n441), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n744), .A2(new_n745), .A3(new_n627), .A4(new_n668), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n741), .B1(new_n746), .B2(new_n735), .ZN(new_n747));
  NOR4_X1   g561(.A1(new_n436), .A2(new_n632), .A3(new_n741), .A4(new_n441), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n340), .A2(new_n342), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n356), .A2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT103), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n356), .A2(KEYINPUT103), .A3(new_n749), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n752), .A2(new_n378), .A3(new_n753), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n748), .A2(new_n693), .A3(new_n627), .A4(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n747), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G131), .ZN(G33));
  INV_X1    g571(.A(new_n666), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n746), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(new_n253), .ZN(G36));
  INV_X1    g574(.A(KEYINPUT104), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n619), .A2(new_n761), .A3(new_n620), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n619), .A2(new_n620), .A3(new_n733), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT43), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n547), .B(new_n733), .C1(new_n761), .C2(KEYINPUT43), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n736), .B1(new_n625), .B2(new_n626), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n767), .A2(KEYINPUT44), .A3(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n745), .B(KEYINPUT105), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n769), .A2(KEYINPUT106), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n767), .A2(new_n768), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT44), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n771), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(KEYINPUT106), .B1(new_n769), .B2(new_n770), .ZN(new_n776));
  OAI21_X1  g590(.A(KEYINPUT107), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n769), .A2(new_n770), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT106), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT107), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n780), .A2(new_n781), .A3(new_n774), .A4(new_n771), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n473), .A2(new_n478), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT45), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n473), .A2(new_n478), .A3(KEYINPUT45), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n785), .A2(G469), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n630), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT46), .ZN(new_n789));
  AOI22_X1  g603(.A1(new_n788), .A2(new_n789), .B1(new_n444), .B2(new_n470), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n444), .B1(new_n783), .B2(new_n784), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n445), .B1(new_n791), .B2(new_n786), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(KEYINPUT46), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n439), .B1(new_n790), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n672), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n777), .A2(new_n782), .A3(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(KEYINPUT108), .B(G137), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(KEYINPUT109), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n797), .B(new_n799), .ZN(G39));
  XOR2_X1   g614(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n788), .A2(new_n789), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n629), .B1(new_n792), .B2(KEYINPUT46), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n438), .B(new_n802), .C1(new_n803), .C2(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n805), .B1(new_n794), .B2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n745), .A2(new_n251), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n809), .A2(new_n735), .A3(new_n744), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G140), .ZN(G42));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n729), .A2(new_n659), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n379), .B(new_n699), .C1(new_n621), .C2(new_n640), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n436), .A2(new_n593), .A3(new_n480), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n816), .A2(new_n628), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n719), .A2(new_n639), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n547), .A2(new_n612), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n817), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n815), .A2(new_n601), .A3(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n814), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n638), .A2(new_n528), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT113), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n715), .A2(new_n665), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n744), .A2(new_n668), .A3(new_n657), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n824), .B1(new_n823), .B2(new_n825), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n693), .A2(new_n668), .A3(new_n737), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n745), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n759), .B1(new_n747), .B2(new_n755), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n822), .A2(new_n713), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n693), .A2(new_n708), .A3(new_n737), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n694), .A2(new_n669), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n357), .A2(new_n689), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n632), .A2(new_n665), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n836), .A2(new_n736), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n838), .B1(new_n720), .B2(new_n718), .ZN(new_n839));
  OAI21_X1  g653(.A(KEYINPUT52), .B1(new_n835), .B2(new_n839), .ZN(new_n840));
  AND4_X1   g654(.A1(new_n744), .A2(new_n667), .A3(new_n657), .A4(new_n668), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n739), .B1(new_n666), .B2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT52), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n721), .A2(new_n690), .A3(new_n837), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n842), .A2(new_n843), .A3(new_n844), .A4(new_n694), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n840), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n813), .B1(new_n833), .B2(new_n846), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n840), .A2(new_n845), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n815), .A2(new_n601), .A3(new_n820), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n481), .B1(new_n646), .B2(new_n647), .ZN(new_n850));
  AOI22_X1  g664(.A1(new_n850), .A2(new_n658), .B1(new_n721), .B2(new_n728), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n713), .A2(new_n849), .A3(new_n851), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n831), .A2(new_n832), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n848), .A2(KEYINPUT53), .A3(new_n852), .A4(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(KEYINPUT114), .B1(new_n847), .B2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT114), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n713), .A2(new_n849), .A3(new_n851), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n831), .A2(new_n832), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(new_n848), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n856), .B1(new_n860), .B2(new_n813), .ZN(new_n861));
  OAI21_X1  g675(.A(KEYINPUT54), .B1(new_n855), .B2(new_n861), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n586), .B(KEYINPUT118), .ZN(new_n863));
  INV_X1    g677(.A(new_n698), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n745), .A2(new_n627), .A3(new_n587), .A4(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n865), .A2(new_n836), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n863), .B1(new_n866), .B2(new_n819), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n767), .A2(new_n587), .A3(new_n864), .A4(new_n724), .ZN(new_n868));
  AND4_X1   g682(.A1(new_n587), .A2(new_n767), .A3(new_n864), .A4(new_n745), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n754), .A2(new_n627), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n871), .A2(KEYINPUT48), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n871), .A2(KEYINPUT48), .ZN(new_n873));
  OAI221_X1 g687(.A(new_n867), .B1(new_n707), .B2(new_n868), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT115), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n807), .A2(new_n875), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n805), .B(KEYINPUT115), .C1(new_n794), .C2(new_n806), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n697), .A2(new_n629), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n878), .A2(new_n438), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n876), .A2(new_n877), .A3(new_n880), .ZN(new_n881));
  AND4_X1   g695(.A1(new_n587), .A2(new_n770), .A3(new_n767), .A4(new_n724), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT51), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT116), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n886), .A2(KEYINPUT50), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n683), .B(new_n441), .C1(new_n886), .C2(KEYINPUT50), .ZN(new_n888));
  OR3_X1    g702(.A1(new_n868), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n887), .B1(new_n868), .B2(new_n888), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI22_X1  g705(.A1(new_n885), .A2(new_n891), .B1(KEYINPUT117), .B2(new_n884), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n719), .A2(new_n733), .ZN(new_n893));
  AOI22_X1  g707(.A1(new_n869), .A2(new_n737), .B1(new_n866), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n882), .B1(new_n808), .B2(new_n879), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT117), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n896), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(KEYINPUT51), .B1(new_n898), .B2(new_n891), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n874), .B1(new_n895), .B2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT54), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n847), .A2(new_n854), .A3(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n862), .A2(new_n900), .A3(new_n903), .ZN(new_n904));
  OR2_X1    g718(.A1(G952), .A2(G953), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n627), .A2(new_n442), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT111), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n908), .A2(new_n547), .A3(new_n733), .ZN(new_n909));
  OR2_X1    g723(.A1(new_n909), .A2(KEYINPUT112), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(KEYINPUT112), .ZN(new_n911));
  INV_X1    g725(.A(new_n683), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n878), .B(KEYINPUT49), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n912), .A2(new_n836), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n910), .A2(new_n911), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n906), .A2(new_n915), .ZN(G75));
  NOR2_X1   g730(.A1(new_n189), .A2(G952), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n187), .B1(new_n847), .B2(new_n854), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT56), .B1(new_n919), .B2(G210), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n428), .A2(new_n429), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(new_n424), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n922), .B(KEYINPUT55), .Z(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n918), .B1(new_n920), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n925), .B1(new_n920), .B2(new_n924), .ZN(G51));
  XNOR2_X1  g740(.A(new_n445), .B(KEYINPUT57), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n901), .B1(new_n847), .B2(new_n854), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n927), .B1(new_n902), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n460), .A2(new_n469), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n919), .A2(new_n786), .A3(new_n791), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n917), .B1(new_n931), .B2(new_n932), .ZN(G54));
  AND2_X1   g747(.A1(KEYINPUT58), .A2(G475), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n919), .A2(new_n934), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n935), .A2(new_n615), .A3(new_n616), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n637), .B1(new_n919), .B2(new_n934), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n936), .A2(new_n917), .A3(new_n937), .ZN(G60));
  XNOR2_X1  g752(.A(new_n731), .B(KEYINPUT119), .ZN(new_n939));
  NAND2_X1  g753(.A1(G478), .A2(G902), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT59), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n939), .B(new_n941), .C1(new_n902), .C2(new_n928), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n918), .ZN(new_n943));
  AOI21_X1  g757(.A(KEYINPUT53), .B1(new_n859), .B2(new_n848), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n833), .A2(new_n813), .A3(new_n846), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n856), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n847), .A2(KEYINPUT114), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n901), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n941), .B1(new_n948), .B2(new_n902), .ZN(new_n949));
  INV_X1    g763(.A(new_n939), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n943), .B1(new_n949), .B2(new_n950), .ZN(G63));
  XNOR2_X1  g765(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n952));
  NAND2_X1  g766(.A1(G217), .A2(G902), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT121), .Z(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT122), .ZN(new_n955));
  XNOR2_X1  g769(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n957), .B1(new_n944), .B2(new_n945), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n232), .A2(new_n236), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n917), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(new_n651), .ZN(new_n961));
  INV_X1    g775(.A(new_n957), .ZN(new_n962));
  AOI211_X1 g776(.A(new_n961), .B(new_n962), .C1(new_n847), .C2(new_n854), .ZN(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n952), .B1(new_n960), .B2(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n962), .B1(new_n847), .B2(new_n854), .ZN(new_n966));
  INV_X1    g780(.A(new_n959), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n918), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(new_n952), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n968), .A2(new_n969), .A3(new_n963), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n965), .A2(new_n970), .ZN(G66));
  AOI21_X1  g785(.A(KEYINPUT124), .B1(new_n822), .B2(new_n713), .ZN(new_n972));
  AND4_X1   g786(.A1(KEYINPUT124), .A2(new_n713), .A3(new_n849), .A4(new_n851), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(new_n189), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n589), .A2(G224), .A3(G953), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n921), .B1(G898), .B2(new_n189), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n977), .B(new_n978), .Z(G69));
  NAND2_X1  g793(.A1(G227), .A2(G900), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n664), .A2(G953), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(KEYINPUT126), .Z(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n759), .B1(new_n808), .B2(new_n810), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n796), .A2(new_n721), .A3(new_n870), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n984), .A2(new_n756), .A3(new_n985), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n986), .A2(new_n835), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n797), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n983), .B1(new_n988), .B2(new_n189), .ZN(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n323), .A2(new_n325), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(KEYINPUT125), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n992), .B(new_n532), .ZN(new_n993));
  OAI211_X1 g807(.A(G953), .B(new_n980), .C1(new_n990), .C2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(new_n691), .ZN(new_n995));
  OAI21_X1  g809(.A(KEYINPUT62), .B1(new_n995), .B2(new_n835), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT62), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n691), .A2(new_n842), .A3(new_n997), .A4(new_n694), .ZN(new_n998));
  OR2_X1    g812(.A1(new_n818), .A2(new_n819), .ZN(new_n999));
  AND4_X1   g813(.A1(new_n379), .A2(new_n675), .A3(new_n679), .A4(new_n745), .ZN(new_n1000));
  AOI22_X1  g814(.A1(new_n808), .A2(new_n810), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  AND3_X1   g815(.A1(new_n996), .A2(new_n998), .A3(new_n1001), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n797), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n993), .B1(new_n1003), .B2(G953), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n980), .A2(G953), .ZN(new_n1005));
  OAI211_X1 g819(.A(new_n1004), .B(new_n1005), .C1(new_n993), .C2(new_n989), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n994), .A2(new_n1006), .ZN(G72));
  INV_X1    g821(.A(KEYINPUT127), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n797), .A2(new_n974), .A3(new_n1002), .ZN(new_n1009));
  NAND2_X1  g823(.A1(G472), .A2(G902), .ZN(new_n1010));
  XOR2_X1   g824(.A(new_n1010), .B(KEYINPUT63), .Z(new_n1011));
  NAND2_X1  g825(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n371), .A2(new_n329), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1008), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g828(.A(new_n1013), .ZN(new_n1015));
  AOI211_X1 g829(.A(KEYINPUT127), .B(new_n1015), .C1(new_n1009), .C2(new_n1011), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n797), .A2(new_n974), .A3(new_n987), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1018), .A2(new_n1011), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n1019), .A2(new_n329), .A3(new_n371), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n366), .A2(new_n685), .ZN(new_n1021));
  OAI211_X1 g835(.A(new_n1011), .B(new_n1021), .C1(new_n855), .C2(new_n861), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n1020), .A2(new_n1022), .A3(new_n918), .ZN(new_n1023));
  NOR2_X1   g837(.A1(new_n1017), .A2(new_n1023), .ZN(G57));
endmodule


