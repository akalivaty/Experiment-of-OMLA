//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 0 0 0 0 1 1 1 0 1 0 0 0 1 1 0 0 1 1 1 0 0 0 0 1 0 0 0 1 0 1 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 1 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:26 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1237,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT64), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  INV_X1    g0005(.A(G264), .ZN(new_n206));
  INV_X1    g0006(.A(G116), .ZN(new_n207));
  INV_X1    g0007(.A(G270), .ZN(new_n208));
  OAI22_X1  g0008(.A1(new_n205), .A2(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(G68), .ZN(new_n210));
  INV_X1    g0010(.A(G238), .ZN(new_n211));
  INV_X1    g0011(.A(G87), .ZN(new_n212));
  INV_X1    g0012(.A(G250), .ZN(new_n213));
  OAI22_X1  g0013(.A1(new_n210), .A2(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g0014(.A(KEYINPUT66), .B(G244), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n209), .B(new_n214), .C1(G77), .C2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G58), .ZN(new_n217));
  INV_X1    g0017(.A(G232), .ZN(new_n218));
  INV_X1    g0018(.A(G97), .ZN(new_n219));
  INV_X1    g0019(.A(G257), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G50), .ZN(new_n222));
  INV_X1    g0022(.A(G226), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n204), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT1), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n204), .A2(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT0), .Z(new_n229));
  OR2_X1    g0029(.A1(KEYINPUT65), .A2(G20), .ZN(new_n230));
  NAND2_X1  g0030(.A1(KEYINPUT65), .A2(G20), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n217), .A2(new_n210), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n233), .A2(G50), .ZN(new_n234));
  NAND2_X1  g0034(.A1(G1), .A2(G13), .ZN(new_n235));
  NOR3_X1   g0035(.A1(new_n232), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  NOR3_X1   g0036(.A1(new_n226), .A2(new_n229), .A3(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(new_n218), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G264), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(new_n208), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G358));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT67), .ZN(new_n247));
  XOR2_X1   g0047(.A(G68), .B(G77), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G87), .B(G97), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G107), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  INV_X1    g0053(.A(KEYINPUT77), .ZN(new_n254));
  INV_X1    g0054(.A(G1), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G20), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n256), .B(KEYINPUT71), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT74), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n255), .A2(G13), .A3(G20), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(new_n235), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n258), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  NAND4_X1  g0063(.A1(new_n259), .A2(KEYINPUT74), .A3(new_n235), .A4(new_n261), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n257), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G68), .ZN(new_n266));
  NAND4_X1  g0066(.A1(new_n255), .A2(new_n210), .A3(G13), .A4(G20), .ZN(new_n267));
  XNOR2_X1  g0067(.A(new_n267), .B(KEYINPUT12), .ZN(new_n268));
  NOR2_X1   g0068(.A1(G20), .A2(G33), .ZN(new_n269));
  AOI22_X1  g0069(.A1(new_n269), .A2(G50), .B1(G20), .B2(new_n210), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n232), .A2(G33), .ZN(new_n271));
  INV_X1    g0071(.A(G77), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT70), .ZN(new_n274));
  AND3_X1   g0074(.A1(new_n261), .A2(new_n274), .A3(new_n235), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n274), .B1(new_n261), .B2(new_n235), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  AND2_X1   g0078(.A1(new_n278), .A2(KEYINPUT11), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n278), .A2(KEYINPUT11), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n266), .B(new_n268), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G169), .ZN(new_n283));
  INV_X1    g0083(.A(G33), .ZN(new_n284));
  INV_X1    g0084(.A(G41), .ZN(new_n285));
  OAI211_X1 g0085(.A(G1), .B(G13), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n255), .B1(G41), .B2(G45), .ZN(new_n287));
  AND2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G238), .ZN(new_n289));
  INV_X1    g0089(.A(G274), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G226), .A2(G1698), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n293), .B1(new_n218), .B2(G1698), .ZN(new_n294));
  XNOR2_X1  g0094(.A(KEYINPUT3), .B(G33), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT75), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n296), .A2(G33), .A3(G97), .ZN(new_n297));
  NAND2_X1  g0097(.A1(G33), .A2(G97), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(KEYINPUT75), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n294), .A2(new_n295), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n289), .B(new_n292), .C1(new_n286), .C2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT13), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n294), .A2(new_n295), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n299), .A2(new_n297), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n235), .B1(G33), .B2(G41), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n291), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT13), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n307), .A2(new_n308), .A3(new_n289), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n283), .B1(new_n302), .B2(new_n309), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n310), .B(KEYINPUT14), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n302), .A2(new_n309), .A3(KEYINPUT76), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT76), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n301), .A2(new_n313), .A3(KEYINPUT13), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G179), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n282), .B1(new_n311), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n315), .A2(G190), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n302), .A2(new_n309), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G200), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n318), .A2(new_n282), .A3(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n254), .B1(new_n317), .B2(new_n322), .ZN(new_n323));
  NOR2_X1   g0123(.A1(G222), .A2(G1698), .ZN(new_n324));
  INV_X1    g0124(.A(G1698), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n325), .A2(G223), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n295), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n327), .B1(G77), .B2(new_n295), .ZN(new_n328));
  OR2_X1    g0128(.A1(new_n328), .A2(KEYINPUT69), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(KEYINPUT69), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n329), .A2(new_n306), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n286), .A2(new_n287), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n292), .B1(new_n332), .B2(new_n223), .ZN(new_n333));
  XNOR2_X1  g0133(.A(new_n333), .B(KEYINPUT68), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n335), .A2(G179), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n336), .B1(new_n283), .B2(new_n335), .ZN(new_n337));
  OAI21_X1  g0137(.A(G20), .B1(new_n233), .B2(G50), .ZN(new_n338));
  INV_X1    g0138(.A(G150), .ZN(new_n339));
  INV_X1    g0139(.A(new_n269), .ZN(new_n340));
  XNOR2_X1  g0140(.A(KEYINPUT8), .B(G58), .ZN(new_n341));
  OAI221_X1 g0141(.A(new_n338), .B1(new_n339), .B2(new_n340), .C1(new_n271), .C2(new_n341), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n342), .A2(new_n277), .B1(new_n222), .B2(new_n260), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n277), .A2(new_n260), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n257), .A2(new_n222), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n337), .A2(new_n347), .ZN(new_n348));
  OAI22_X1  g0148(.A1(new_n232), .A2(new_n272), .B1(new_n341), .B2(new_n340), .ZN(new_n349));
  XNOR2_X1  g0149(.A(new_n349), .B(KEYINPUT72), .ZN(new_n350));
  XOR2_X1   g0150(.A(KEYINPUT15), .B(G87), .Z(new_n351));
  OR2_X1    g0151(.A1(new_n351), .A2(KEYINPUT73), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(KEYINPUT73), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n350), .B1(new_n271), .B2(new_n354), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n355), .A2(new_n262), .B1(new_n272), .B2(new_n260), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n265), .A2(G77), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(G238), .A2(G1698), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n295), .B(new_n359), .C1(new_n218), .C2(G1698), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n360), .B(new_n306), .C1(G107), .C2(new_n295), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n288), .A2(new_n215), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n361), .A2(new_n292), .A3(new_n362), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n363), .A2(G179), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n364), .B1(new_n283), .B2(new_n363), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n358), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n363), .A2(G200), .ZN(new_n367));
  INV_X1    g0167(.A(G190), .ZN(new_n368));
  OR2_X1    g0168(.A1(new_n363), .A2(new_n368), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n356), .A2(new_n357), .A3(new_n367), .A4(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  AND3_X1   g0172(.A1(new_n323), .A2(new_n348), .A3(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT79), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT7), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n284), .A2(KEYINPUT3), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT3), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(G33), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT78), .ZN(new_n379));
  AND3_X1   g0179(.A1(new_n376), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n379), .B1(new_n376), .B2(new_n378), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n375), .B(new_n232), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(KEYINPUT7), .B1(new_n295), .B2(G20), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n382), .A2(G68), .A3(new_n383), .ZN(new_n384));
  XNOR2_X1  g0184(.A(G58), .B(G68), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n385), .A2(G20), .B1(G159), .B2(new_n269), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n384), .A2(KEYINPUT16), .A3(new_n386), .ZN(new_n387));
  AND2_X1   g0187(.A1(KEYINPUT65), .A2(G20), .ZN(new_n388));
  NOR2_X1   g0188(.A1(KEYINPUT65), .A2(G20), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(KEYINPUT7), .B1(new_n390), .B2(new_n295), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n376), .A2(new_n378), .ZN(new_n392));
  INV_X1    g0192(.A(G20), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n392), .A2(new_n375), .A3(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n391), .A2(G68), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n386), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT16), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n387), .A2(new_n398), .A3(new_n262), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n257), .A2(new_n341), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n344), .A2(new_n400), .B1(new_n260), .B2(new_n341), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  OR2_X1    g0202(.A1(G223), .A2(G1698), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n223), .A2(G1698), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n295), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G33), .A2(G87), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n306), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n291), .B1(new_n288), .B2(G232), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n408), .A2(G179), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n286), .B1(new_n405), .B2(new_n406), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n292), .B1(new_n332), .B2(new_n218), .ZN(new_n412));
  OAI21_X1  g0212(.A(G169), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n402), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT18), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n411), .A2(new_n412), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n368), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(G200), .B2(new_n417), .ZN(new_n419));
  AND3_X1   g0219(.A1(new_n399), .A2(new_n419), .A3(new_n401), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(KEYINPUT17), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT18), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n402), .A2(new_n414), .A3(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n399), .A2(new_n419), .A3(new_n401), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT17), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n416), .A2(new_n421), .A3(new_n423), .A4(new_n426), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n317), .A2(new_n322), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n427), .B1(new_n428), .B2(KEYINPUT77), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT9), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n335), .A2(G200), .B1(new_n430), .B2(new_n347), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n343), .A2(KEYINPUT9), .A3(new_n346), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n331), .A2(G190), .A3(new_n334), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  XNOR2_X1  g0234(.A(new_n434), .B(KEYINPUT10), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n373), .A2(new_n374), .A3(new_n429), .A4(new_n435), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n323), .A2(new_n435), .A3(new_n348), .A4(new_n372), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n416), .A2(new_n423), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  AND2_X1   g0239(.A1(new_n421), .A2(new_n426), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT14), .ZN(new_n441));
  XNOR2_X1  g0241(.A(new_n310), .B(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n316), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n281), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n321), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n439), .B(new_n440), .C1(new_n445), .C2(new_n254), .ZN(new_n446));
  OAI21_X1  g0246(.A(KEYINPUT79), .B1(new_n437), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n436), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT23), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n230), .A2(new_n449), .A3(new_n205), .A4(new_n231), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n284), .A2(new_n207), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n393), .ZN(new_n452));
  OAI21_X1  g0252(.A(KEYINPUT23), .B1(new_n393), .B2(G107), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n450), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n376), .B(new_n378), .C1(new_n388), .C2(new_n389), .ZN(new_n455));
  OAI21_X1  g0255(.A(KEYINPUT22), .B1(new_n455), .B2(new_n212), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT22), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n232), .A2(new_n295), .A3(new_n457), .A4(G87), .ZN(new_n458));
  AOI211_X1 g0258(.A(KEYINPUT24), .B(new_n454), .C1(new_n456), .C2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT24), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n456), .A2(new_n458), .ZN(new_n461));
  INV_X1    g0261(.A(new_n454), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n262), .B1(new_n459), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT81), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n465), .B1(new_n284), .B2(G1), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n255), .A2(KEYINPUT81), .A3(G33), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n259), .B(new_n468), .C1(new_n275), .C2(new_n276), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G107), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n259), .A2(G107), .ZN(new_n472));
  XNOR2_X1  g0272(.A(new_n472), .B(KEYINPUT25), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n464), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n213), .A2(new_n325), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n220), .A2(G1698), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n376), .A2(new_n475), .A3(new_n378), .A4(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(G294), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n477), .B1(new_n284), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n255), .A2(G45), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT82), .ZN(new_n481));
  OAI21_X1  g0281(.A(KEYINPUT5), .B1(new_n481), .B2(G41), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT5), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n483), .A2(new_n285), .A3(KEYINPUT82), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n480), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n479), .A2(new_n306), .B1(G274), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n482), .A2(new_n484), .ZN(new_n487));
  INV_X1    g0287(.A(new_n480), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n306), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(G264), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(KEYINPUT90), .B1(new_n489), .B2(G264), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT90), .ZN(new_n494));
  NOR4_X1   g0294(.A1(new_n485), .A2(new_n494), .A3(new_n306), .A4(new_n206), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n486), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(G200), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n492), .A2(new_n368), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n474), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT89), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n474), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n464), .A2(KEYINPUT89), .A3(new_n471), .A4(new_n473), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(G179), .ZN(new_n504));
  OAI22_X1  g0304(.A1(new_n492), .A2(new_n283), .B1(new_n496), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n499), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(G33), .B(G97), .C1(new_n388), .C2(new_n389), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  OAI21_X1  g0308(.A(KEYINPUT84), .B1(new_n508), .B2(KEYINPUT19), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n299), .A2(new_n297), .A3(KEYINPUT19), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n232), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n212), .A2(new_n219), .A3(new_n205), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n232), .A2(new_n295), .A3(G68), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT84), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT19), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n507), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n509), .A2(new_n513), .A3(new_n514), .A4(new_n517), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n518), .A2(new_n262), .B1(new_n260), .B2(new_n354), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n470), .A2(new_n352), .A3(new_n353), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(KEYINPUT85), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n488), .A2(G274), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n286), .A2(G250), .A3(new_n480), .ZN(new_n524));
  NAND2_X1  g0324(.A1(G244), .A2(G1698), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(new_n211), .B2(G1698), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n451), .B1(new_n295), .B2(new_n526), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n523), .B(new_n524), .C1(new_n527), .C2(new_n286), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n528), .A2(new_n504), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(G169), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT85), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n519), .A2(new_n533), .A3(new_n520), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n522), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n518), .A2(new_n262), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n354), .A2(new_n260), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n470), .A2(G87), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n528), .A2(G200), .ZN(new_n541));
  OR2_X1    g0341(.A1(new_n528), .A2(new_n368), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AND2_X1   g0343(.A1(new_n535), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n284), .A2(G97), .ZN(new_n545));
  NAND2_X1  g0345(.A1(G33), .A2(G283), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n545), .B(new_n546), .C1(new_n388), .C2(new_n389), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n261), .A2(new_n235), .B1(G20), .B2(new_n207), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT20), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n547), .A2(KEYINPUT20), .A3(new_n548), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n551), .A2(KEYINPUT87), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n263), .A2(new_n264), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n554), .A2(G116), .A3(new_n468), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n255), .A2(new_n207), .A3(G13), .A4(G20), .ZN(new_n556));
  XOR2_X1   g0356(.A(new_n556), .B(KEYINPUT86), .Z(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT87), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n549), .A2(new_n559), .A3(new_n550), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n553), .A2(new_n555), .A3(new_n558), .A4(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT88), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n487), .A2(new_n488), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n564), .A2(G270), .A3(new_n286), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n485), .A2(G274), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n325), .A2(G257), .ZN(new_n567));
  NAND2_X1  g0367(.A1(G264), .A2(G1698), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n376), .A2(new_n378), .A3(new_n567), .A4(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n569), .B(new_n306), .C1(G303), .C2(new_n295), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n565), .A2(new_n566), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(G200), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n565), .A2(new_n570), .A3(G190), .A4(new_n566), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n562), .A2(new_n563), .A3(new_n572), .A4(new_n573), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n263), .A2(new_n264), .B1(new_n466), .B2(new_n467), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n557), .B1(new_n575), .B2(G116), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n576), .A2(new_n560), .A3(new_n573), .A4(new_n553), .ZN(new_n577));
  INV_X1    g0377(.A(new_n572), .ZN(new_n578));
  OAI21_X1  g0378(.A(KEYINPUT88), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n574), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n561), .A2(G169), .A3(new_n571), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(KEYINPUT21), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT21), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n561), .A2(new_n583), .A3(G169), .A4(new_n571), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n562), .A2(new_n571), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(G179), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n580), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n376), .A2(new_n378), .A3(G244), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT4), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n590), .A2(G1698), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n592), .A2(new_n376), .A3(new_n378), .A4(G244), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n591), .A2(new_n546), .A3(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n376), .A2(new_n378), .A3(G250), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n325), .B1(new_n595), .B2(KEYINPUT4), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n306), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n489), .A2(G257), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n599), .A2(KEYINPUT83), .A3(new_n504), .A4(new_n566), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n469), .A2(new_n219), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n391), .A2(G107), .A3(new_n394), .ZN(new_n602));
  XOR2_X1   g0402(.A(KEYINPUT80), .B(G107), .Z(new_n603));
  OR2_X1    g0403(.A1(KEYINPUT6), .A2(G97), .ZN(new_n604));
  OAI21_X1  g0404(.A(KEYINPUT6), .B1(G97), .B2(G107), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g0407(.A(KEYINPUT80), .B(G107), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n608), .A2(new_n605), .A3(new_n604), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n607), .A2(new_n390), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n269), .A2(G77), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n602), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n601), .B1(new_n612), .B2(new_n262), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(G97), .B2(new_n259), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT83), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n597), .A2(new_n566), .A3(new_n598), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n615), .B1(new_n616), .B2(G179), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n283), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n600), .A2(new_n614), .A3(new_n617), .A4(new_n618), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n259), .A2(G97), .ZN(new_n620));
  AOI211_X1 g0420(.A(new_n620), .B(new_n601), .C1(new_n612), .C2(new_n262), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n616), .A2(G200), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n597), .A2(G190), .A3(new_n566), .A4(new_n598), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n619), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n588), .A2(new_n625), .ZN(new_n626));
  AND4_X1   g0426(.A1(new_n448), .A2(new_n506), .A3(new_n544), .A4(new_n626), .ZN(G372));
  NAND2_X1  g0427(.A1(new_n541), .A2(KEYINPUT91), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT91), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n528), .A2(new_n629), .A3(G200), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n628), .A2(new_n542), .A3(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n539), .A2(new_n631), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n519), .A2(new_n520), .B1(new_n531), .B2(new_n530), .ZN(new_n633));
  OAI21_X1  g0433(.A(KEYINPUT92), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n521), .A2(new_n532), .ZN(new_n635));
  INV_X1    g0435(.A(new_n528), .ZN(new_n636));
  AOI22_X1  g0436(.A1(KEYINPUT91), .A2(new_n541), .B1(new_n636), .B2(G190), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n637), .A2(new_n519), .A3(new_n538), .A4(new_n630), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT92), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n635), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(KEYINPUT26), .B1(new_n634), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n624), .B1(new_n474), .B2(new_n498), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n582), .A2(new_n584), .B1(new_n586), .B2(G179), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n474), .A2(new_n505), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n642), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n619), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n641), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n646), .A2(new_n535), .A3(new_n543), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n633), .B1(new_n648), .B2(KEYINPUT26), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n448), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT93), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n435), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n435), .A2(new_n652), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n444), .B1(new_n322), .B2(new_n366), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n438), .B1(new_n656), .B2(new_n440), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n348), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n651), .A2(new_n659), .ZN(G369));
  INV_X1    g0460(.A(new_n505), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n661), .B1(new_n501), .B2(new_n502), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n232), .A2(G13), .ZN(new_n663));
  OAI21_X1  g0463(.A(KEYINPUT27), .B1(new_n663), .B2(G1), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT27), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n232), .A2(new_n665), .A3(new_n255), .A4(G13), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n664), .A2(G213), .A3(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(G343), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AOI211_X1 g0469(.A(new_n499), .B(new_n662), .C1(new_n503), .C2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n503), .A2(new_n505), .ZN(new_n671));
  INV_X1    g0471(.A(new_n669), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n585), .A2(new_n587), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n562), .A2(new_n672), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n588), .B2(new_n676), .ZN(new_n678));
  XOR2_X1   g0478(.A(KEYINPUT94), .B(G330), .Z(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n674), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n675), .A2(new_n672), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT95), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n684), .B1(new_n670), .B2(new_n673), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n644), .A2(new_n669), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n682), .A2(new_n688), .ZN(G399));
  INV_X1    g0489(.A(new_n227), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(G41), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n512), .A2(G116), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(G1), .A3(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n694), .B1(new_n234), .B2(new_n692), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n695), .B(KEYINPUT28), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n626), .A2(new_n506), .A3(new_n544), .A4(new_n672), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT98), .ZN(new_n698));
  AND3_X1   g0498(.A1(new_n616), .A2(new_n698), .A3(new_n496), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n698), .B1(new_n616), .B2(new_n496), .ZN(new_n700));
  OAI211_X1 g0500(.A(new_n504), .B(new_n528), .C1(new_n699), .C2(new_n700), .ZN(new_n701));
  AND3_X1   g0501(.A1(new_n565), .A2(new_n566), .A3(new_n570), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n493), .A2(new_n495), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n616), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n571), .B1(new_n306), .B2(new_n479), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n705), .A2(new_n529), .A3(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT97), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(KEYINPUT30), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n709), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n705), .A2(new_n529), .A3(new_n711), .A4(new_n706), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n669), .B1(new_n703), .B2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT31), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  XOR2_X1   g0516(.A(KEYINPUT96), .B(KEYINPUT31), .Z(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n697), .B(new_n716), .C1(new_n714), .C2(new_n718), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n719), .A2(new_n679), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n634), .A2(new_n640), .ZN(new_n721));
  INV_X1    g0521(.A(new_n642), .ZN(new_n722));
  OAI211_X1 g0522(.A(new_n721), .B(new_n722), .C1(new_n662), .C2(new_n675), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT26), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n646), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n646), .A2(new_n535), .A3(new_n724), .A4(new_n543), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n634), .A2(new_n640), .A3(KEYINPUT26), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n726), .A2(new_n727), .A3(new_n635), .ZN(new_n728));
  OAI211_X1 g0528(.A(KEYINPUT29), .B(new_n672), .C1(new_n725), .C2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(KEYINPUT99), .ZN(new_n730));
  INV_X1    g0530(.A(new_n728), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n671), .A2(new_n643), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n642), .B1(new_n634), .B2(new_n640), .ZN(new_n733));
  AOI21_X1  g0533(.A(KEYINPUT26), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n731), .B1(new_n734), .B2(new_n646), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT99), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n735), .A2(new_n736), .A3(KEYINPUT29), .A4(new_n672), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n730), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n669), .B1(new_n647), .B2(new_n649), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(KEYINPUT29), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n720), .B1(new_n738), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n696), .B1(new_n742), .B2(G1), .ZN(G364));
  AOI21_X1  g0543(.A(new_n235), .B1(G20), .B2(new_n283), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n232), .A2(G190), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n746), .A2(G179), .A3(new_n497), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n295), .B1(new_n747), .B2(new_n272), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT100), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  NOR3_X1   g0550(.A1(new_n232), .A2(KEYINPUT100), .A3(G190), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n497), .A2(G179), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n205), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n746), .A2(G179), .A3(G200), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI211_X1 g0559(.A(new_n748), .B(new_n757), .C1(G68), .C2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G179), .A2(G200), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G190), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n390), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n219), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n232), .A2(new_n504), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n766), .A2(G190), .A3(G200), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n754), .A2(new_n393), .A3(new_n368), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n767), .A2(new_n222), .B1(new_n769), .B2(new_n212), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n766), .A2(G190), .A3(new_n497), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI211_X1 g0572(.A(new_n765), .B(new_n770), .C1(G58), .C2(new_n772), .ZN(new_n773));
  NOR3_X1   g0573(.A1(new_n752), .A2(G179), .A3(G200), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(G159), .ZN(new_n776));
  OAI21_X1  g0576(.A(KEYINPUT32), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OR3_X1    g0577(.A1(new_n775), .A2(KEYINPUT32), .A3(new_n776), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n760), .A2(new_n773), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n774), .A2(G329), .B1(new_n755), .B2(G283), .ZN(new_n780));
  INV_X1    g0580(.A(G322), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n771), .A2(new_n781), .ZN(new_n782));
  XOR2_X1   g0582(.A(KEYINPUT33), .B(G317), .Z(new_n783));
  OAI21_X1  g0583(.A(new_n392), .B1(new_n758), .B2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n767), .ZN(new_n785));
  XOR2_X1   g0585(.A(KEYINPUT101), .B(G326), .Z(new_n786));
  AOI211_X1 g0586(.A(new_n782), .B(new_n784), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n747), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G311), .ZN(new_n789));
  AND3_X1   g0589(.A1(new_n780), .A2(new_n787), .A3(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G303), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n790), .B1(new_n478), .B2(new_n764), .C1(new_n791), .C2(new_n769), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n745), .B1(new_n779), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(G13), .A2(G33), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(G20), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n744), .ZN(new_n797));
  OR2_X1    g0597(.A1(new_n380), .A2(new_n381), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(new_n690), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(G45), .B2(new_n234), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n801), .B1(G45), .B2(new_n249), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n802), .B1(new_n207), .B2(new_n690), .ZN(new_n803));
  INV_X1    g0603(.A(G355), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n227), .A2(new_n295), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n793), .B1(new_n797), .B2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n663), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(G45), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(G1), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n691), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n796), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n807), .B(new_n811), .C1(new_n678), .C2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n811), .B1(new_n678), .B2(new_n679), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n814), .B1(new_n679), .B2(new_n678), .ZN(new_n815));
  AND2_X1   g0615(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(G396));
  NAND2_X1  g0617(.A1(new_n358), .A2(new_n669), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(new_n370), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(new_n366), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n366), .A2(new_n669), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n739), .B(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n824), .A2(new_n720), .ZN(new_n825));
  XOR2_X1   g0625(.A(new_n825), .B(KEYINPUT104), .Z(new_n826));
  AOI21_X1  g0626(.A(new_n811), .B1(new_n824), .B2(new_n720), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n755), .A2(G87), .B1(G294), .B2(new_n772), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(new_n205), .B2(new_n769), .ZN(new_n830));
  OR3_X1    g0630(.A1(new_n830), .A2(new_n295), .A3(new_n765), .ZN(new_n831));
  INV_X1    g0631(.A(G283), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n207), .A2(new_n747), .B1(new_n758), .B2(new_n832), .ZN(new_n833));
  OR2_X1    g0633(.A1(new_n833), .A2(KEYINPUT102), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(KEYINPUT102), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n834), .B(new_n835), .C1(new_n791), .C2(new_n767), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n836), .B(KEYINPUT103), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n831), .B(new_n837), .C1(G311), .C2(new_n774), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n772), .A2(G143), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n788), .A2(G159), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n785), .A2(G137), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n759), .A2(G150), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n839), .A2(new_n840), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT34), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(G132), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n845), .B(new_n799), .C1(new_n846), .C2(new_n775), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n764), .A2(new_n217), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n756), .A2(new_n210), .ZN(new_n849));
  OAI22_X1  g0649(.A1(new_n843), .A2(new_n844), .B1(new_n222), .B2(new_n769), .ZN(new_n850));
  NOR4_X1   g0650(.A1(new_n847), .A2(new_n848), .A3(new_n849), .A4(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n744), .B1(new_n838), .B2(new_n851), .ZN(new_n852));
  AND2_X1   g0652(.A1(new_n852), .A2(new_n811), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n744), .A2(new_n794), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n823), .ZN(new_n856));
  OAI221_X1 g0656(.A(new_n853), .B1(G77), .B2(new_n855), .C1(new_n795), .C2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n828), .A2(new_n857), .ZN(G384));
  INV_X1    g0658(.A(KEYINPUT38), .ZN(new_n859));
  AND3_X1   g0659(.A1(new_n410), .A2(new_n413), .A3(new_n667), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n402), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT37), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n862), .A2(new_n863), .A3(new_n424), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(KEYINPUT106), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT108), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT106), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n862), .A2(new_n867), .A3(new_n863), .A4(new_n424), .ZN(new_n868));
  AND3_X1   g0668(.A1(new_n865), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n866), .B1(new_n865), .B2(new_n868), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n860), .B1(new_n401), .B2(new_n399), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n420), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n872), .A2(new_n863), .ZN(new_n873));
  NOR3_X1   g0673(.A1(new_n869), .A2(new_n870), .A3(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n667), .ZN(new_n875));
  AND3_X1   g0675(.A1(new_n427), .A2(new_n402), .A3(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n859), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT39), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n384), .A2(new_n386), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n397), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n880), .A2(new_n277), .A3(new_n387), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n860), .B1(new_n881), .B2(new_n401), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT37), .B1(new_n882), .B2(new_n420), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n867), .B1(new_n872), .B2(new_n863), .ZN(new_n884));
  INV_X1    g0684(.A(new_n868), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n881), .A2(new_n401), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n427), .A2(new_n875), .A3(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n886), .A2(KEYINPUT38), .A3(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n877), .A2(new_n878), .A3(new_n889), .ZN(new_n890));
  AND3_X1   g0690(.A1(new_n886), .A2(KEYINPUT38), .A3(new_n888), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT38), .B1(new_n886), .B2(new_n888), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT39), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT107), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n886), .A2(new_n888), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n859), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n889), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n898), .A2(KEYINPUT107), .A3(KEYINPUT39), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n890), .A2(new_n895), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n317), .A2(new_n672), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n438), .A2(new_n667), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n821), .B1(new_n739), .B2(new_n856), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n281), .A2(new_n669), .ZN(new_n907));
  AND3_X1   g0707(.A1(new_n444), .A2(new_n321), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n907), .B1(new_n444), .B2(new_n321), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n906), .A2(new_n898), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n903), .A2(new_n904), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n740), .B1(new_n436), .B2(new_n447), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n658), .B1(new_n738), .B2(new_n914), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n913), .B(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT40), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n714), .A2(new_n718), .ZN(new_n918));
  OAI211_X1 g0718(.A(KEYINPUT31), .B(new_n669), .C1(new_n703), .C2(new_n713), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n697), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT109), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n697), .A2(new_n918), .A3(KEYINPUT109), .A4(new_n919), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n856), .B1(new_n908), .B2(new_n909), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n924), .A2(new_n898), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n917), .B1(new_n877), .B2(new_n889), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n925), .B1(new_n922), .B2(new_n923), .ZN(new_n929));
  AOI22_X1  g0729(.A1(new_n917), .A2(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n448), .A2(new_n924), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n930), .B(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n679), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n916), .B(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n255), .B2(new_n808), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n607), .A2(new_n609), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT35), .ZN(new_n937));
  AOI211_X1 g0737(.A(new_n235), .B(new_n232), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n938), .B(G116), .C1(new_n937), .C2(new_n936), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT36), .ZN(new_n940));
  OAI21_X1  g0740(.A(G77), .B1(new_n217), .B2(new_n210), .ZN(new_n941));
  OAI22_X1  g0741(.A1(new_n234), .A2(new_n941), .B1(G50), .B2(new_n210), .ZN(new_n942));
  INV_X1    g0742(.A(G13), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n942), .A2(G1), .A3(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT105), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n935), .A2(new_n940), .A3(new_n945), .ZN(G367));
  NOR2_X1   g0746(.A1(new_n619), .A2(new_n672), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT110), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n619), .B(new_n624), .C1(new_n621), .C2(new_n672), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  OR3_X1    g0751(.A1(new_n685), .A2(new_n951), .A3(KEYINPUT42), .ZN(new_n952));
  OAI21_X1  g0752(.A(KEYINPUT42), .B1(new_n685), .B2(new_n951), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n646), .B1(new_n950), .B2(new_n662), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n952), .B(new_n953), .C1(new_n669), .C2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n681), .A2(new_n950), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n634), .A2(new_n640), .B1(new_n539), .B2(new_n669), .ZN(new_n957));
  NOR3_X1   g0757(.A1(new_n635), .A2(new_n540), .A3(new_n672), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(KEYINPUT43), .ZN(new_n961));
  AND3_X1   g0761(.A1(new_n955), .A2(new_n956), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n956), .B1(new_n955), .B2(new_n961), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n960), .A2(KEYINPUT43), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  OR3_X1    g0765(.A1(new_n962), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n965), .B1(new_n962), .B2(new_n963), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n691), .B(KEYINPUT41), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n685), .A2(new_n687), .A3(new_n950), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT45), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n685), .A2(KEYINPUT45), .A3(new_n687), .A4(new_n950), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(KEYINPUT44), .B1(new_n688), .B2(new_n950), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n685), .A2(new_n687), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT44), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n976), .A2(new_n977), .A3(new_n951), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n974), .A2(new_n975), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n681), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n674), .A2(new_n680), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n682), .A2(new_n981), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(new_n684), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n974), .A2(new_n975), .A3(new_n682), .A4(new_n978), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n980), .A2(new_n983), .A3(new_n742), .A4(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n969), .B1(new_n985), .B2(new_n742), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n966), .B(new_n967), .C1(new_n986), .C2(new_n810), .ZN(new_n987));
  INV_X1    g0787(.A(new_n800), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n797), .B1(new_n227), .B2(new_n354), .C1(new_n988), .C2(new_n244), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n768), .A2(G116), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n990), .B(KEYINPUT46), .Z(new_n991));
  NOR2_X1   g0791(.A1(new_n756), .A2(new_n219), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(G294), .B2(new_n759), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n774), .A2(G317), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n785), .A2(G311), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n799), .B1(new_n788), .B2(G283), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n993), .A2(new_n994), .A3(new_n995), .A4(new_n996), .ZN(new_n997));
  AOI211_X1 g0797(.A(new_n991), .B(new_n997), .C1(G303), .C2(new_n772), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n763), .A2(G107), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n756), .A2(new_n272), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(G143), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n295), .B1(new_n767), .B2(new_n1002), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n339), .A2(new_n771), .B1(new_n758), .B2(new_n776), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n1003), .B(new_n1004), .C1(new_n774), .C2(G137), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n1005), .B1(new_n222), .B2(new_n747), .C1(new_n210), .C2(new_n764), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1006), .B1(G58), .B2(new_n768), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n998), .A2(new_n999), .B1(new_n1001), .B2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT47), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n811), .B(new_n989), .C1(new_n1009), .C2(new_n745), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(new_n796), .B2(new_n959), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT111), .Z(new_n1012));
  NAND2_X1  g0812(.A1(new_n987), .A2(new_n1012), .ZN(G387));
  OR2_X1    g0813(.A1(new_n983), .A2(new_n742), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n983), .A2(new_n742), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1014), .A2(new_n691), .A3(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n769), .A2(new_n272), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n799), .B1(new_n341), .B2(new_n758), .C1(new_n775), .C2(new_n339), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n1017), .B(new_n1018), .C1(G50), .C2(new_n772), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n992), .B1(G68), .B2(new_n788), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n354), .A2(new_n764), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(G159), .B2(new_n785), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1019), .A2(new_n1020), .A3(new_n1022), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(G311), .A2(new_n759), .B1(new_n772), .B2(G317), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1024), .B1(new_n791), .B2(new_n747), .C1(new_n781), .C2(new_n767), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT48), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1026), .B1(new_n832), .B2(new_n764), .C1(new_n478), .C2(new_n769), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT49), .Z(new_n1028));
  NAND2_X1  g0828(.A1(new_n774), .A2(new_n786), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1029), .B(new_n798), .C1(new_n207), .C2(new_n756), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1023), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n744), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n811), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(new_n674), .B2(new_n796), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n241), .A2(G45), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT112), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n341), .A2(G50), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT50), .ZN(new_n1039));
  AOI21_X1  g0839(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1039), .A2(new_n693), .A3(new_n1040), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1037), .A2(new_n800), .A3(new_n1041), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(G107), .B2(new_n227), .C1(new_n693), .C2(new_n805), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT113), .Z(new_n1044));
  AOI21_X1  g0844(.A(new_n1035), .B1(new_n797), .B2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(new_n810), .B2(new_n983), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1016), .A2(new_n1046), .ZN(G393));
  NAND2_X1  g0847(.A1(new_n980), .A2(new_n984), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n692), .B1(new_n1048), .B2(new_n1015), .ZN(new_n1049));
  AND2_X1   g0849(.A1(new_n1049), .A2(new_n985), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n950), .A2(new_n812), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT114), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n758), .A2(new_n222), .B1(new_n769), .B2(new_n210), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n339), .A2(new_n767), .B1(new_n771), .B2(new_n776), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT51), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1055), .B1(new_n212), .B2(new_n756), .C1(new_n1002), .C2(new_n775), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n1053), .B(new_n1056), .C1(G77), .C2(new_n763), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1057), .B(new_n799), .C1(new_n341), .C2(new_n747), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n775), .A2(new_n781), .B1(new_n832), .B2(new_n769), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT116), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n392), .B1(new_n791), .B2(new_n758), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(G116), .B2(new_n763), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n747), .A2(new_n478), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n1063), .B(new_n757), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(G311), .A2(new_n772), .B1(new_n785), .B2(G317), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT115), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n1066), .B(KEYINPUT52), .Z(new_n1067));
  NAND3_X1  g0867(.A1(new_n1062), .A2(new_n1064), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n745), .B1(new_n1058), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n797), .B1(new_n227), .B2(new_n219), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n800), .B2(new_n252), .ZN(new_n1071));
  OR4_X1    g0871(.A1(new_n1033), .A2(new_n1052), .A3(new_n1069), .A4(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n810), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1072), .B1(new_n1048), .B2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1050), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(G390));
  AOI21_X1  g0876(.A(new_n392), .B1(new_n774), .B2(G125), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n222), .B2(new_n756), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT118), .ZN(new_n1079));
  XOR2_X1   g0879(.A(KEYINPUT54), .B(G143), .Z(new_n1080));
  NAND2_X1  g0880(.A1(new_n788), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n768), .A2(G150), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT53), .Z(new_n1083));
  INV_X1    g0883(.A(G128), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n1084), .A2(new_n767), .B1(new_n771), .B2(new_n846), .ZN(new_n1085));
  INV_X1    g0885(.A(G137), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n758), .A2(new_n1086), .B1(new_n776), .B2(new_n764), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1079), .A2(new_n1081), .A3(new_n1083), .A4(new_n1088), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n758), .A2(new_n205), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n1090), .B(new_n849), .C1(G294), .C2(new_n774), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n763), .A2(G77), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n788), .A2(G97), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n767), .A2(new_n832), .B1(new_n769), .B2(new_n212), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n295), .B(new_n1094), .C1(G116), .C2(new_n772), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .A4(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n745), .B1(new_n1089), .B2(new_n1096), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n1033), .B(new_n1097), .C1(new_n341), .C2(new_n854), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1098), .B1(new_n900), .B2(new_n795), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n901), .B1(new_n905), .B2(new_n910), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n890), .A2(new_n1100), .A3(new_n895), .A4(new_n899), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n902), .B1(new_n877), .B2(new_n889), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n672), .B(new_n820), .C1(new_n725), .C2(new_n728), .ZN(new_n1103));
  AND2_X1   g0903(.A1(new_n1103), .A2(new_n822), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1102), .B1(new_n1104), .B2(new_n910), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n720), .A2(new_n856), .A3(new_n911), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  AND3_X1   g0907(.A1(new_n1101), .A2(new_n1105), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(G330), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n1109), .B(new_n925), .C1(new_n922), .C2(new_n923), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(new_n1101), .B2(new_n1105), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1099), .B1(new_n1112), .B2(new_n1073), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n738), .A2(new_n914), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n448), .A2(G330), .A3(new_n924), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1114), .A2(new_n659), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(KEYINPUT117), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n915), .A2(new_n1118), .A3(new_n1115), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n1109), .B(new_n823), .C1(new_n922), .C2(new_n923), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1104), .B(new_n1106), .C1(new_n1121), .C2(new_n911), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n719), .A2(new_n679), .A3(new_n856), .ZN(new_n1123));
  AND2_X1   g0923(.A1(new_n1123), .A2(new_n910), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n906), .B1(new_n1110), .B2(new_n1124), .ZN(new_n1125));
  AND2_X1   g0925(.A1(new_n1122), .A2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1120), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1101), .A2(new_n1105), .A3(new_n1107), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n1101), .A2(new_n1105), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1128), .B1(new_n1129), .B2(new_n1110), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n692), .B1(new_n1127), .B2(new_n1130), .ZN(new_n1131));
  AND4_X1   g0931(.A1(new_n1118), .A2(new_n1114), .A3(new_n659), .A4(new_n1115), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1118), .B1(new_n915), .B2(new_n1115), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1122), .A2(new_n1125), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n1112), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1113), .B1(new_n1131), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(G378));
  INV_X1    g0939(.A(KEYINPUT57), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n927), .A2(new_n917), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n928), .A2(new_n929), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1141), .A2(new_n1142), .A3(G330), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n347), .A2(new_n875), .ZN(new_n1144));
  XOR2_X1   g0944(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1145));
  XOR2_X1   g0945(.A(new_n1144), .B(new_n1145), .Z(new_n1146));
  AND2_X1   g0946(.A1(new_n653), .A2(new_n654), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1146), .B1(new_n1147), .B2(new_n348), .ZN(new_n1148));
  AND4_X1   g0948(.A1(new_n348), .A2(new_n653), .A3(new_n654), .A4(new_n1146), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1143), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n930), .A2(G330), .A3(new_n1150), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n912), .A2(new_n904), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(new_n902), .B2(new_n900), .ZN(new_n1155));
  AND3_X1   g0955(.A1(new_n1152), .A2(new_n1153), .A3(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1155), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1120), .B1(new_n1130), .B2(new_n1135), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1140), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1150), .B1(new_n930), .B2(G330), .ZN(new_n1161));
  AND4_X1   g0961(.A1(G330), .A2(new_n1141), .A3(new_n1142), .A4(new_n1150), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n913), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1152), .A2(new_n1153), .A3(new_n1155), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1163), .A2(KEYINPUT124), .A3(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT124), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1157), .A2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1134), .B1(new_n1112), .B2(new_n1126), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1165), .A2(KEYINPUT57), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1160), .A2(new_n1169), .A3(new_n691), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n284), .A2(new_n285), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT119), .ZN(new_n1172));
  AOI211_X1 g0972(.A(G50), .B(new_n1172), .C1(new_n798), .C2(new_n285), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n755), .A2(G58), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n772), .A2(G107), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n759), .A2(G97), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1177), .A2(new_n1017), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n285), .B(new_n798), .C1(new_n354), .C2(new_n747), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n767), .A2(new_n207), .B1(new_n210), .B2(new_n764), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1178), .B(new_n1181), .C1(new_n832), .C2(new_n775), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT120), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1173), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT122), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1185), .B(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n774), .A2(G124), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1188), .B(new_n1172), .C1(new_n776), .C2(new_n756), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n758), .A2(new_n846), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1080), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n769), .A2(new_n1191), .B1(new_n339), .B2(new_n764), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1190), .B(new_n1192), .C1(G125), .C2(new_n785), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n1193), .B1(new_n1084), .B2(new_n771), .C1(new_n1086), .C2(new_n747), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1194), .B(KEYINPUT59), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1187), .B1(new_n1183), .B2(new_n1184), .C1(new_n1189), .C2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1196), .A2(new_n744), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1033), .B1(new_n222), .B2(new_n854), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1197), .B(new_n1198), .C1(new_n795), .C2(new_n1150), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT123), .ZN(new_n1200));
  AND2_X1   g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n1158), .A2(new_n1073), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1170), .A2(new_n1204), .ZN(G375));
  NAND2_X1  g1005(.A1(new_n910), .A2(new_n794), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n855), .A2(G68), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n392), .B1(new_n219), .B2(new_n769), .C1(new_n354), .C2(new_n764), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1001), .B1(new_n205), .B2(new_n747), .C1(new_n791), .C2(new_n775), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n1208), .B(new_n1209), .C1(G294), .C2(new_n785), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1210), .B1(new_n207), .B2(new_n758), .C1(new_n832), .C2(new_n771), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1174), .B1(new_n222), .B2(new_n764), .C1(new_n758), .C2(new_n1191), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(G128), .B2(new_n774), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n768), .A2(G159), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n788), .A2(G150), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n798), .B1(new_n772), .B2(G137), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n767), .A2(new_n846), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1211), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n1033), .B(new_n1207), .C1(new_n1219), .C2(new_n744), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n1135), .A2(new_n810), .B1(new_n1206), .B2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1126), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(new_n968), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1221), .B1(new_n1223), .B2(new_n1127), .ZN(G381));
  NOR2_X1   g1024(.A1(G375), .A2(G378), .ZN(new_n1225));
  INV_X1    g1025(.A(G384), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1075), .A2(new_n987), .A3(new_n1012), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(G393), .A2(G396), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  NOR3_X1   g1031(.A1(new_n1227), .A2(G381), .A3(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT125), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NOR4_X1   g1034(.A1(new_n1227), .A2(KEYINPUT125), .A3(G381), .A4(new_n1231), .ZN(new_n1235));
  OR2_X1    g1035(.A1(new_n1234), .A2(new_n1235), .ZN(G407));
  NAND2_X1  g1036(.A1(new_n1225), .A2(new_n668), .ZN(new_n1237));
  OAI211_X1 g1037(.A(G213), .B(new_n1237), .C1(new_n1234), .C2(new_n1235), .ZN(G409));
  INV_X1    g1038(.A(G213), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1239), .A2(G343), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1242), .A2(new_n1168), .A3(new_n968), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1165), .A2(new_n810), .A3(new_n1167), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1138), .A2(new_n1199), .A3(new_n1243), .A4(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1242), .A2(new_n1168), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n692), .B1(new_n1246), .B2(new_n1140), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1203), .B1(new_n1247), .B2(new_n1169), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1241), .B(new_n1245), .C1(new_n1248), .C2(new_n1138), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1135), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT126), .ZN(new_n1251));
  OAI21_X1  g1051(.A(KEYINPUT60), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT60), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1222), .A2(KEYINPUT126), .A3(new_n1253), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1252), .A2(new_n1254), .A3(new_n691), .A4(new_n1136), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n1255), .A2(G384), .A3(new_n1221), .ZN(new_n1256));
  AOI21_X1  g1056(.A(G384), .B1(new_n1255), .B2(new_n1221), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  OAI21_X1  g1059(.A(KEYINPUT62), .B1(new_n1249), .B2(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1240), .B1(G375), .B2(G378), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT62), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1261), .A2(new_n1262), .A3(new_n1258), .A4(new_n1245), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1255), .A2(new_n1221), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(new_n1226), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1255), .A2(G384), .A3(new_n1221), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1240), .A2(G2897), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1265), .A2(new_n1266), .A3(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1267), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1269), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1249), .A2(new_n1268), .A3(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT61), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1260), .A2(new_n1263), .A3(new_n1271), .A4(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(G390), .A2(G387), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n1228), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n816), .B1(new_n1016), .B2(new_n1046), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1230), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1275), .A2(new_n1277), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1274), .B(new_n1228), .C1(new_n1230), .C2(new_n1276), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1273), .A2(new_n1280), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1280), .A2(KEYINPUT61), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT63), .ZN(new_n1283));
  AND2_X1   g1083(.A1(new_n1270), .A2(new_n1268), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1283), .B1(new_n1284), .B2(new_n1249), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1249), .A2(new_n1259), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1282), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1286), .A2(KEYINPUT127), .A3(KEYINPUT63), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1261), .A2(KEYINPUT63), .A3(new_n1258), .A4(new_n1245), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT127), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1288), .A2(new_n1291), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1281), .B1(new_n1287), .B2(new_n1292), .ZN(G405));
  NAND2_X1  g1093(.A1(new_n1248), .A2(new_n1138), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(G375), .A2(G378), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1280), .A2(new_n1294), .A3(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1294), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1297), .A2(new_n1278), .A3(new_n1279), .ZN(new_n1298));
  AND3_X1   g1098(.A1(new_n1296), .A2(new_n1258), .A3(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1258), .B1(new_n1296), .B2(new_n1298), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1299), .A2(new_n1300), .ZN(G402));
endmodule


