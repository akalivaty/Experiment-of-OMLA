//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 1 0 1 1 0 1 0 1 0 1 0 0 1 1 0 1 1 0 1 0 0 1 0 0 0 0 1 1 0 0 0 0 0 1 1 0 0 1 1 1 1 1 0 1 0 1 0 1 0 0 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n797, new_n798, new_n800,
    new_n801, new_n803, new_n804, new_n805, new_n806, new_n807, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202));
  XOR2_X1   g001(.A(new_n202), .B(KEYINPUT13), .Z(new_n203));
  INV_X1    g002(.A(KEYINPUT91), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n204), .A2(G8gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(G15gat), .B(G22gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT90), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G1gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT16), .ZN(new_n210));
  AOI22_X1  g009(.A1(new_n208), .A2(new_n209), .B1(new_n210), .B2(new_n206), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n206), .A2(new_n207), .A3(G1gat), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n205), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n204), .A2(G8gat), .ZN(new_n214));
  OR2_X1    g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n214), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G29gat), .ZN(new_n218));
  INV_X1    g017(.A(G36gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT14), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT14), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(G29gat), .B2(G36gat), .ZN(new_n222));
  OAI211_X1 g021(.A(new_n220), .B(new_n222), .C1(new_n218), .C2(new_n219), .ZN(new_n223));
  INV_X1    g022(.A(G50gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(G43gat), .ZN(new_n225));
  INV_X1    g024(.A(G43gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(G50gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT89), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT15), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  OR3_X1    g029(.A1(new_n223), .A2(new_n228), .A3(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n228), .B1(new_n223), .B2(new_n230), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT15), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n223), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n231), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n217), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT92), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n235), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n215), .A2(new_n239), .A3(new_n216), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n236), .A2(new_n237), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n203), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n235), .A2(KEYINPUT17), .ZN(new_n244));
  OR2_X1    g043(.A1(new_n235), .A2(KEYINPUT17), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n217), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n246), .A2(new_n202), .A3(new_n240), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT18), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  AND2_X1   g048(.A1(new_n246), .A2(new_n240), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n250), .A2(KEYINPUT18), .A3(new_n202), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n243), .A2(new_n249), .A3(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(G113gat), .B(G141gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(KEYINPUT11), .ZN(new_n254));
  INV_X1    g053(.A(G169gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n256), .B(G197gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n257), .B(KEYINPUT12), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n252), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n243), .A2(new_n251), .A3(new_n258), .A4(new_n249), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(G228gat), .A2(G233gat), .ZN(new_n264));
  XOR2_X1   g063(.A(KEYINPUT76), .B(KEYINPUT3), .Z(new_n265));
  OR2_X1    g064(.A1(KEYINPUT70), .A2(KEYINPUT22), .ZN(new_n266));
  NAND2_X1  g065(.A1(G211gat), .A2(G218gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(KEYINPUT70), .A2(KEYINPUT22), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G197gat), .B(G204gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(G211gat), .B(G218gat), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n269), .A2(new_n272), .A3(new_n270), .ZN(new_n275));
  AND3_X1   g074(.A1(new_n274), .A2(KEYINPUT80), .A3(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT29), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n277), .B1(new_n275), .B2(KEYINPUT80), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n265), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  OR2_X1    g078(.A1(G155gat), .A2(G162gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(G155gat), .A2(G162gat), .ZN(new_n281));
  AND2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G141gat), .B(G148gat), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n282), .B(KEYINPUT72), .C1(KEYINPUT2), .C2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT72), .ZN(new_n285));
  INV_X1    g084(.A(G148gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(G141gat), .ZN(new_n287));
  INV_X1    g086(.A(G141gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(G148gat), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT2), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n280), .A2(new_n281), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n285), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n284), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n281), .B1(new_n280), .B2(KEYINPUT2), .ZN(new_n294));
  AND2_X1   g093(.A1(KEYINPUT73), .A2(G141gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(KEYINPUT73), .A2(G141gat), .ZN(new_n296));
  NOR3_X1   g095(.A1(new_n295), .A2(new_n296), .A3(new_n286), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT74), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n298), .B1(new_n288), .B2(G148gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n286), .A2(KEYINPUT74), .A3(G141gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  OAI211_X1 g100(.A(KEYINPUT75), .B(new_n294), .C1(new_n297), .C2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT73), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(new_n288), .ZN(new_n305));
  NAND2_X1  g104(.A1(KEYINPUT73), .A2(G141gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n305), .A2(G148gat), .A3(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n307), .A2(new_n299), .A3(new_n300), .ZN(new_n308));
  AOI21_X1  g107(.A(KEYINPUT75), .B1(new_n308), .B2(new_n294), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n293), .B1(new_n303), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n279), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n274), .A2(new_n275), .ZN(new_n312));
  OAI211_X1 g111(.A(new_n293), .B(new_n265), .C1(new_n303), .C2(new_n309), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n312), .B1(new_n313), .B2(new_n277), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT81), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n311), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  AOI211_X1 g115(.A(KEYINPUT81), .B(new_n312), .C1(new_n313), .C2(new_n277), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n264), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT82), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI211_X1 g119(.A(KEYINPUT82), .B(new_n264), .C1(new_n316), .C2(new_n317), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n294), .B1(new_n297), .B2(new_n301), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT75), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI22_X1  g124(.A1(new_n325), .A2(new_n302), .B1(new_n292), .B2(new_n284), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT3), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n312), .A2(new_n277), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n264), .B1(new_n329), .B2(KEYINPUT83), .ZN(new_n330));
  INV_X1    g129(.A(new_n314), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n310), .A2(KEYINPUT3), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT83), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n332), .B(new_n333), .C1(new_n326), .C2(new_n328), .ZN(new_n334));
  AND3_X1   g133(.A1(new_n330), .A2(new_n331), .A3(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n322), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(G22gat), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n335), .B1(new_n320), .B2(new_n321), .ZN(new_n339));
  INV_X1    g138(.A(G22gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(G78gat), .B(G106gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n342), .B(new_n224), .ZN(new_n343));
  XNOR2_X1  g142(.A(KEYINPUT79), .B(KEYINPUT31), .ZN(new_n344));
  XOR2_X1   g143(.A(new_n343), .B(new_n344), .Z(new_n345));
  NAND4_X1  g144(.A1(new_n338), .A2(KEYINPUT84), .A3(new_n341), .A4(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT84), .B1(new_n339), .B2(new_n340), .ZN(new_n347));
  INV_X1    g146(.A(new_n345), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n340), .B1(new_n322), .B2(new_n336), .ZN(new_n349));
  AOI211_X1 g148(.A(G22gat), .B(new_n335), .C1(new_n320), .C2(new_n321), .ZN(new_n350));
  OAI22_X1  g149(.A1(new_n347), .A2(new_n348), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n312), .ZN(new_n352));
  NAND2_X1  g151(.A1(G226gat), .A2(G233gat), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT24), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n355), .A2(G183gat), .A3(G190gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(G183gat), .B(G190gat), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n356), .B1(new_n357), .B2(new_n355), .ZN(new_n358));
  NOR2_X1   g157(.A1(G169gat), .A2(G176gat), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT25), .B1(new_n359), .B2(KEYINPUT23), .ZN(new_n360));
  NAND2_X1  g159(.A1(G169gat), .A2(G176gat), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT23), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n362), .B1(G169gat), .B2(G176gat), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n360), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n358), .A2(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n366));
  INV_X1    g165(.A(G190gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(KEYINPUT27), .B(G183gat), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(G183gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT27), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT27), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(G183gat), .ZN(new_n373));
  NOR2_X1   g172(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n371), .A2(new_n373), .A3(new_n367), .A4(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(G183gat), .A2(G190gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n369), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(G176gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n255), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT26), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT64), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n359), .A2(KEYINPUT64), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n361), .B(new_n381), .C1(new_n385), .C2(KEYINPUT26), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n365), .B1(new_n378), .B2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT65), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n388), .B(new_n356), .C1(new_n357), .C2(new_n355), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n383), .A2(KEYINPUT23), .A3(new_n384), .ZN(new_n390));
  AND2_X1   g189(.A1(new_n363), .A2(new_n361), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n367), .A2(G183gat), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n370), .A2(G190gat), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT24), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n388), .B1(new_n395), .B2(new_n356), .ZN(new_n396));
  OAI21_X1  g195(.A(KEYINPUT25), .B1(new_n392), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n387), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n354), .B1(new_n398), .B2(new_n277), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n353), .B1(new_n387), .B2(new_n397), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n352), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n398), .A2(new_n354), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT29), .B1(new_n387), .B2(new_n397), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n402), .B(new_n312), .C1(new_n354), .C2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(G64gat), .B(G92gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n406), .B(KEYINPUT71), .ZN(new_n407));
  XNOR2_X1  g206(.A(G8gat), .B(G36gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n407), .B(new_n408), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT30), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n405), .A2(new_n409), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT30), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n413), .B1(new_n405), .B2(new_n409), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n411), .A2(new_n412), .A3(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(G134gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(G113gat), .B(G120gat), .ZN(new_n418));
  NOR2_X1   g217(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  NOR3_X1   g219(.A1(new_n418), .A2(G127gat), .A3(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(G127gat), .ZN(new_n422));
  INV_X1    g221(.A(G120gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(G113gat), .ZN(new_n424));
  INV_X1    g223(.A(G113gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(G120gat), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n422), .B1(new_n427), .B2(new_n419), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n417), .B1(new_n421), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(G127gat), .B1(new_n418), .B2(new_n420), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n427), .A2(new_n422), .A3(new_n419), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n430), .A2(new_n431), .A3(G134gat), .ZN(new_n432));
  AND3_X1   g231(.A1(new_n429), .A2(KEYINPUT68), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(KEYINPUT68), .B1(new_n429), .B2(new_n432), .ZN(new_n434));
  OR3_X1    g233(.A1(new_n398), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n398), .B1(new_n433), .B2(new_n434), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(G227gat), .ZN(new_n438));
  INV_X1    g237(.A(G233gat), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n437), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT34), .ZN(new_n443));
  XNOR2_X1  g242(.A(KEYINPUT69), .B(G71gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n444), .B(G99gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(G15gat), .B(G43gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n445), .B(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n435), .A2(new_n440), .A3(new_n436), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT33), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n448), .A2(KEYINPUT32), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT34), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n437), .A2(new_n453), .A3(new_n441), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n448), .B(KEYINPUT32), .C1(new_n449), .C2(new_n447), .ZN(new_n455));
  AND4_X1   g254(.A1(new_n443), .A2(new_n452), .A3(new_n454), .A4(new_n455), .ZN(new_n456));
  AOI22_X1  g255(.A1(new_n452), .A2(new_n455), .B1(new_n443), .B2(new_n454), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AND4_X1   g257(.A1(new_n346), .A2(new_n351), .A3(new_n416), .A4(new_n458), .ZN(new_n459));
  OAI211_X1 g258(.A(KEYINPUT4), .B(new_n326), .C1(new_n433), .C2(new_n434), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n429), .A2(new_n432), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n313), .B(new_n461), .C1(new_n326), .C2(new_n327), .ZN(new_n462));
  NAND2_X1  g261(.A1(G225gat), .A2(G233gat), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT4), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n464), .B1(new_n310), .B2(new_n461), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n460), .A2(new_n462), .A3(new_n463), .A4(new_n465), .ZN(new_n466));
  XNOR2_X1  g265(.A(KEYINPUT77), .B(KEYINPUT5), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n310), .A2(new_n461), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n430), .A2(new_n431), .A3(G134gat), .ZN(new_n469));
  AOI21_X1  g268(.A(G134gat), .B1(new_n430), .B2(new_n431), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n326), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n463), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n467), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n466), .A2(new_n475), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n464), .B(new_n326), .C1(new_n433), .C2(new_n434), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n472), .A2(KEYINPUT4), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n471), .B1(new_n310), .B2(KEYINPUT3), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n474), .B1(new_n480), .B2(new_n313), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n479), .A2(new_n481), .A3(new_n467), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n476), .A2(new_n482), .ZN(new_n483));
  XOR2_X1   g282(.A(G57gat), .B(G85gat), .Z(new_n484));
  XNOR2_X1  g283(.A(G1gat), .B(G29gat), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n484), .B(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n486), .B(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n483), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT6), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n476), .A2(new_n488), .A3(new_n482), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  AOI211_X1 g292(.A(new_n491), .B(new_n488), .C1(new_n476), .C2(new_n482), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT35), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AND3_X1   g298(.A1(new_n462), .A2(new_n463), .A3(new_n467), .ZN(new_n500));
  AOI22_X1  g299(.A1(new_n466), .A2(new_n475), .B1(new_n500), .B2(new_n479), .ZN(new_n501));
  XOR2_X1   g300(.A(new_n488), .B(KEYINPUT85), .Z(new_n502));
  OAI211_X1 g301(.A(new_n492), .B(new_n491), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT86), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n494), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OR2_X1    g304(.A1(new_n501), .A2(new_n502), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n506), .A2(KEYINPUT86), .A3(new_n491), .A4(new_n492), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n415), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n508), .A2(new_n351), .A3(new_n346), .A4(new_n458), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n459), .A2(new_n499), .B1(new_n509), .B2(new_n498), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT37), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n401), .A2(new_n511), .A3(new_n404), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(new_n409), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n511), .B1(new_n401), .B2(new_n404), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT38), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT88), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI211_X1 g316(.A(KEYINPUT88), .B(KEYINPUT38), .C1(new_n513), .C2(new_n514), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(KEYINPUT87), .B1(new_n405), .B2(KEYINPUT37), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT87), .ZN(new_n521));
  AOI211_X1 g320(.A(new_n521), .B(new_n511), .C1(new_n401), .C2(new_n404), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n513), .A2(KEYINPUT38), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n410), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n519), .A2(new_n507), .A3(new_n505), .A4(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n479), .A2(new_n462), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(new_n474), .ZN(new_n528));
  OR2_X1    g327(.A1(new_n528), .A2(KEYINPUT39), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n468), .A2(new_n472), .A3(new_n463), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n528), .A2(KEYINPUT39), .A3(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n529), .A2(new_n502), .A3(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT40), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n529), .A2(KEYINPUT40), .A3(new_n531), .A4(new_n502), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n534), .A2(new_n415), .A3(new_n506), .A4(new_n535), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n526), .A2(new_n346), .A3(new_n351), .A4(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n351), .A2(new_n346), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n416), .A2(new_n496), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n458), .A2(KEYINPUT36), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT36), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n542), .B1(new_n456), .B2(new_n457), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n537), .A2(new_n540), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n263), .B1(new_n510), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT21), .ZN(new_n547));
  XNOR2_X1  g346(.A(G71gat), .B(G78gat), .ZN(new_n548));
  OR2_X1    g347(.A1(new_n548), .A2(KEYINPUT95), .ZN(new_n549));
  INV_X1    g348(.A(G64gat), .ZN(new_n550));
  INV_X1    g349(.A(G57gat), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n550), .B1(new_n551), .B2(KEYINPUT94), .ZN(new_n552));
  NAND2_X1  g351(.A1(G57gat), .A2(G64gat), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n553), .A2(KEYINPUT94), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT9), .ZN(new_n555));
  NAND2_X1  g354(.A1(G71gat), .A2(G78gat), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n548), .A2(KEYINPUT95), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n549), .A2(new_n552), .A3(new_n557), .A4(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT93), .ZN(new_n560));
  OR2_X1    g359(.A1(new_n548), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n556), .A2(new_n555), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n551), .A2(new_n550), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n562), .A2(new_n553), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n560), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n561), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n559), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n217), .B1(new_n547), .B2(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(G183gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n547), .ZN(new_n570));
  NAND2_X1  g369(.A1(G231gat), .A2(G233gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(G127gat), .B(G155gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(KEYINPUT96), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n572), .B(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n569), .B(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(G211gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n576), .B(new_n578), .ZN(new_n579));
  AND2_X1   g378(.A1(G232gat), .A2(G233gat), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n580), .A2(KEYINPUT41), .ZN(new_n581));
  XNOR2_X1  g380(.A(G134gat), .B(G162gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G190gat), .B(G218gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT100), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  AOI22_X1  g386(.A1(new_n587), .A2(KEYINPUT101), .B1(KEYINPUT41), .B2(new_n580), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  XOR2_X1   g388(.A(KEYINPUT97), .B(G92gat), .Z(new_n590));
  INV_X1    g389(.A(G85gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(G99gat), .A2(G106gat), .ZN(new_n592));
  AOI22_X1  g391(.A1(new_n590), .A2(new_n591), .B1(KEYINPUT8), .B2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT98), .ZN(new_n594));
  XOR2_X1   g393(.A(G99gat), .B(G106gat), .Z(new_n595));
  NAND2_X1  g394(.A1(G85gat), .A2(G92gat), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n596), .A2(KEYINPUT7), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(KEYINPUT7), .ZN(new_n598));
  AOI22_X1  g397(.A1(new_n595), .A2(KEYINPUT99), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n594), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n595), .A2(KEYINPUT99), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI211_X1 g401(.A(new_n594), .B(new_n599), .C1(KEYINPUT99), .C2(new_n595), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n589), .B1(new_n604), .B2(new_n239), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n587), .A2(KEYINPUT101), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n602), .A2(new_n244), .A3(new_n603), .A4(new_n245), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n605), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n607), .B1(new_n605), .B2(new_n608), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n584), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n611), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n613), .A2(new_n583), .A3(new_n609), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n579), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n567), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n604), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT10), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n602), .A2(new_n567), .A3(new_n603), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n604), .A2(KEYINPUT10), .A3(new_n618), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(G230gat), .A2(G233gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n619), .A2(new_n621), .ZN(new_n627));
  INV_X1    g426(.A(new_n625), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(G120gat), .B(G148gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(G176gat), .ZN(new_n632));
  INV_X1    g431(.A(G204gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n630), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n626), .A2(new_n629), .A3(new_n634), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  AND3_X1   g438(.A1(new_n546), .A2(new_n617), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(new_n497), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n415), .ZN(new_n643));
  XNOR2_X1  g442(.A(KEYINPUT16), .B(G8gat), .ZN(new_n644));
  OR2_X1    g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT42), .ZN(new_n646));
  OR2_X1    g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n643), .A2(G8gat), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n645), .A2(new_n646), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(G1325gat));
  AOI21_X1  g449(.A(G15gat), .B1(new_n640), .B2(new_n458), .ZN(new_n651));
  INV_X1    g450(.A(new_n544), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(G15gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT102), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n651), .B1(new_n640), .B2(new_n654), .ZN(G1326gat));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n538), .ZN(new_n656));
  XNOR2_X1  g455(.A(KEYINPUT43), .B(G22gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(G1327gat));
  OR2_X1    g457(.A1(new_n639), .A2(KEYINPUT103), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n639), .A2(KEYINPUT103), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NOR3_X1   g460(.A1(new_n661), .A2(new_n263), .A3(new_n579), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n509), .A2(new_n498), .ZN(new_n664));
  AND2_X1   g463(.A1(new_n351), .A2(new_n346), .ZN(new_n665));
  NAND4_X1  g464(.A1(new_n665), .A2(new_n416), .A3(new_n458), .A4(new_n499), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n545), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n615), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(KEYINPUT44), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n615), .B1(new_n510), .B2(new_n545), .ZN(new_n671));
  XOR2_X1   g470(.A(KEYINPUT104), .B(KEYINPUT44), .Z(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n663), .B1(new_n670), .B2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(G29gat), .B1(new_n675), .B2(new_n496), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n579), .A2(new_n615), .A3(new_n638), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n546), .A2(new_n218), .A3(new_n497), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT45), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n676), .A2(new_n679), .ZN(G1328gat));
  OAI21_X1  g479(.A(G36gat), .B1(new_n675), .B2(new_n416), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n546), .A2(new_n219), .A3(new_n415), .A4(new_n677), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n682), .B(KEYINPUT46), .Z(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(G1329gat));
  NAND4_X1  g483(.A1(new_n546), .A2(new_n226), .A3(new_n458), .A4(new_n677), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n674), .A2(new_n652), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n685), .B1(new_n687), .B2(new_n226), .ZN(new_n688));
  XNOR2_X1  g487(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  OAI211_X1 g490(.A(new_n689), .B(new_n685), .C1(new_n687), .C2(new_n226), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(G1330gat));
  INV_X1    g492(.A(new_n672), .ZN(new_n694));
  AOI211_X1 g493(.A(new_n615), .B(new_n694), .C1(new_n510), .C2(new_n545), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n696), .B1(new_n667), .B2(new_n668), .ZN(new_n697));
  OAI211_X1 g496(.A(new_n538), .B(new_n662), .C1(new_n695), .C2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(G50gat), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n546), .A2(new_n224), .A3(new_n538), .A4(new_n677), .ZN(new_n700));
  AOI22_X1  g499(.A1(new_n699), .A2(new_n700), .B1(KEYINPUT106), .B2(KEYINPUT48), .ZN(new_n701));
  NOR2_X1   g500(.A1(KEYINPUT106), .A2(KEYINPUT48), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(G1331gat));
  AND4_X1   g502(.A1(new_n667), .A2(new_n263), .A3(new_n617), .A4(new_n661), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(new_n497), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g505(.A1(new_n704), .A2(new_n415), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n707), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n708));
  XOR2_X1   g507(.A(KEYINPUT49), .B(G64gat), .Z(new_n709));
  OAI21_X1  g508(.A(new_n708), .B1(new_n707), .B2(new_n709), .ZN(G1333gat));
  NAND2_X1  g509(.A1(new_n704), .A2(new_n652), .ZN(new_n711));
  INV_X1    g510(.A(new_n458), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n712), .A2(G71gat), .ZN(new_n713));
  AOI22_X1  g512(.A1(new_n711), .A2(G71gat), .B1(new_n704), .B2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g514(.A1(new_n704), .A2(new_n538), .ZN(new_n716));
  XOR2_X1   g515(.A(KEYINPUT107), .B(G78gat), .Z(new_n717));
  XNOR2_X1  g516(.A(new_n716), .B(new_n717), .ZN(G1335gat));
  NOR2_X1   g517(.A1(new_n579), .A2(new_n262), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n638), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n720), .B1(new_n670), .B2(new_n673), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(G85gat), .B1(new_n722), .B2(new_n496), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT51), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT108), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n719), .B1(new_n671), .B2(new_n725), .ZN(new_n726));
  AOI211_X1 g525(.A(KEYINPUT108), .B(new_n615), .C1(new_n510), .C2(new_n545), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n724), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n669), .A2(KEYINPUT108), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n671), .A2(new_n725), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n729), .A2(KEYINPUT51), .A3(new_n730), .A4(new_n719), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n638), .A2(new_n591), .A3(new_n497), .ZN(new_n733));
  XOR2_X1   g532(.A(new_n733), .B(KEYINPUT109), .Z(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n723), .A2(new_n735), .ZN(G1336gat));
  INV_X1    g535(.A(new_n661), .ZN(new_n737));
  OR3_X1    g536(.A1(new_n737), .A2(G92gat), .A3(new_n416), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n719), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n740), .B1(new_n669), .B2(KEYINPUT108), .ZN(new_n741));
  AOI21_X1  g540(.A(KEYINPUT51), .B1(new_n741), .B2(new_n730), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n726), .A2(new_n724), .A3(new_n727), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n739), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(new_n720), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n415), .B(new_n745), .C1(new_n695), .C2(new_n697), .ZN(new_n746));
  INV_X1    g545(.A(new_n590), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT110), .ZN(new_n749));
  OAI211_X1 g548(.A(new_n744), .B(new_n748), .C1(new_n749), .C2(KEYINPUT52), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n749), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT52), .ZN(new_n752));
  INV_X1    g551(.A(new_n748), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n738), .B1(new_n728), .B2(new_n731), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n751), .B(new_n752), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  AND2_X1   g554(.A1(new_n750), .A2(new_n755), .ZN(G1337gat));
  OAI21_X1  g555(.A(G99gat), .B1(new_n722), .B2(new_n544), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n712), .A2(new_n639), .A3(G99gat), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n732), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n757), .A2(new_n759), .ZN(G1338gat));
  INV_X1    g559(.A(G106gat), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n661), .A2(new_n761), .A3(new_n538), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n762), .B1(new_n728), .B2(new_n731), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n761), .B1(new_n721), .B2(new_n538), .ZN(new_n764));
  OR3_X1    g563(.A1(new_n763), .A2(new_n764), .A3(KEYINPUT53), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT53), .B1(new_n763), .B2(new_n764), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(G1339gat));
  INV_X1    g566(.A(new_n579), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n769));
  AND3_X1   g568(.A1(new_n622), .A2(new_n623), .A3(new_n628), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n628), .B1(new_n622), .B2(new_n623), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT54), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n624), .A2(new_n772), .A3(new_n625), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(new_n635), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n769), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n622), .A2(new_n623), .A3(new_n628), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n626), .A2(KEYINPUT54), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n634), .B1(new_n771), .B2(new_n772), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n778), .A2(KEYINPUT55), .A3(new_n779), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n776), .A2(new_n262), .A3(new_n637), .A4(new_n780), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n241), .A2(new_n203), .A3(new_n242), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n250), .A2(new_n202), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n257), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n638), .A2(new_n261), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n668), .B1(new_n781), .B2(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n776), .A2(new_n637), .A3(new_n780), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n668), .A2(new_n261), .A3(new_n784), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n768), .B1(new_n786), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n617), .A2(new_n263), .A3(new_n639), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n496), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n792), .A2(new_n459), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n262), .ZN(new_n794));
  XNOR2_X1  g593(.A(KEYINPUT111), .B(G113gat), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n794), .B(new_n795), .ZN(G1340gat));
  AOI21_X1  g595(.A(G120gat), .B1(new_n793), .B2(new_n638), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n737), .A2(new_n423), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n797), .B1(new_n793), .B2(new_n798), .ZN(G1341gat));
  NAND2_X1  g598(.A1(new_n793), .A2(new_n579), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n422), .A2(KEYINPUT112), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n800), .B(new_n801), .ZN(G1342gat));
  NAND2_X1  g601(.A1(new_n793), .A2(new_n668), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(G134gat), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n793), .A2(new_n417), .A3(new_n668), .ZN(new_n805));
  AND3_X1   g604(.A1(new_n805), .A2(KEYINPUT113), .A3(KEYINPUT56), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT113), .B1(new_n805), .B2(KEYINPUT56), .ZN(new_n807));
  OAI221_X1 g606(.A(new_n804), .B1(KEYINPUT56), .B2(new_n805), .C1(new_n806), .C2(new_n807), .ZN(G1343gat));
  INV_X1    g607(.A(new_n792), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n544), .A2(new_n538), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n810), .A2(KEYINPUT115), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n810), .A2(KEYINPUT115), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n416), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n262), .A2(new_n288), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n814), .B(KEYINPUT116), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n809), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n652), .A2(new_n496), .A3(new_n415), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n665), .B1(new_n790), .B2(new_n791), .ZN(new_n819));
  XOR2_X1   g618(.A(KEYINPUT114), .B(KEYINPUT57), .Z(new_n820));
  OAI21_X1  g619(.A(new_n818), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  AOI211_X1 g620(.A(KEYINPUT57), .B(new_n665), .C1(new_n790), .C2(new_n791), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n821), .A2(new_n822), .A3(new_n263), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n295), .A2(new_n296), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n817), .B(KEYINPUT118), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT117), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n825), .A2(new_n826), .A3(KEYINPUT58), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n790), .A2(new_n791), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n538), .ZN(new_n829));
  INV_X1    g628(.A(new_n820), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT57), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n819), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n831), .A2(new_n262), .A3(new_n833), .A4(new_n818), .ZN(new_n834));
  INV_X1    g633(.A(new_n824), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n816), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(KEYINPUT117), .B1(new_n836), .B2(KEYINPUT118), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT58), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n838), .B1(new_n836), .B2(KEYINPUT117), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n827), .B1(new_n837), .B2(new_n839), .ZN(G1344gat));
  XOR2_X1   g639(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n841));
  NAND2_X1  g640(.A1(new_n818), .A2(new_n638), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n829), .A2(new_n832), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n819), .A2(new_n830), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n842), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n841), .B1(new_n845), .B2(new_n286), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n831), .A2(new_n638), .A3(new_n833), .A4(new_n818), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n286), .A2(KEYINPUT59), .ZN(new_n848));
  AND3_X1   g647(.A1(new_n847), .A2(KEYINPUT119), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(KEYINPUT119), .B1(new_n847), .B2(new_n848), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n846), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n809), .A2(new_n813), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n852), .A2(new_n286), .A3(new_n638), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(new_n853), .ZN(G1345gat));
  NAND3_X1  g653(.A1(new_n831), .A2(new_n833), .A3(new_n818), .ZN(new_n855));
  OAI21_X1  g654(.A(G155gat), .B1(new_n855), .B2(new_n768), .ZN(new_n856));
  INV_X1    g655(.A(new_n852), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n768), .A2(G155gat), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n856), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT121), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n856), .B(KEYINPUT121), .C1(new_n857), .C2(new_n859), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(G1346gat));
  OAI21_X1  g663(.A(G162gat), .B1(new_n855), .B2(new_n615), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n615), .A2(G162gat), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n865), .B1(new_n857), .B2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT122), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n865), .B(KEYINPUT122), .C1(new_n857), .C2(new_n867), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(G1347gat));
  AOI21_X1  g671(.A(new_n497), .B1(new_n790), .B2(new_n791), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n538), .A2(new_n712), .A3(new_n416), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(G169gat), .B1(new_n875), .B2(new_n263), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n876), .A2(KEYINPUT124), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n876), .A2(KEYINPUT124), .ZN(new_n878));
  INV_X1    g677(.A(new_n875), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(KEYINPUT123), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT123), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n875), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n262), .A2(new_n255), .ZN(new_n884));
  OAI22_X1  g683(.A1(new_n877), .A2(new_n878), .B1(new_n883), .B2(new_n884), .ZN(G1348gat));
  NOR3_X1   g684(.A1(new_n875), .A2(new_n379), .A3(new_n737), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n880), .A2(new_n638), .A3(new_n882), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(new_n379), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(KEYINPUT125), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT125), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n887), .A2(new_n890), .A3(new_n379), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n886), .B1(new_n889), .B2(new_n891), .ZN(G1349gat));
  NAND2_X1  g691(.A1(new_n879), .A2(new_n579), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n893), .A2(new_n368), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT60), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n893), .A2(new_n370), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n895), .B1(new_n894), .B2(new_n896), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n897), .A2(new_n898), .ZN(G1350gat));
  NAND2_X1  g698(.A1(new_n879), .A2(new_n668), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(G190gat), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(KEYINPUT126), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT126), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n900), .A2(new_n903), .A3(G190gat), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n902), .A2(KEYINPUT61), .A3(new_n904), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n880), .A2(new_n367), .A3(new_n668), .A4(new_n882), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n905), .B(new_n906), .C1(KEYINPUT61), .C2(new_n902), .ZN(G1351gat));
  AND4_X1   g706(.A1(new_n538), .A2(new_n873), .A3(new_n415), .A4(new_n544), .ZN(new_n908));
  INV_X1    g707(.A(G197gat), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n908), .A2(new_n909), .A3(new_n262), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT127), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n843), .A2(new_n844), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n652), .A2(new_n497), .A3(new_n416), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n911), .B1(new_n914), .B2(new_n263), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(G197gat), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n914), .A2(new_n911), .A3(new_n263), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n910), .B1(new_n916), .B2(new_n917), .ZN(G1352gat));
  NAND3_X1  g717(.A1(new_n908), .A2(new_n633), .A3(new_n638), .ZN(new_n919));
  XOR2_X1   g718(.A(new_n919), .B(KEYINPUT62), .Z(new_n920));
  OAI21_X1  g719(.A(G204gat), .B1(new_n914), .B2(new_n737), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1353gat));
  INV_X1    g721(.A(G211gat), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n908), .A2(new_n923), .A3(new_n579), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n912), .A2(new_n579), .A3(new_n913), .ZN(new_n925));
  AND3_X1   g724(.A1(new_n925), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n926));
  AOI21_X1  g725(.A(KEYINPUT63), .B1(new_n925), .B2(G211gat), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n924), .B1(new_n926), .B2(new_n927), .ZN(G1354gat));
  AOI21_X1  g727(.A(G218gat), .B1(new_n908), .B2(new_n668), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n912), .A2(new_n913), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n668), .A2(G218gat), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n929), .B1(new_n930), .B2(new_n931), .ZN(G1355gat));
endmodule


