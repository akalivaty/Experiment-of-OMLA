

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754;

  NOR2_X2 U377 ( .A1(n372), .A2(n615), .ZN(n388) );
  XNOR2_X2 U378 ( .A(n618), .B(KEYINPUT82), .ZN(n372) );
  XNOR2_X2 U379 ( .A(n422), .B(KEYINPUT45), .ZN(n655) );
  INV_X1 U380 ( .A(n634), .ZN(n646) );
  NOR2_X1 U381 ( .A1(n542), .A2(n459), .ZN(n634) );
  NAND2_X1 U382 ( .A1(n542), .A2(n459), .ZN(n642) );
  INV_X1 U383 ( .A(n549), .ZN(n576) );
  NOR2_X1 U384 ( .A1(n355), .A2(n356), .ZN(n392) );
  NAND2_X1 U385 ( .A1(n646), .A2(n642), .ZN(n664) );
  INV_X1 U386 ( .A(KEYINPUT32), .ZN(n554) );
  NOR2_X1 U387 ( .A1(n725), .A2(n623), .ZN(n624) );
  NOR2_X1 U388 ( .A1(n725), .A2(n717), .ZN(n718) );
  NOR2_X1 U389 ( .A1(n725), .A2(n704), .ZN(n705) );
  NAND2_X1 U390 ( .A1(n381), .A2(n386), .ZN(n716) );
  NAND2_X1 U391 ( .A1(n393), .A2(n392), .ZN(n391) );
  XNOR2_X1 U392 ( .A(n547), .B(KEYINPUT22), .ZN(n553) );
  OR2_X1 U393 ( .A1(n546), .A2(n545), .ZN(n547) );
  NAND2_X1 U394 ( .A1(n662), .A2(n544), .ZN(n545) );
  XNOR2_X1 U395 ( .A(n581), .B(KEYINPUT1), .ZN(n611) );
  XNOR2_X1 U396 ( .A(n714), .B(n713), .ZN(n715) );
  NAND2_X1 U397 ( .A1(n446), .A2(n445), .ZN(n460) );
  INV_X2 U398 ( .A(G953), .ZN(n514) );
  NAND2_X2 U399 ( .A1(n387), .A2(n365), .ZN(n386) );
  NAND2_X1 U400 ( .A1(n388), .A2(n655), .ZN(n387) );
  AND2_X1 U401 ( .A1(n561), .A2(n364), .ZN(n423) );
  NAND2_X1 U402 ( .A1(n655), .A2(n390), .ZN(n389) );
  NOR2_X1 U403 ( .A1(n410), .A2(n557), .ZN(n407) );
  NOR2_X1 U404 ( .A1(G953), .A2(G237), .ZN(n462) );
  INV_X1 U405 ( .A(KEYINPUT48), .ZN(n395) );
  XNOR2_X1 U406 ( .A(G134), .B(G131), .ZN(n737) );
  XOR2_X1 U407 ( .A(G140), .B(G137), .Z(n521) );
  XNOR2_X1 U408 ( .A(n737), .B(n414), .ZN(n517) );
  INV_X1 U409 ( .A(G146), .ZN(n414) );
  XNOR2_X1 U410 ( .A(n520), .B(n516), .ZN(n415) );
  XNOR2_X1 U411 ( .A(n371), .B(n370), .ZN(n528) );
  INV_X1 U412 ( .A(KEYINPUT95), .ZN(n370) );
  OR2_X1 U413 ( .A1(G237), .A2(G902), .ZN(n502) );
  INV_X1 U414 ( .A(KEYINPUT0), .ZN(n512) );
  XNOR2_X1 U415 ( .A(n379), .B(n357), .ZN(n562) );
  OR2_X1 U416 ( .A1(n620), .A2(G902), .ZN(n379) );
  XNOR2_X1 U417 ( .A(n534), .B(n533), .ZN(n694) );
  XNOR2_X1 U418 ( .A(n532), .B(n531), .ZN(n533) );
  NAND2_X1 U419 ( .A1(n611), .A2(n530), .ZN(n534) );
  INV_X1 U420 ( .A(KEYINPUT72), .ZN(n531) );
  XNOR2_X1 U421 ( .A(n574), .B(n398), .ZN(n397) );
  INV_X1 U422 ( .A(KEYINPUT39), .ZN(n398) );
  NOR2_X1 U423 ( .A1(n596), .A2(n573), .ZN(n574) );
  XNOR2_X1 U424 ( .A(n412), .B(n358), .ZN(n581) );
  OR2_X1 U425 ( .A1(n706), .A2(G902), .ZN(n412) );
  XNOR2_X1 U426 ( .A(n483), .B(KEYINPUT25), .ZN(n484) );
  NOR2_X1 U427 ( .A1(n722), .A2(G902), .ZN(n485) );
  NOR2_X1 U428 ( .A1(G952), .A2(n514), .ZN(n725) );
  INV_X1 U429 ( .A(n389), .ZN(n659) );
  OR2_X1 U430 ( .A1(KEYINPUT2), .A2(n655), .ZN(n656) );
  INV_X1 U431 ( .A(G143), .ZN(n444) );
  NOR2_X1 U432 ( .A1(n609), .A2(n648), .ZN(n377) );
  XOR2_X1 U433 ( .A(KEYINPUT88), .B(G104), .Z(n519) );
  XNOR2_X1 U434 ( .A(G107), .B(G110), .ZN(n518) );
  NAND2_X1 U435 ( .A1(n754), .A2(n407), .ZN(n406) );
  XNOR2_X1 U436 ( .A(G119), .B(G113), .ZN(n466) );
  INV_X1 U437 ( .A(G137), .ZN(n465) );
  XOR2_X1 U438 ( .A(G113), .B(G104), .Z(n494) );
  XNOR2_X1 U439 ( .A(G122), .B(G107), .ZN(n498) );
  XOR2_X1 U440 ( .A(G119), .B(G110), .Z(n495) );
  XOR2_X1 U441 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n448) );
  XNOR2_X1 U442 ( .A(G116), .B(G134), .ZN(n447) );
  XNOR2_X1 U443 ( .A(G143), .B(G122), .ZN(n437) );
  XOR2_X1 U444 ( .A(G140), .B(G131), .Z(n433) );
  XNOR2_X1 U445 ( .A(KEYINPUT89), .B(KEYINPUT84), .ZN(n486) );
  NAND2_X1 U446 ( .A1(G237), .A2(G234), .ZN(n505) );
  NAND2_X1 U447 ( .A1(n394), .A2(n363), .ZN(n618) );
  INV_X1 U448 ( .A(n653), .ZN(n614) );
  INV_X1 U449 ( .A(KEYINPUT38), .ZN(n572) );
  XNOR2_X1 U450 ( .A(n378), .B(n563), .ZN(n568) );
  XNOR2_X1 U451 ( .A(G128), .B(KEYINPUT23), .ZN(n477) );
  XNOR2_X1 U452 ( .A(n415), .B(n413), .ZN(n524) );
  INV_X1 U453 ( .A(n517), .ZN(n413) );
  XNOR2_X1 U454 ( .A(n611), .B(n411), .ZN(n595) );
  INV_X1 U455 ( .A(KEYINPUT86), .ZN(n411) );
  NAND2_X1 U456 ( .A1(n592), .A2(n660), .ZN(n610) );
  XNOR2_X1 U457 ( .A(n504), .B(n503), .ZN(n601) );
  XNOR2_X1 U458 ( .A(n562), .B(n425), .ZN(n529) );
  XNOR2_X1 U459 ( .A(n426), .B(KEYINPUT101), .ZN(n425) );
  INV_X1 U460 ( .A(KEYINPUT6), .ZN(n426) );
  NAND2_X1 U461 ( .A1(n380), .A2(n386), .ZN(n720) );
  AND2_X1 U462 ( .A1(n389), .A2(G217), .ZN(n380) );
  AND2_X1 U463 ( .A1(n389), .A2(G475), .ZN(n381) );
  AND2_X2 U464 ( .A1(n386), .A2(n389), .ZN(n382) );
  AND2_X1 U465 ( .A1(n397), .A2(n639), .ZN(n575) );
  XNOR2_X1 U466 ( .A(n540), .B(KEYINPUT35), .ZN(n749) );
  INV_X1 U467 ( .A(KEYINPUT107), .ZN(n384) );
  NOR2_X1 U468 ( .A1(n596), .A2(n597), .ZN(n385) );
  NAND2_X1 U469 ( .A1(n393), .A2(n403), .ZN(n556) );
  NOR2_X1 U470 ( .A1(n611), .A2(n359), .ZN(n403) );
  OR2_X1 U471 ( .A1(n526), .A2(n367), .ZN(n525) );
  NAND2_X1 U472 ( .A1(n368), .A2(n581), .ZN(n367) );
  INV_X1 U473 ( .A(n555), .ZN(n368) );
  INV_X1 U474 ( .A(KEYINPUT124), .ZN(n416) );
  AND2_X1 U475 ( .A1(n699), .A2(n514), .ZN(n369) );
  XOR2_X1 U476 ( .A(KEYINPUT102), .B(n552), .Z(n355) );
  XNOR2_X1 U477 ( .A(KEYINPUT78), .B(n590), .ZN(n356) );
  XOR2_X1 U478 ( .A(KEYINPUT73), .B(G472), .Z(n357) );
  XOR2_X1 U479 ( .A(KEYINPUT69), .B(G469), .Z(n358) );
  OR2_X1 U480 ( .A1(n555), .A2(n549), .ZN(n359) );
  AND2_X1 U481 ( .A1(n751), .A2(n407), .ZN(n360) );
  AND2_X1 U482 ( .A1(n389), .A2(G472), .ZN(n361) );
  AND2_X1 U483 ( .A1(n389), .A2(G210), .ZN(n362) );
  AND2_X1 U484 ( .A1(n614), .A2(n652), .ZN(n363) );
  AND2_X1 U485 ( .A1(n551), .A2(n626), .ZN(n364) );
  OR2_X1 U486 ( .A1(n617), .A2(n616), .ZN(n365) );
  XNOR2_X1 U487 ( .A(G902), .B(KEYINPUT15), .ZN(n615) );
  XOR2_X1 U488 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n366) );
  INV_X1 U489 ( .A(KEYINPUT65), .ZN(n410) );
  XNOR2_X1 U490 ( .A(n369), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U491 ( .A1(n630), .A2(n645), .ZN(n371) );
  NAND2_X1 U492 ( .A1(n424), .A2(n423), .ZN(n422) );
  NAND2_X1 U493 ( .A1(n406), .A2(n405), .ZN(n402) );
  AND2_X1 U494 ( .A1(n409), .A2(n560), .ZN(n424) );
  INV_X1 U495 ( .A(n553), .ZN(n393) );
  XNOR2_X1 U496 ( .A(n421), .B(n420), .ZN(n419) );
  NAND2_X1 U497 ( .A1(n372), .A2(n617), .ZN(n654) );
  XNOR2_X1 U498 ( .A(n372), .B(n744), .ZN(n743) );
  XNOR2_X1 U499 ( .A(n373), .B(n395), .ZN(n394) );
  NAND2_X1 U500 ( .A1(n376), .A2(n374), .ZN(n373) );
  XNOR2_X1 U501 ( .A(n375), .B(n366), .ZN(n374) );
  NAND2_X1 U502 ( .A1(n753), .A2(n752), .ZN(n375) );
  XNOR2_X1 U503 ( .A(n377), .B(n396), .ZN(n376) );
  NAND2_X1 U504 ( .A1(n562), .A2(n660), .ZN(n378) );
  NAND2_X1 U505 ( .A1(n361), .A2(n386), .ZN(n622) );
  NAND2_X1 U506 ( .A1(n362), .A2(n386), .ZN(n703) );
  NAND2_X1 U507 ( .A1(n382), .A2(G478), .ZN(n421) );
  NAND2_X1 U508 ( .A1(n382), .A2(G469), .ZN(n709) );
  NAND2_X1 U509 ( .A1(n599), .A2(n638), .ZN(n600) );
  NAND2_X1 U510 ( .A1(n383), .A2(n598), .ZN(n638) );
  XNOR2_X1 U511 ( .A(n385), .B(n384), .ZN(n383) );
  NOR2_X1 U512 ( .A1(n618), .A2(n617), .ZN(n390) );
  XNOR2_X2 U513 ( .A(n391), .B(n554), .ZN(n754) );
  INV_X1 U514 ( .A(KEYINPUT67), .ZN(n396) );
  NAND2_X1 U515 ( .A1(n397), .A2(n634), .ZN(n652) );
  NAND2_X1 U516 ( .A1(n401), .A2(n399), .ZN(n409) );
  NAND2_X1 U517 ( .A1(n400), .A2(n408), .ZN(n399) );
  NOR2_X1 U518 ( .A1(n751), .A2(KEYINPUT65), .ZN(n400) );
  NOR2_X1 U519 ( .A1(n360), .A2(n402), .ZN(n401) );
  NOR2_X1 U520 ( .A1(n553), .A2(n611), .ZN(n404) );
  NAND2_X1 U521 ( .A1(n404), .A2(n529), .ZN(n548) );
  NOR2_X1 U522 ( .A1(n751), .A2(n754), .ZN(n559) );
  NAND2_X1 U523 ( .A1(n410), .A2(n557), .ZN(n405) );
  INV_X1 U524 ( .A(n754), .ZN(n408) );
  XNOR2_X1 U525 ( .A(n417), .B(n416), .ZN(G63) );
  NAND2_X1 U526 ( .A1(n419), .A2(n418), .ZN(n417) );
  INV_X1 U527 ( .A(n725), .ZN(n418) );
  INV_X1 U528 ( .A(n719), .ZN(n420) );
  XNOR2_X1 U529 ( .A(n703), .B(n428), .ZN(n704) );
  NAND2_X1 U530 ( .A1(n571), .A2(n660), .ZN(n504) );
  AND2_X1 U531 ( .A1(G210), .A2(n502), .ZN(n427) );
  XOR2_X1 U532 ( .A(n702), .B(n701), .Z(n428) );
  AND2_X1 U533 ( .A1(n581), .A2(n569), .ZN(n429) );
  XNOR2_X1 U534 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U535 ( .A(n515), .B(KEYINPUT76), .ZN(n516) );
  INV_X1 U536 ( .A(n543), .ZN(n544) );
  INV_X1 U537 ( .A(KEYINPUT108), .ZN(n583) );
  INV_X1 U538 ( .A(n577), .ZN(n567) );
  INV_X1 U539 ( .A(n712), .ZN(n714) );
  INV_X1 U540 ( .A(KEYINPUT19), .ZN(n503) );
  XNOR2_X1 U541 ( .A(n716), .B(n715), .ZN(n717) );
  INV_X1 U542 ( .A(KEYINPUT63), .ZN(n625) );
  XNOR2_X1 U543 ( .A(KEYINPUT13), .B(G475), .ZN(n442) );
  XOR2_X1 U544 ( .A(KEYINPUT97), .B(KEYINPUT12), .Z(n431) );
  XNOR2_X1 U545 ( .A(KEYINPUT11), .B(KEYINPUT96), .ZN(n430) );
  XNOR2_X1 U546 ( .A(n431), .B(n430), .ZN(n435) );
  NAND2_X1 U547 ( .A1(n462), .A2(G214), .ZN(n432) );
  XNOR2_X1 U548 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U549 ( .A(n435), .B(n434), .ZN(n440) );
  XNOR2_X1 U550 ( .A(G125), .B(G146), .ZN(n489) );
  XNOR2_X1 U551 ( .A(KEYINPUT10), .B(n489), .ZN(n739) );
  INV_X1 U552 ( .A(n739), .ZN(n436) );
  XNOR2_X1 U553 ( .A(n436), .B(n494), .ZN(n438) );
  XNOR2_X1 U554 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U555 ( .A(n440), .B(n439), .ZN(n712) );
  NOR2_X1 U556 ( .A1(G902), .A2(n712), .ZN(n441) );
  XNOR2_X1 U557 ( .A(n442), .B(n441), .ZN(n542) );
  INV_X1 U558 ( .A(G128), .ZN(n443) );
  NAND2_X1 U559 ( .A1(G143), .A2(n443), .ZN(n446) );
  NAND2_X1 U560 ( .A1(n444), .A2(G128), .ZN(n445) );
  XOR2_X1 U561 ( .A(n460), .B(n498), .Z(n450) );
  XNOR2_X1 U562 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U563 ( .A(n450), .B(n449), .ZN(n456) );
  XOR2_X1 U564 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n454) );
  XOR2_X1 U565 ( .A(KEYINPUT66), .B(KEYINPUT8), .Z(n452) );
  NAND2_X1 U566 ( .A1(G234), .A2(n514), .ZN(n451) );
  XNOR2_X1 U567 ( .A(n452), .B(n451), .ZN(n474) );
  NAND2_X1 U568 ( .A1(G217), .A2(n474), .ZN(n453) );
  XNOR2_X1 U569 ( .A(n454), .B(n453), .ZN(n455) );
  XOR2_X1 U570 ( .A(n456), .B(n455), .Z(n719) );
  NOR2_X1 U571 ( .A1(n719), .A2(G902), .ZN(n457) );
  XNOR2_X1 U572 ( .A(G478), .B(n457), .ZN(n458) );
  XOR2_X1 U573 ( .A(n458), .B(KEYINPUT100), .Z(n541) );
  INV_X1 U574 ( .A(n541), .ZN(n459) );
  XNOR2_X2 U575 ( .A(n460), .B(KEYINPUT4), .ZN(n741) );
  XNOR2_X2 U576 ( .A(n741), .B(G101), .ZN(n522) );
  XOR2_X1 U577 ( .A(G116), .B(KEYINPUT3), .Z(n461) );
  XNOR2_X1 U578 ( .A(KEYINPUT70), .B(n461), .ZN(n731) );
  XNOR2_X2 U579 ( .A(n522), .B(n731), .ZN(n493) );
  XOR2_X1 U580 ( .A(KEYINPUT75), .B(KEYINPUT5), .Z(n464) );
  NAND2_X1 U581 ( .A1(n462), .A2(G210), .ZN(n463) );
  XNOR2_X1 U582 ( .A(n464), .B(n463), .ZN(n468) );
  XNOR2_X1 U583 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U584 ( .A(n469), .B(n517), .ZN(n470) );
  XNOR2_X1 U585 ( .A(n493), .B(n470), .ZN(n620) );
  BUF_X1 U586 ( .A(n562), .Z(n555) );
  NAND2_X1 U587 ( .A1(n615), .A2(G234), .ZN(n472) );
  XNOR2_X1 U588 ( .A(KEYINPUT92), .B(KEYINPUT20), .ZN(n471) );
  XNOR2_X1 U589 ( .A(n472), .B(n471), .ZN(n482) );
  NAND2_X1 U590 ( .A1(n482), .A2(G221), .ZN(n473) );
  XOR2_X1 U591 ( .A(KEYINPUT21), .B(n473), .Z(n670) );
  XNOR2_X1 U592 ( .A(KEYINPUT93), .B(n670), .ZN(n543) );
  NAND2_X1 U593 ( .A1(G221), .A2(n474), .ZN(n476) );
  XOR2_X1 U594 ( .A(n521), .B(n495), .Z(n475) );
  XNOR2_X1 U595 ( .A(n476), .B(n475), .ZN(n481) );
  XOR2_X1 U596 ( .A(KEYINPUT71), .B(KEYINPUT24), .Z(n478) );
  XNOR2_X1 U597 ( .A(n478), .B(n477), .ZN(n479) );
  XOR2_X1 U598 ( .A(n479), .B(n739), .Z(n480) );
  XNOR2_X1 U599 ( .A(n481), .B(n480), .ZN(n722) );
  NAND2_X1 U600 ( .A1(G217), .A2(n482), .ZN(n483) );
  XNOR2_X2 U601 ( .A(n485), .B(n484), .ZN(n549) );
  NOR2_X1 U602 ( .A1(n543), .A2(n576), .ZN(n569) );
  XOR2_X1 U603 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n487) );
  XNOR2_X1 U604 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U605 ( .A(n489), .B(n488), .ZN(n491) );
  NAND2_X1 U606 ( .A1(G224), .A2(n514), .ZN(n490) );
  XNOR2_X1 U607 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U608 ( .A(n493), .B(n492), .ZN(n500) );
  XOR2_X1 U609 ( .A(KEYINPUT88), .B(KEYINPUT16), .Z(n497) );
  XNOR2_X1 U610 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U611 ( .A(n497), .B(n496), .ZN(n499) );
  XNOR2_X1 U612 ( .A(n499), .B(n498), .ZN(n730) );
  XNOR2_X1 U613 ( .A(n500), .B(n730), .ZN(n700) );
  NAND2_X1 U614 ( .A1(n700), .A2(n615), .ZN(n501) );
  XNOR2_X2 U615 ( .A(n501), .B(n427), .ZN(n571) );
  NAND2_X1 U616 ( .A1(G214), .A2(n502), .ZN(n660) );
  XNOR2_X1 U617 ( .A(n505), .B(KEYINPUT14), .ZN(n506) );
  XNOR2_X1 U618 ( .A(KEYINPUT74), .B(n506), .ZN(n507) );
  NAND2_X1 U619 ( .A1(G952), .A2(n507), .ZN(n691) );
  NOR2_X1 U620 ( .A1(G953), .A2(n691), .ZN(n566) );
  AND2_X1 U621 ( .A1(n507), .A2(G953), .ZN(n508) );
  NAND2_X1 U622 ( .A1(G902), .A2(n508), .ZN(n564) );
  NOR2_X1 U623 ( .A1(G898), .A2(n564), .ZN(n509) );
  NOR2_X1 U624 ( .A1(n566), .A2(n509), .ZN(n510) );
  XNOR2_X1 U625 ( .A(n510), .B(KEYINPUT90), .ZN(n511) );
  NOR2_X1 U626 ( .A1(n601), .A2(n511), .ZN(n513) );
  XNOR2_X1 U627 ( .A(n513), .B(n512), .ZN(n546) );
  INV_X1 U628 ( .A(n546), .ZN(n535) );
  NAND2_X1 U629 ( .A1(n569), .A2(n535), .ZN(n526) );
  NAND2_X1 U630 ( .A1(G227), .A2(n514), .ZN(n515) );
  XNOR2_X1 U631 ( .A(n519), .B(n518), .ZN(n520) );
  XOR2_X1 U632 ( .A(KEYINPUT91), .B(n521), .Z(n738) );
  XNOR2_X1 U633 ( .A(n522), .B(n738), .ZN(n523) );
  XNOR2_X1 U634 ( .A(n524), .B(n523), .ZN(n706) );
  XNOR2_X1 U635 ( .A(n525), .B(KEYINPUT94), .ZN(n630) );
  NAND2_X1 U636 ( .A1(n555), .A2(n611), .ZN(n680) );
  NOR2_X1 U637 ( .A1(n526), .A2(n680), .ZN(n527) );
  XNOR2_X1 U638 ( .A(n527), .B(KEYINPUT31), .ZN(n645) );
  NAND2_X1 U639 ( .A1(n664), .A2(n528), .ZN(n561) );
  INV_X1 U640 ( .A(n611), .ZN(n674) );
  INV_X1 U641 ( .A(n529), .ZN(n590) );
  INV_X1 U642 ( .A(n569), .ZN(n681) );
  NOR2_X1 U643 ( .A1(n529), .A2(n681), .ZN(n530) );
  XOR2_X1 U644 ( .A(KEYINPUT104), .B(KEYINPUT33), .Z(n532) );
  AND2_X1 U645 ( .A1(n535), .A2(n694), .ZN(n536) );
  XNOR2_X1 U646 ( .A(n536), .B(KEYINPUT34), .ZN(n539) );
  NAND2_X1 U647 ( .A1(n541), .A2(n542), .ZN(n537) );
  XNOR2_X1 U648 ( .A(n537), .B(KEYINPUT105), .ZN(n598) );
  XOR2_X1 U649 ( .A(n598), .B(KEYINPUT77), .Z(n538) );
  NAND2_X1 U650 ( .A1(n539), .A2(n538), .ZN(n540) );
  NAND2_X1 U651 ( .A1(n749), .A2(KEYINPUT44), .ZN(n551) );
  NOR2_X1 U652 ( .A1(n542), .A2(n541), .ZN(n662) );
  XNOR2_X1 U653 ( .A(KEYINPUT83), .B(n548), .ZN(n550) );
  NAND2_X1 U654 ( .A1(n550), .A2(n549), .ZN(n626) );
  NOR2_X1 U655 ( .A1(n595), .A2(n549), .ZN(n552) );
  XNOR2_X2 U656 ( .A(KEYINPUT103), .B(n556), .ZN(n751) );
  INV_X1 U657 ( .A(KEYINPUT44), .ZN(n557) );
  NOR2_X1 U658 ( .A1(n749), .A2(KEYINPUT44), .ZN(n558) );
  NAND2_X1 U659 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U660 ( .A(KEYINPUT106), .B(KEYINPUT30), .Z(n563) );
  NOR2_X1 U661 ( .A1(G900), .A2(n564), .ZN(n565) );
  NOR2_X1 U662 ( .A1(n566), .A2(n565), .ZN(n577) );
  AND2_X1 U663 ( .A1(n568), .A2(n567), .ZN(n570) );
  NAND2_X1 U664 ( .A1(n570), .A2(n429), .ZN(n596) );
  XNOR2_X1 U665 ( .A(n571), .B(n572), .ZN(n661) );
  INV_X1 U666 ( .A(n661), .ZN(n573) );
  INV_X1 U667 ( .A(n642), .ZN(n639) );
  XOR2_X1 U668 ( .A(KEYINPUT40), .B(n575), .Z(n752) );
  NAND2_X1 U669 ( .A1(n576), .A2(n670), .ZN(n578) );
  NOR2_X1 U670 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U671 ( .A(n579), .B(KEYINPUT68), .ZN(n589) );
  NAND2_X1 U672 ( .A1(n589), .A2(n555), .ZN(n580) );
  XOR2_X1 U673 ( .A(n580), .B(KEYINPUT28), .Z(n582) );
  NAND2_X1 U674 ( .A1(n582), .A2(n581), .ZN(n602) );
  INV_X1 U675 ( .A(n602), .ZN(n587) );
  XOR2_X1 U676 ( .A(KEYINPUT41), .B(KEYINPUT109), .Z(n586) );
  NAND2_X1 U677 ( .A1(n660), .A2(n661), .ZN(n584) );
  XNOR2_X2 U678 ( .A(n584), .B(n583), .ZN(n665) );
  NAND2_X1 U679 ( .A1(n665), .A2(n662), .ZN(n585) );
  XNOR2_X2 U680 ( .A(n586), .B(n585), .ZN(n693) );
  NAND2_X1 U681 ( .A1(n587), .A2(n693), .ZN(n588) );
  XNOR2_X1 U682 ( .A(n588), .B(KEYINPUT42), .ZN(n753) );
  INV_X1 U683 ( .A(n571), .ZN(n597) );
  NAND2_X1 U684 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U685 ( .A1(n642), .A2(n591), .ZN(n592) );
  NOR2_X1 U686 ( .A1(n597), .A2(n610), .ZN(n593) );
  XOR2_X1 U687 ( .A(KEYINPUT36), .B(n593), .Z(n594) );
  NOR2_X1 U688 ( .A1(n595), .A2(n594), .ZN(n648) );
  INV_X1 U689 ( .A(KEYINPUT47), .ZN(n603) );
  OR2_X1 U690 ( .A1(n603), .A2(n664), .ZN(n599) );
  XNOR2_X1 U691 ( .A(n600), .B(KEYINPUT79), .ZN(n608) );
  NOR2_X1 U692 ( .A1(n602), .A2(n601), .ZN(n640) );
  NAND2_X1 U693 ( .A1(n664), .A2(n640), .ZN(n604) );
  NAND2_X1 U694 ( .A1(n604), .A2(n603), .ZN(n606) );
  NAND2_X1 U695 ( .A1(n640), .A2(KEYINPUT47), .ZN(n605) );
  NAND2_X1 U696 ( .A1(n606), .A2(n605), .ZN(n607) );
  NAND2_X1 U697 ( .A1(n608), .A2(n607), .ZN(n609) );
  NOR2_X1 U698 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U699 ( .A(n612), .B(KEYINPUT43), .ZN(n613) );
  NOR2_X1 U700 ( .A1(n571), .A2(n613), .ZN(n653) );
  INV_X1 U701 ( .A(KEYINPUT2), .ZN(n617) );
  XOR2_X1 U702 ( .A(KEYINPUT81), .B(n615), .Z(n616) );
  XOR2_X1 U703 ( .A(KEYINPUT62), .B(KEYINPUT85), .Z(n619) );
  XNOR2_X1 U704 ( .A(n620), .B(n619), .ZN(n621) );
  XNOR2_X1 U705 ( .A(n622), .B(n621), .ZN(n623) );
  XNOR2_X1 U706 ( .A(n625), .B(n624), .ZN(G57) );
  XNOR2_X1 U707 ( .A(G101), .B(n626), .ZN(G3) );
  NOR2_X1 U708 ( .A1(n630), .A2(n642), .ZN(n628) );
  XNOR2_X1 U709 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n627) );
  XNOR2_X1 U710 ( .A(n628), .B(n627), .ZN(n629) );
  XNOR2_X1 U711 ( .A(G104), .B(n629), .ZN(G6) );
  NOR2_X1 U712 ( .A1(n630), .A2(n646), .ZN(n632) );
  XNOR2_X1 U713 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n631) );
  XNOR2_X1 U714 ( .A(n632), .B(n631), .ZN(n633) );
  XNOR2_X1 U715 ( .A(G107), .B(n633), .ZN(G9) );
  XOR2_X1 U716 ( .A(KEYINPUT112), .B(KEYINPUT29), .Z(n636) );
  NAND2_X1 U717 ( .A1(n640), .A2(n634), .ZN(n635) );
  XNOR2_X1 U718 ( .A(n636), .B(n635), .ZN(n637) );
  XNOR2_X1 U719 ( .A(G128), .B(n637), .ZN(G30) );
  XNOR2_X1 U720 ( .A(n638), .B(G143), .ZN(G45) );
  NAND2_X1 U721 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U722 ( .A(n641), .B(G146), .ZN(G48) );
  NOR2_X1 U723 ( .A1(n642), .A2(n645), .ZN(n644) );
  XNOR2_X1 U724 ( .A(G113), .B(KEYINPUT113), .ZN(n643) );
  XNOR2_X1 U725 ( .A(n644), .B(n643), .ZN(G15) );
  NOR2_X1 U726 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U727 ( .A(G116), .B(n647), .Z(G18) );
  XNOR2_X1 U728 ( .A(n648), .B(KEYINPUT37), .ZN(n649) );
  XNOR2_X1 U729 ( .A(n649), .B(KEYINPUT114), .ZN(n650) );
  XNOR2_X1 U730 ( .A(G125), .B(n650), .ZN(G27) );
  XOR2_X1 U731 ( .A(G134), .B(KEYINPUT115), .Z(n651) );
  XNOR2_X1 U732 ( .A(n652), .B(n651), .ZN(G36) );
  XOR2_X1 U733 ( .A(G140), .B(n653), .Z(G42) );
  XNOR2_X1 U734 ( .A(n654), .B(KEYINPUT80), .ZN(n657) );
  NAND2_X1 U735 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U736 ( .A1(n659), .A2(n658), .ZN(n698) );
  OR2_X1 U737 ( .A1(n661), .A2(n660), .ZN(n663) );
  NAND2_X1 U738 ( .A1(n663), .A2(n662), .ZN(n667) );
  NAND2_X1 U739 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U740 ( .A1(n667), .A2(n666), .ZN(n668) );
  XOR2_X1 U741 ( .A(KEYINPUT119), .B(n668), .Z(n669) );
  NAND2_X1 U742 ( .A1(n669), .A2(n694), .ZN(n687) );
  NOR2_X1 U743 ( .A1(n670), .A2(n549), .ZN(n671) );
  XOR2_X1 U744 ( .A(KEYINPUT49), .B(n671), .Z(n672) );
  NOR2_X1 U745 ( .A1(n555), .A2(n672), .ZN(n673) );
  XOR2_X1 U746 ( .A(KEYINPUT116), .B(n673), .Z(n678) );
  NAND2_X1 U747 ( .A1(n681), .A2(n674), .ZN(n675) );
  XNOR2_X1 U748 ( .A(n675), .B(KEYINPUT117), .ZN(n676) );
  XNOR2_X1 U749 ( .A(KEYINPUT50), .B(n676), .ZN(n677) );
  NOR2_X1 U750 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U751 ( .A(n679), .B(KEYINPUT118), .ZN(n683) );
  NOR2_X1 U752 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U753 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U754 ( .A(KEYINPUT51), .B(n684), .ZN(n685) );
  NAND2_X1 U755 ( .A1(n685), .A2(n693), .ZN(n686) );
  NAND2_X1 U756 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U757 ( .A(n688), .B(KEYINPUT52), .ZN(n689) );
  XOR2_X1 U758 ( .A(KEYINPUT120), .B(n689), .Z(n690) );
  NOR2_X1 U759 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U760 ( .A(n692), .B(KEYINPUT121), .ZN(n696) );
  NAND2_X1 U761 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U762 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U763 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U764 ( .A(KEYINPUT122), .B(KEYINPUT54), .Z(n702) );
  XNOR2_X1 U765 ( .A(n700), .B(KEYINPUT55), .ZN(n701) );
  XNOR2_X1 U766 ( .A(KEYINPUT56), .B(n705), .ZN(G51) );
  XOR2_X1 U767 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n708) );
  XNOR2_X1 U768 ( .A(n706), .B(KEYINPUT123), .ZN(n707) );
  XNOR2_X1 U769 ( .A(n708), .B(n707), .ZN(n710) );
  XOR2_X1 U770 ( .A(n710), .B(n709), .Z(n711) );
  NOR2_X1 U771 ( .A1(n725), .A2(n711), .ZN(G54) );
  XOR2_X1 U772 ( .A(KEYINPUT59), .B(KEYINPUT87), .Z(n713) );
  XNOR2_X1 U773 ( .A(KEYINPUT60), .B(n718), .ZN(G60) );
  XOR2_X1 U774 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n721) );
  XNOR2_X1 U775 ( .A(n721), .B(n720), .ZN(n723) );
  XNOR2_X1 U776 ( .A(n723), .B(n722), .ZN(n724) );
  NOR2_X1 U777 ( .A1(n725), .A2(n724), .ZN(G66) );
  NAND2_X1 U778 ( .A1(n514), .A2(n655), .ZN(n729) );
  NAND2_X1 U779 ( .A1(G953), .A2(G224), .ZN(n726) );
  XNOR2_X1 U780 ( .A(KEYINPUT61), .B(n726), .ZN(n727) );
  NAND2_X1 U781 ( .A1(n727), .A2(G898), .ZN(n728) );
  NAND2_X1 U782 ( .A1(n729), .A2(n728), .ZN(n736) );
  XNOR2_X1 U783 ( .A(G101), .B(n730), .ZN(n732) );
  XNOR2_X1 U784 ( .A(n732), .B(n731), .ZN(n734) );
  NOR2_X1 U785 ( .A1(G898), .A2(n514), .ZN(n733) );
  NOR2_X1 U786 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U787 ( .A(n736), .B(n735), .ZN(G69) );
  XNOR2_X1 U788 ( .A(n738), .B(n737), .ZN(n740) );
  XOR2_X1 U789 ( .A(n740), .B(n739), .Z(n742) );
  XNOR2_X1 U790 ( .A(n741), .B(n742), .ZN(n744) );
  NAND2_X1 U791 ( .A1(n743), .A2(n514), .ZN(n748) );
  XNOR2_X1 U792 ( .A(G227), .B(n744), .ZN(n745) );
  NAND2_X1 U793 ( .A1(n745), .A2(G900), .ZN(n746) );
  NAND2_X1 U794 ( .A1(n746), .A2(G953), .ZN(n747) );
  NAND2_X1 U795 ( .A1(n748), .A2(n747), .ZN(G72) );
  XNOR2_X1 U796 ( .A(G122), .B(n749), .ZN(n750) );
  XNOR2_X1 U797 ( .A(n750), .B(KEYINPUT127), .ZN(G24) );
  XOR2_X1 U798 ( .A(n751), .B(G110), .Z(G12) );
  XNOR2_X1 U799 ( .A(G131), .B(n752), .ZN(G33) );
  XNOR2_X1 U800 ( .A(n753), .B(G137), .ZN(G39) );
  XOR2_X1 U801 ( .A(n754), .B(G119), .Z(G21) );
endmodule

