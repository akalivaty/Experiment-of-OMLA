//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 1 0 0 1 0 1 0 0 1 0 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 0 1 1 0 0 1 1 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:18 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1287, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(new_n201));
  XNOR2_X1  g0001(.A(new_n201), .B(KEYINPUT64), .ZN(G353));
  NOR2_X1   g0002(.A1(G97), .A2(G107), .ZN(new_n203));
  INV_X1    g0003(.A(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT65), .Z(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  AND2_X1   g0013(.A1(G68), .A2(G238), .ZN(new_n214));
  INV_X1    g0014(.A(G87), .ZN(new_n215));
  INV_X1    g0015(.A(G250), .ZN(new_n216));
  INV_X1    g0016(.A(G97), .ZN(new_n217));
  INV_X1    g0017(.A(G257), .ZN(new_n218));
  OAI22_X1  g0018(.A1(new_n215), .A2(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AOI211_X1 g0019(.A(new_n214), .B(new_n219), .C1(G107), .C2(G264), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G116), .A2(G270), .ZN(new_n221));
  AND2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G50), .ZN(new_n223));
  INV_X1    g0023(.A(G226), .ZN(new_n224));
  INV_X1    g0024(.A(G77), .ZN(new_n225));
  INV_X1    g0025(.A(G244), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(G58), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n209), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT1), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n233), .A2(new_n207), .ZN(new_n234));
  INV_X1    g0034(.A(G68), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n228), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g0036(.A1(new_n236), .A2(G50), .ZN(new_n237));
  INV_X1    g0037(.A(new_n237), .ZN(new_n238));
  AOI211_X1 g0038(.A(new_n213), .B(new_n232), .C1(new_n234), .C2(new_n238), .ZN(G361));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G264), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n241), .B(G270), .Z(new_n242));
  XNOR2_X1  g0042(.A(G238), .B(G244), .ZN(new_n243));
  XNOR2_X1  g0043(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G226), .B(G232), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n242), .B(new_n247), .ZN(G358));
  XOR2_X1   g0048(.A(G68), .B(G77), .Z(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G58), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G107), .B(G116), .Z(new_n252));
  XNOR2_X1  g0052(.A(G87), .B(G97), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  INV_X1    g0055(.A(KEYINPUT14), .ZN(new_n256));
  AND2_X1   g0056(.A1(KEYINPUT67), .A2(G41), .ZN(new_n257));
  NOR2_X1   g0057(.A1(KEYINPUT67), .A2(G41), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  OAI211_X1 g0059(.A(KEYINPUT68), .B(new_n206), .C1(new_n259), .C2(G45), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G33), .A2(G41), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(G1), .A3(G13), .ZN(new_n262));
  AND2_X1   g0062(.A1(new_n262), .A2(G274), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT67), .ZN(new_n264));
  INV_X1    g0064(.A(G41), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(KEYINPUT67), .A2(G41), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n266), .A2(new_n206), .A3(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT68), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n206), .A2(G45), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n260), .A2(new_n263), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G97), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n229), .A2(G1698), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n274), .B1(G226), .B2(G1698), .ZN(new_n275));
  INV_X1    g0075(.A(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT3), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT3), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n273), .B1(new_n275), .B2(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n233), .B1(G33), .B2(G41), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n262), .A2(G238), .A3(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n272), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  OR2_X1    g0086(.A1(new_n286), .A2(KEYINPUT13), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(KEYINPUT13), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n256), .B1(new_n289), .B2(G169), .ZN(new_n290));
  INV_X1    g0090(.A(G169), .ZN(new_n291));
  AOI211_X1 g0091(.A(KEYINPUT14), .B(new_n291), .C1(new_n287), .C2(new_n288), .ZN(new_n292));
  INV_X1    g0092(.A(G179), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n289), .A2(new_n293), .ZN(new_n294));
  NOR3_X1   g0094(.A1(new_n290), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(G20), .A2(G33), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n297), .A2(G50), .B1(G20), .B2(new_n235), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n207), .A2(G33), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n298), .B1(new_n225), .B2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(new_n233), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  XOR2_X1   g0103(.A(new_n303), .B(KEYINPUT11), .Z(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G13), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n306), .A2(G1), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n307), .A2(G20), .A3(new_n235), .ZN(new_n308));
  XOR2_X1   g0108(.A(new_n308), .B(KEYINPUT12), .Z(new_n309));
  AOI21_X1  g0109(.A(new_n302), .B1(new_n206), .B2(G20), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n309), .B1(G68), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n305), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n296), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n312), .ZN(new_n315));
  INV_X1    g0115(.A(G190), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n315), .B1(new_n316), .B2(new_n289), .ZN(new_n317));
  INV_X1    g0117(.A(G200), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n318), .B1(new_n287), .B2(new_n288), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n314), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g0121(.A(KEYINPUT3), .B(G33), .ZN(new_n322));
  INV_X1    g0122(.A(G1698), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(G222), .ZN(new_n324));
  INV_X1    g0124(.A(G223), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n322), .B(new_n324), .C1(new_n325), .C2(new_n323), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n326), .B(new_n282), .C1(G77), .C2(new_n322), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n262), .A2(new_n284), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n327), .B(new_n272), .C1(new_n224), .C2(new_n328), .ZN(new_n329));
  OR2_X1    g0129(.A1(new_n329), .A2(KEYINPUT69), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(KEYINPUT69), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n332), .A2(G169), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n223), .A2(new_n228), .A3(new_n235), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n334), .A2(G20), .B1(G150), .B2(new_n297), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n228), .A2(KEYINPUT70), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT70), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(G58), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n336), .A2(new_n338), .A3(KEYINPUT8), .ZN(new_n339));
  OR2_X1    g0139(.A1(KEYINPUT8), .A2(G58), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n335), .B1(new_n341), .B2(new_n299), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n302), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT71), .ZN(new_n344));
  XNOR2_X1  g0144(.A(new_n343), .B(new_n344), .ZN(new_n345));
  NOR3_X1   g0145(.A1(new_n306), .A2(new_n207), .A3(G1), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n223), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n310), .A2(G50), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n345), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(G179), .B1(new_n330), .B2(new_n331), .ZN(new_n351));
  NOR3_X1   g0151(.A1(new_n333), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n332), .A2(G190), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT9), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n349), .A2(new_n354), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n345), .A2(KEYINPUT9), .A3(new_n347), .A4(new_n348), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n330), .A2(G200), .A3(new_n331), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n353), .A2(new_n355), .A3(new_n356), .A4(new_n357), .ZN(new_n358));
  OR2_X1    g0158(.A1(new_n358), .A2(KEYINPUT10), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(KEYINPUT10), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n352), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(G238), .A2(G1698), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n322), .B(new_n362), .C1(new_n229), .C2(G1698), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n363), .B(new_n282), .C1(G107), .C2(new_n322), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n364), .B(new_n272), .C1(new_n226), .C2(new_n328), .ZN(new_n365));
  OR2_X1    g0165(.A1(new_n365), .A2(new_n316), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(G200), .ZN(new_n367));
  NAND2_X1  g0167(.A1(G20), .A2(G77), .ZN(new_n368));
  XNOR2_X1  g0168(.A(new_n297), .B(KEYINPUT72), .ZN(new_n369));
  XNOR2_X1  g0169(.A(KEYINPUT8), .B(G58), .ZN(new_n370));
  XOR2_X1   g0170(.A(KEYINPUT15), .B(G87), .Z(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  OAI221_X1 g0172(.A(new_n368), .B1(new_n369), .B2(new_n370), .C1(new_n372), .C2(new_n299), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n373), .A2(new_n302), .B1(new_n225), .B2(new_n346), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n310), .A2(G77), .ZN(new_n375));
  XNOR2_X1  g0175(.A(new_n375), .B(KEYINPUT73), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n366), .A2(new_n367), .A3(new_n374), .A4(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n206), .A2(G20), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n339), .A2(new_n378), .A3(new_n340), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT75), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n346), .A2(new_n302), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT75), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n339), .A2(new_n382), .A3(new_n378), .A4(new_n340), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n380), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n341), .A2(new_n346), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n325), .A2(new_n323), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n224), .A2(G1698), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n277), .A2(new_n387), .A3(new_n279), .A4(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(G33), .A2(G87), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n282), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n262), .A2(G232), .A3(new_n284), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT76), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n262), .A2(new_n284), .A3(KEYINPUT76), .A4(G232), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AND4_X1   g0197(.A1(G190), .A2(new_n272), .A3(new_n392), .A4(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n302), .ZN(new_n399));
  AOI21_X1  g0199(.A(KEYINPUT7), .B1(new_n280), .B2(new_n207), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT7), .ZN(new_n401));
  AOI211_X1 g0201(.A(new_n401), .B(G20), .C1(new_n277), .C2(new_n279), .ZN(new_n402));
  OAI21_X1  g0202(.A(G68), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(G159), .ZN(new_n404));
  NOR3_X1   g0204(.A1(new_n404), .A2(G20), .A3(G33), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n336), .A2(new_n338), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n236), .B1(new_n406), .B2(new_n235), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n405), .B1(new_n407), .B2(G20), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n403), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT16), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n399), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  AND3_X1   g0211(.A1(new_n277), .A2(new_n279), .A3(KEYINPUT74), .ZN(new_n412));
  AOI21_X1  g0212(.A(KEYINPUT74), .B1(new_n277), .B2(new_n279), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n207), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n402), .B1(new_n414), .B2(new_n401), .ZN(new_n415));
  OAI211_X1 g0215(.A(KEYINPUT16), .B(new_n408), .C1(new_n415), .C2(new_n235), .ZN(new_n416));
  AOI211_X1 g0216(.A(new_n386), .B(new_n398), .C1(new_n411), .C2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(KEYINPUT77), .A2(KEYINPUT17), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n272), .A2(new_n392), .A3(new_n397), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(G200), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT77), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT17), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n417), .A2(new_n418), .A3(new_n420), .A4(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n411), .A2(new_n416), .ZN(new_n425));
  INV_X1    g0225(.A(new_n386), .ZN(new_n426));
  INV_X1    g0226(.A(new_n398), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n425), .A2(new_n426), .A3(new_n420), .A4(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n428), .A2(new_n421), .A3(new_n422), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n424), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n425), .A2(new_n426), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n419), .A2(G169), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n272), .A2(new_n397), .A3(new_n392), .A4(G179), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n431), .A2(KEYINPUT18), .A3(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT18), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n386), .B1(new_n411), .B2(new_n416), .ZN(new_n437));
  AND2_X1   g0237(.A1(new_n432), .A2(new_n433), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n435), .A2(new_n439), .ZN(new_n440));
  OR2_X1    g0240(.A1(new_n365), .A2(G179), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n374), .A2(new_n376), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n365), .A2(new_n291), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  AND3_X1   g0244(.A1(new_n430), .A2(new_n440), .A3(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n321), .A2(new_n361), .A3(new_n377), .A4(new_n445), .ZN(new_n446));
  NOR3_X1   g0246(.A1(new_n257), .A2(new_n258), .A3(KEYINPUT5), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT5), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n206), .B(G45), .C1(new_n448), .C2(G41), .ZN(new_n449));
  OAI211_X1 g0249(.A(G270), .B(new_n262), .C1(new_n447), .C2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT84), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n449), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n266), .A2(new_n448), .A3(new_n267), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n453), .A2(new_n454), .A3(G274), .A4(new_n262), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(new_n454), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n456), .A2(KEYINPUT84), .A3(G270), .A4(new_n262), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n452), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT85), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(G264), .A2(G1698), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n322), .B(new_n461), .C1(new_n218), .C2(G1698), .ZN(new_n462));
  XOR2_X1   g0262(.A(KEYINPUT86), .B(G303), .Z(new_n463));
  OAI211_X1 g0263(.A(new_n462), .B(new_n282), .C1(new_n322), .C2(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n452), .A2(KEYINPUT85), .A3(new_n455), .A4(new_n457), .ZN(new_n465));
  AND3_X1   g0265(.A1(new_n460), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n307), .A2(G20), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n206), .A2(G33), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n399), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(G116), .ZN(new_n470));
  OAI21_X1  g0270(.A(KEYINPUT87), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT87), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n381), .A2(new_n472), .A3(G116), .A4(new_n468), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G33), .A2(G283), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n474), .B(new_n207), .C1(G33), .C2(new_n217), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n470), .A2(G20), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n475), .A2(new_n302), .A3(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT20), .ZN(new_n478));
  OR2_X1    g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n477), .A2(new_n478), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n471), .A2(new_n473), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n346), .A2(new_n470), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n466), .A2(KEYINPUT88), .A3(G179), .A4(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT88), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n460), .A2(G179), .A3(new_n464), .A4(new_n465), .ZN(new_n486));
  INV_X1    g0286(.A(new_n483), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n484), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT21), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n460), .A2(new_n464), .A3(new_n465), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n291), .B1(new_n481), .B2(new_n482), .ZN(new_n492));
  AOI211_X1 g0292(.A(KEYINPUT89), .B(new_n490), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n491), .A2(new_n492), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT89), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n490), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n489), .B1(new_n494), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n467), .A2(G97), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n469), .A2(new_n217), .ZN(new_n501));
  OAI21_X1  g0301(.A(G107), .B1(new_n400), .B2(new_n402), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n297), .A2(G77), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT6), .ZN(new_n504));
  INV_X1    g0304(.A(G107), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n217), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n504), .B1(new_n506), .B2(new_n203), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n505), .A2(KEYINPUT6), .A3(G97), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G20), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n502), .A2(new_n503), .A3(new_n510), .ZN(new_n511));
  AOI211_X1 g0311(.A(new_n500), .B(new_n501), .C1(new_n511), .C2(new_n302), .ZN(new_n512));
  OAI211_X1 g0312(.A(G257), .B(new_n262), .C1(new_n447), .C2(new_n449), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n455), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT78), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT4), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(new_n280), .B2(new_n226), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n516), .A2(G1698), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n322), .A2(G244), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n517), .A2(new_n474), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n322), .A2(G250), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n323), .B1(new_n521), .B2(KEYINPUT4), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n282), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT78), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n513), .A2(new_n524), .A3(new_n455), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n515), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G200), .ZN(new_n527));
  INV_X1    g0327(.A(new_n514), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n523), .A2(new_n528), .A3(G190), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n512), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n511), .A2(new_n302), .ZN(new_n531));
  INV_X1    g0331(.A(new_n500), .ZN(new_n532));
  INV_X1    g0332(.A(new_n501), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n523), .A2(new_n528), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n291), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n515), .A2(new_n523), .A3(new_n293), .A4(new_n525), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n534), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n530), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n322), .A2(new_n207), .A3(G68), .ZN(new_n540));
  AND2_X1   g0340(.A1(KEYINPUT80), .A2(KEYINPUT19), .ZN(new_n541));
  NOR2_X1   g0341(.A1(KEYINPUT80), .A2(KEYINPUT19), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n273), .ZN(new_n544));
  AOI21_X1  g0344(.A(G20), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n204), .A2(G87), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n540), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n299), .A2(new_n217), .ZN(new_n548));
  OAI21_X1  g0348(.A(KEYINPUT81), .B1(new_n548), .B2(new_n543), .ZN(new_n549));
  XNOR2_X1  g0349(.A(KEYINPUT80), .B(KEYINPUT19), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT81), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n550), .B(new_n551), .C1(new_n217), .C2(new_n299), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n302), .B1(new_n547), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n372), .A2(new_n346), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT82), .ZN(new_n556));
  INV_X1    g0356(.A(new_n469), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n556), .B1(new_n557), .B2(new_n371), .ZN(new_n558));
  NOR3_X1   g0358(.A1(new_n469), .A2(new_n372), .A3(KEYINPUT82), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n554), .B(new_n555), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n262), .A2(G250), .A3(new_n270), .ZN(new_n561));
  XNOR2_X1  g0361(.A(new_n561), .B(KEYINPUT79), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n206), .A2(G45), .A3(G274), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n276), .A2(new_n470), .ZN(new_n564));
  NOR2_X1   g0364(.A1(G238), .A2(G1698), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n565), .B1(new_n226), .B2(G1698), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n564), .B1(new_n566), .B2(new_n322), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n563), .B1(new_n567), .B2(new_n262), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n291), .B1(new_n562), .B2(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n562), .A2(new_n568), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n293), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n560), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n207), .B1(new_n550), .B2(new_n273), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(G87), .B2(new_n204), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n574), .A2(new_n540), .A3(new_n549), .A4(new_n552), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n575), .A2(new_n302), .B1(new_n346), .B2(new_n372), .ZN(new_n576));
  OR2_X1    g0376(.A1(new_n567), .A2(new_n262), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT79), .ZN(new_n578));
  XNOR2_X1  g0378(.A(new_n561), .B(new_n578), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n577), .A2(new_n579), .A3(G190), .A4(new_n563), .ZN(new_n580));
  OAI21_X1  g0380(.A(G200), .B1(new_n562), .B2(new_n568), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n557), .A2(G87), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n576), .A2(new_n580), .A3(new_n581), .A4(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n572), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(KEYINPUT83), .B1(new_n539), .B2(new_n584), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n572), .A2(new_n583), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT83), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n586), .A2(new_n587), .A3(new_n538), .A4(new_n530), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n491), .A2(G200), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n460), .A2(G190), .A3(new_n464), .A4(new_n465), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n590), .A2(new_n487), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(KEYINPUT90), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT90), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n590), .A2(new_n594), .A3(new_n487), .A4(new_n591), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n282), .B1(new_n453), .B2(new_n454), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n449), .B1(new_n259), .B2(new_n448), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n597), .A2(G264), .B1(new_n598), .B2(new_n263), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n216), .A2(new_n323), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n218), .A2(G1698), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n277), .A2(new_n600), .A3(new_n279), .A4(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(G33), .A2(G294), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n282), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n599), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n318), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT91), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n604), .A2(KEYINPUT91), .A3(new_n282), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n609), .A2(new_n599), .A3(new_n316), .A4(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n277), .A2(new_n279), .A3(new_n207), .A4(G87), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(KEYINPUT22), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT22), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n322), .A2(new_n615), .A3(new_n207), .A4(G87), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n614), .A2(new_n616), .B1(new_n207), .B2(new_n564), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT24), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n207), .A2(G107), .ZN(new_n619));
  XNOR2_X1  g0419(.A(new_n619), .B(KEYINPUT23), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n617), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n618), .B1(new_n617), .B2(new_n620), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n302), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n469), .A2(new_n505), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n307), .A2(new_n619), .ZN(new_n625));
  XNOR2_X1  g0425(.A(new_n625), .B(KEYINPUT25), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n612), .A2(new_n623), .A3(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n609), .A2(new_n599), .A3(new_n610), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(G169), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n599), .A2(G179), .A3(new_n605), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n623), .A2(new_n627), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NOR3_X1   g0432(.A1(new_n628), .A2(new_n632), .A3(KEYINPUT92), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT92), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n630), .A2(new_n631), .ZN(new_n635));
  INV_X1    g0435(.A(new_n622), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n617), .A2(new_n618), .A3(new_n620), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n399), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n627), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n635), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n612), .A2(new_n623), .A3(new_n627), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n634), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n633), .A2(new_n642), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n499), .A2(new_n589), .A3(new_n596), .A4(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n446), .A2(new_n644), .ZN(G372));
  INV_X1    g0445(.A(KEYINPUT93), .ZN(new_n646));
  AOI21_X1  g0446(.A(KEYINPUT18), .B1(new_n431), .B2(new_n434), .ZN(new_n647));
  NOR3_X1   g0447(.A1(new_n437), .A2(new_n438), .A3(new_n436), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n435), .A2(KEYINPUT93), .A3(new_n439), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n313), .B1(new_n320), .B2(new_n444), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n651), .B1(new_n652), .B2(new_n430), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT94), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n653), .A2(new_n654), .B1(new_n360), .B2(new_n359), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n352), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n530), .A2(new_n538), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n658), .A2(new_n641), .A3(new_n583), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n659), .B1(new_n499), .B2(new_n640), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT26), .ZN(new_n661));
  OR3_X1    g0461(.A1(new_n584), .A2(new_n661), .A3(new_n538), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n661), .B1(new_n584), .B2(new_n538), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n572), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n657), .B1(new_n446), .B2(new_n666), .ZN(new_n667));
  XOR2_X1   g0467(.A(new_n667), .B(KEYINPUT95), .Z(G369));
  AOI21_X1  g0468(.A(KEYINPUT21), .B1(new_n495), .B2(new_n496), .ZN(new_n669));
  OAI211_X1 g0469(.A(new_n488), .B(new_n484), .C1(new_n669), .C2(new_n493), .ZN(new_n670));
  INV_X1    g0470(.A(new_n307), .ZN(new_n671));
  OR3_X1    g0471(.A1(new_n671), .A2(KEYINPUT27), .A3(G20), .ZN(new_n672));
  OAI21_X1  g0472(.A(KEYINPUT27), .B1(new_n671), .B2(G20), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(G213), .A3(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(G343), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n670), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(KEYINPUT92), .B1(new_n628), .B2(new_n632), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n640), .A2(new_n634), .A3(new_n641), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n676), .B1(new_n638), .B2(new_n639), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n632), .A2(new_n676), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT97), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n682), .A2(KEYINPUT97), .A3(new_n683), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n678), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n640), .A2(new_n676), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(G330), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n483), .A2(new_n676), .ZN(new_n692));
  XOR2_X1   g0492(.A(new_n692), .B(KEYINPUT96), .Z(new_n693));
  NAND3_X1  g0493(.A1(new_n499), .A2(new_n596), .A3(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n693), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n670), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n691), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n686), .A2(new_n687), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n690), .A2(new_n699), .ZN(G399));
  INV_X1    g0500(.A(new_n210), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(new_n259), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n546), .A2(new_n470), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n702), .A2(new_n206), .A3(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n704), .B1(new_n238), .B2(new_n702), .ZN(new_n705));
  XOR2_X1   g0505(.A(new_n705), .B(KEYINPUT28), .Z(new_n706));
  OAI21_X1  g0506(.A(new_n677), .B1(new_n660), .B2(new_n665), .ZN(new_n707));
  XNOR2_X1  g0507(.A(KEYINPUT101), .B(KEYINPUT29), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n707), .A2(KEYINPUT102), .A3(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT102), .ZN(new_n711));
  AND3_X1   g0511(.A1(new_n658), .A2(new_n641), .A3(new_n583), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(new_n670), .B2(new_n632), .ZN(new_n713));
  INV_X1    g0513(.A(new_n572), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n714), .B1(new_n662), .B2(new_n663), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n676), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n711), .B1(new_n716), .B2(new_n708), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(KEYINPUT29), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n710), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n679), .A2(new_n680), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n720), .B1(new_n585), .B2(new_n588), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n721), .A2(new_n499), .A3(new_n596), .A4(new_n677), .ZN(new_n722));
  AND2_X1   g0522(.A1(new_n523), .A2(new_n528), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n597), .A2(G264), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n723), .A2(new_n724), .A3(new_n605), .A4(new_n570), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(new_n486), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT30), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(KEYINPUT98), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n570), .A2(G179), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n491), .A2(new_n730), .A3(new_n606), .A4(new_n526), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(KEYINPUT99), .ZN(new_n732));
  OAI211_X1 g0532(.A(KEYINPUT98), .B(new_n727), .C1(new_n725), .C2(new_n486), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n730), .A2(new_n526), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT99), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n734), .A2(new_n735), .A3(new_n491), .A4(new_n606), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n729), .A2(new_n732), .A3(new_n733), .A4(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n676), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT31), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT100), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n729), .A2(new_n733), .A3(new_n731), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n743), .A2(KEYINPUT31), .A3(new_n676), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n738), .A2(KEYINPUT100), .A3(new_n739), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n722), .A2(new_n742), .A3(new_n744), .A4(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G330), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n719), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n706), .B1(new_n749), .B2(G1), .ZN(G364));
  NAND3_X1  g0550(.A1(new_n210), .A2(G355), .A3(new_n322), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n412), .A2(new_n413), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n701), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(G45), .B2(new_n237), .ZN(new_n754));
  INV_X1    g0554(.A(G45), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n251), .A2(new_n755), .ZN(new_n756));
  OAI221_X1 g0556(.A(new_n751), .B1(G116), .B2(new_n210), .C1(new_n754), .C2(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n207), .B1(KEYINPUT103), .B2(new_n291), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n758), .B1(KEYINPUT103), .B2(new_n291), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n759), .A2(G1), .A3(G13), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G13), .A2(G33), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(G20), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  AND2_X1   g0565(.A1(new_n757), .A2(new_n765), .ZN(new_n766));
  XOR2_X1   g0566(.A(KEYINPUT33), .B(G317), .Z(new_n767));
  NOR2_X1   g0567(.A1(new_n293), .A2(new_n318), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n207), .A2(G190), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n767), .A2(new_n770), .ZN(new_n771));
  OR2_X1    g0571(.A1(new_n769), .A2(KEYINPUT104), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G179), .A2(G200), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n769), .A2(KEYINPUT104), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n772), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT107), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AND2_X1   g0577(.A1(new_n777), .A2(G329), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n293), .A2(G200), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n769), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G311), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n207), .B1(new_n773), .B2(G190), .ZN(new_n783));
  INV_X1    g0583(.A(G294), .ZN(new_n784));
  NAND2_X1  g0584(.A1(G20), .A2(G190), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n768), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(G326), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n280), .B1(new_n783), .B2(new_n784), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  OR4_X1    g0589(.A1(new_n771), .A2(new_n778), .A3(new_n782), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n779), .A2(new_n786), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n790), .B1(G322), .B2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G283), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n318), .A2(G179), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n772), .A2(new_n774), .A3(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(G303), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n795), .A2(new_n786), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n793), .B1(new_n794), .B2(new_n796), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n796), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(G107), .ZN(new_n801));
  INV_X1    g0601(.A(KEYINPUT105), .ZN(new_n802));
  INV_X1    g0602(.A(new_n798), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n280), .B1(new_n803), .B2(G87), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n801), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n783), .B(KEYINPUT106), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(G97), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT32), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n775), .A2(new_n404), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n808), .B1(new_n809), .B2(new_n810), .C1(new_n225), .C2(new_n780), .ZN(new_n811));
  AOI211_X1 g0611(.A(new_n805), .B(new_n811), .C1(new_n802), .C2(new_n804), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n810), .A2(new_n809), .ZN(new_n813));
  INV_X1    g0613(.A(new_n406), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n792), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n770), .ZN(new_n816));
  INV_X1    g0616(.A(new_n787), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n816), .A2(G68), .B1(new_n817), .B2(G50), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n812), .A2(new_n813), .A3(new_n815), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n799), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT108), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n766), .B1(new_n821), .B2(new_n761), .ZN(new_n822));
  INV_X1    g0622(.A(new_n702), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n306), .A2(G20), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(G45), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n823), .A2(G1), .A3(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n694), .A2(new_n696), .ZN(new_n828));
  INV_X1    g0628(.A(new_n764), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n822), .B(new_n827), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n697), .A2(new_n827), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(G330), .B2(new_n828), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n830), .A2(new_n832), .ZN(G396));
  NOR2_X1   g0633(.A1(new_n444), .A2(new_n676), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n442), .A2(new_n676), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n377), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n834), .B1(new_n444), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n707), .A2(new_n838), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n677), .B(new_n837), .C1(new_n660), .C2(new_n665), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n747), .B2(KEYINPUT109), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n747), .A2(KEYINPUT109), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n827), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n747), .A2(new_n841), .A3(KEYINPUT109), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n780), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n847), .A2(G159), .B1(new_n792), .B2(G143), .ZN(new_n848));
  INV_X1    g0648(.A(G137), .ZN(new_n849));
  INV_X1    g0649(.A(G150), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n848), .B1(new_n849), .B2(new_n787), .C1(new_n850), .C2(new_n770), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT34), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n223), .B2(new_n798), .ZN(new_n854));
  INV_X1    g0654(.A(new_n783), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n854), .B1(new_n814), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(G132), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n856), .B1(new_n235), .B2(new_n796), .C1(new_n857), .C2(new_n776), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n752), .B1(new_n851), .B2(new_n852), .ZN(new_n859));
  OAI22_X1  g0659(.A1(new_n776), .A2(new_n781), .B1(new_n797), .B2(new_n787), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(G107), .B2(new_n803), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n861), .B1(new_n215), .B2(new_n796), .C1(new_n784), .C2(new_n791), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n322), .B1(new_n816), .B2(G283), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n808), .B(new_n863), .C1(new_n470), .C2(new_n780), .ZN(new_n864));
  OAI22_X1  g0664(.A1(new_n858), .A2(new_n859), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n761), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n866), .B(new_n827), .C1(new_n763), .C2(new_n837), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n761), .A2(new_n762), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n867), .B1(new_n225), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n846), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(G384));
  OAI211_X1 g0671(.A(G116), .B(new_n234), .C1(new_n509), .C2(KEYINPUT35), .ZN(new_n872));
  XOR2_X1   g0672(.A(new_n872), .B(KEYINPUT110), .Z(new_n873));
  NAND2_X1  g0673(.A1(new_n509), .A2(KEYINPUT35), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n875), .B(KEYINPUT36), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n238), .B1(new_n406), .B2(new_n235), .ZN(new_n877));
  OAI22_X1  g0677(.A1(new_n877), .A2(new_n225), .B1(G50), .B2(new_n235), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n878), .A2(G1), .A3(new_n306), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT38), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n408), .B1(new_n415), .B2(new_n235), .ZN(new_n881));
  NOR2_X1   g0681(.A1(KEYINPUT111), .A2(KEYINPUT16), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n882), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n408), .B(new_n884), .C1(new_n415), .C2(new_n235), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n883), .A2(new_n302), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n426), .ZN(new_n887));
  INV_X1    g0687(.A(new_n674), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n889), .B1(new_n430), .B2(new_n440), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n411), .A2(new_n416), .ZN(new_n891));
  OAI22_X1  g0691(.A1(new_n891), .A2(new_n386), .B1(new_n434), .B2(new_n888), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT37), .ZN(new_n893));
  AND3_X1   g0693(.A1(new_n892), .A2(new_n893), .A3(new_n428), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n887), .A2(new_n434), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n889), .A2(new_n895), .A3(new_n428), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n894), .B1(new_n896), .B2(KEYINPUT37), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n880), .B1(new_n890), .B2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n894), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n674), .B1(new_n886), .B2(new_n426), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n438), .B1(new_n886), .B2(new_n426), .ZN(new_n901));
  INV_X1    g0701(.A(new_n428), .ZN(new_n902));
  NOR3_X1   g0702(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n899), .B1(new_n903), .B2(new_n893), .ZN(new_n904));
  INV_X1    g0704(.A(new_n440), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n424), .A2(new_n429), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n900), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n904), .A2(KEYINPUT38), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n898), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n737), .A2(KEYINPUT31), .A3(new_n676), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n740), .B(new_n910), .C1(new_n644), .C2(new_n676), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n312), .B(new_n676), .C1(new_n296), .C2(new_n320), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n312), .A2(new_n676), .ZN(new_n913));
  OAI221_X1 g0713(.A(new_n913), .B1(new_n319), .B2(new_n317), .C1(new_n295), .C2(new_n315), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n838), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n909), .A2(new_n911), .A3(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT40), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n431), .A2(new_n888), .ZN(new_n919));
  AND3_X1   g0719(.A1(new_n435), .A2(KEYINPUT93), .A3(new_n439), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT93), .B1(new_n435), .B2(new_n439), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n919), .B1(new_n922), .B2(new_n430), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n892), .A2(new_n428), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(KEYINPUT37), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n899), .A2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n880), .B1(new_n923), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n908), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n929), .A2(KEYINPUT40), .A3(new_n911), .A4(new_n915), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n918), .A2(new_n930), .A3(G330), .ZN(new_n931));
  INV_X1    g0731(.A(new_n446), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n932), .A2(G330), .A3(new_n911), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n934), .B(KEYINPUT112), .Z(new_n935));
  AND2_X1   g0735(.A1(new_n911), .A2(new_n915), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n917), .B1(new_n928), .B2(new_n908), .ZN(new_n937));
  AOI22_X1  g0737(.A1(new_n936), .A2(new_n937), .B1(new_n916), .B2(new_n917), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n938), .A2(new_n932), .A3(new_n911), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n935), .A2(new_n939), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n719), .A2(new_n446), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n657), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT39), .ZN(new_n943));
  INV_X1    g0743(.A(new_n919), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n651), .B2(new_n906), .ZN(new_n945));
  AOI21_X1  g0745(.A(KEYINPUT38), .B1(new_n945), .B2(new_n926), .ZN(new_n946));
  NOR3_X1   g0746(.A1(new_n890), .A2(new_n897), .A3(new_n880), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n943), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n314), .A2(new_n677), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n898), .A2(new_n908), .A3(KEYINPUT39), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n948), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n912), .A2(new_n914), .ZN(new_n953));
  INV_X1    g0753(.A(new_n834), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n953), .B1(new_n840), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n909), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n651), .A2(new_n674), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n952), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n942), .B(new_n958), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n940), .A2(new_n959), .B1(new_n206), .B2(new_n824), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT113), .ZN(new_n961));
  AND2_X1   g0761(.A1(new_n940), .A2(new_n959), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n876), .B(new_n879), .C1(new_n961), .C2(new_n962), .ZN(G367));
  NOR2_X1   g0763(.A1(new_n798), .A2(new_n470), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT46), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n796), .A2(new_n217), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(new_n463), .B2(new_n792), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n781), .B2(new_n787), .ZN(new_n968));
  AOI211_X1 g0768(.A(new_n752), .B(new_n968), .C1(G107), .C2(new_n855), .ZN(new_n969));
  INV_X1    g0769(.A(G317), .ZN(new_n970));
  OAI221_X1 g0770(.A(new_n969), .B1(new_n794), .B2(new_n780), .C1(new_n970), .C2(new_n775), .ZN(new_n971));
  AOI211_X1 g0771(.A(new_n965), .B(new_n971), .C1(G294), .C2(new_n816), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n806), .A2(new_n235), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(G143), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n787), .A2(new_n975), .B1(new_n780), .B2(new_n223), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n976), .B1(new_n814), .B2(new_n803), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n404), .B2(new_n770), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n322), .B1(new_n796), .B2(new_n225), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT117), .Z(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n850), .B2(new_n791), .ZN(new_n981));
  INV_X1    g0781(.A(new_n775), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n978), .B(new_n981), .C1(G137), .C2(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n972), .B1(new_n974), .B2(new_n983), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n984), .B(KEYINPUT47), .Z(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n761), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n677), .B1(new_n576), .B2(new_n582), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n714), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n584), .B2(new_n987), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n989), .A2(new_n829), .ZN(new_n990));
  INV_X1    g0790(.A(new_n753), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n765), .B1(new_n210), .B2(new_n372), .C1(new_n242), .C2(new_n991), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n986), .A2(new_n827), .A3(new_n990), .A4(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n825), .A2(G1), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n686), .A2(new_n678), .A3(new_n687), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT116), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n697), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n828), .A2(G330), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n999), .A2(new_n996), .A3(new_n995), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n678), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n687), .ZN(new_n1003));
  AOI21_X1  g0803(.A(KEYINPUT97), .B1(new_n682), .B2(new_n683), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1002), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1001), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n998), .A2(new_n688), .A3(new_n1000), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n748), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT44), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n689), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1005), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n658), .B1(new_n512), .B2(new_n677), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n538), .A2(new_n677), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1009), .B1(new_n1011), .B2(new_n1015), .ZN(new_n1016));
  AOI211_X1 g0816(.A(KEYINPUT44), .B(new_n1014), .C1(new_n1005), .C2(new_n1010), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n699), .A2(KEYINPUT115), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT45), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n1011), .B2(new_n1015), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1005), .A2(KEYINPUT45), .A3(new_n1010), .A4(new_n1014), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1018), .A2(new_n1020), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1008), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1020), .B1(new_n1018), .B2(new_n1024), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n749), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n702), .B(KEYINPUT41), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n994), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n989), .A2(KEYINPUT43), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n698), .A2(new_n1002), .A3(new_n1014), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(KEYINPUT42), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT114), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n632), .A2(new_n530), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n676), .B1(new_n1036), .B2(new_n538), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1034), .A2(new_n1035), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT42), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(new_n688), .B2(new_n1014), .ZN(new_n1041));
  OAI21_X1  g0841(.A(KEYINPUT114), .B1(new_n1041), .B2(new_n1037), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1039), .B(new_n1042), .C1(KEYINPUT42), .C2(new_n1033), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n699), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n1014), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n989), .A2(KEYINPUT43), .ZN(new_n1046));
  AND3_X1   g0846(.A1(new_n1043), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1045), .B1(new_n1043), .B2(new_n1046), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1032), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1045), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1043), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1052), .A2(new_n1031), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1049), .A2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n993), .B1(new_n1030), .B2(new_n1055), .ZN(G387));
  NAND2_X1  g0856(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n749), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1006), .A2(new_n748), .A3(new_n1007), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1058), .A2(new_n702), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1057), .A2(new_n994), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n752), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n788), .B2(new_n775), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n816), .A2(G311), .B1(new_n817), .B2(G322), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n847), .A2(new_n463), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1064), .B(new_n1065), .C1(new_n970), .C2(new_n791), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT48), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1067), .B1(new_n794), .B2(new_n783), .C1(new_n784), .C2(new_n798), .ZN(new_n1068));
  XOR2_X1   g0868(.A(KEYINPUT121), .B(KEYINPUT49), .Z(new_n1069));
  XNOR2_X1  g0869(.A(new_n1068), .B(new_n1069), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n1063), .B(new_n1070), .C1(G116), .C2(new_n800), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n775), .A2(new_n850), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n966), .B(new_n1072), .C1(new_n371), .C2(new_n807), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n803), .A2(G77), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n341), .A2(new_n770), .B1(new_n404), .B2(new_n787), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n1062), .B(new_n1075), .C1(G50), .C2(new_n792), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1073), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(G68), .B2(new_n847), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n761), .B1(new_n1071), .B2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n686), .A2(new_n687), .A3(new_n764), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n703), .A2(new_n210), .A3(new_n322), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(G107), .B2(new_n210), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT118), .Z(new_n1083));
  XNOR2_X1  g0883(.A(KEYINPUT119), .B(KEYINPUT50), .ZN(new_n1084));
  NOR3_X1   g0884(.A1(new_n370), .A2(new_n1084), .A3(G50), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1085), .A2(new_n703), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(G68), .A2(G77), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1084), .B1(new_n370), .B2(G50), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1086), .A2(new_n755), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n753), .B(new_n1089), .C1(new_n247), .C2(new_n755), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1083), .A2(new_n1090), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT120), .Z(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n765), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1079), .A2(new_n827), .A3(new_n1080), .A4(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1060), .A2(new_n1061), .A3(new_n1094), .ZN(G393));
  AND2_X1   g0895(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1096));
  OAI21_X1  g0896(.A(KEYINPUT44), .B1(new_n690), .B2(new_n1014), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1011), .A2(new_n1009), .A3(new_n1015), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NOR3_X1   g0899(.A1(new_n1096), .A2(new_n1099), .A3(new_n1044), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n699), .B1(new_n1018), .B2(new_n1024), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1058), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1019), .B1(new_n1096), .B2(new_n1099), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1103), .A2(new_n1008), .A3(new_n1025), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1102), .A2(new_n702), .A3(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1044), .B1(new_n1096), .B2(new_n1099), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1018), .A2(new_n699), .A3(new_n1024), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1106), .A2(new_n994), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n826), .B1(new_n1015), .B2(new_n764), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n765), .B1(new_n217), .B2(new_n210), .C1(new_n991), .C2(new_n254), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n770), .A2(new_n223), .B1(new_n780), .B2(new_n370), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1111), .B(KEYINPUT122), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n215), .B2(new_n796), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1062), .B1(G143), .B2(new_n982), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n807), .A2(G77), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n787), .A2(new_n850), .B1(new_n791), .B2(new_n404), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT51), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1114), .A2(new_n1115), .A3(new_n1118), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n798), .A2(new_n235), .ZN(new_n1121));
  NOR4_X1   g0921(.A1(new_n1113), .A2(new_n1119), .A3(new_n1120), .A4(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n982), .A2(G322), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n803), .A2(G283), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n322), .B1(new_n816), .B2(new_n463), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n801), .A2(new_n1123), .A3(new_n1124), .A4(new_n1125), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n787), .A2(new_n970), .B1(new_n791), .B2(new_n781), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT52), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n1127), .A2(new_n1128), .B1(new_n470), .B2(new_n783), .ZN(new_n1129));
  AND2_X1   g0929(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n780), .A2(new_n784), .ZN(new_n1131));
  NOR4_X1   g0931(.A1(new_n1126), .A2(new_n1129), .A3(new_n1130), .A4(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n761), .B1(new_n1122), .B2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1109), .A2(new_n1110), .A3(new_n1133), .ZN(new_n1134));
  AND2_X1   g0934(.A1(new_n1108), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1105), .A2(new_n1135), .ZN(G390));
  OAI211_X1 g0936(.A(new_n657), .B(new_n933), .C1(new_n446), .C2(new_n719), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n746), .A2(G330), .A3(new_n837), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n953), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n911), .A2(G330), .A3(new_n915), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n840), .A2(new_n954), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n746), .A2(G330), .A3(new_n915), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(KEYINPUT123), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT123), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n746), .A2(new_n1146), .A3(G330), .A4(new_n915), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n911), .A2(G330), .A3(new_n837), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1142), .B1(new_n1149), .B2(new_n953), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1137), .B1(new_n1143), .B2(new_n1151), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n948), .B(new_n951), .C1(new_n955), .C2(new_n950), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n946), .A2(new_n947), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n834), .B1(new_n716), .B2(new_n837), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1154), .B(new_n949), .C1(new_n1155), .C2(new_n953), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1153), .A2(new_n1156), .A3(new_n1140), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n953), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n950), .B1(new_n1142), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n948), .A2(new_n951), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1156), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1157), .B1(new_n1162), .B2(new_n1148), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n823), .B1(new_n1152), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1143), .A2(new_n1151), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1137), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n1153), .A2(new_n1156), .A3(new_n1140), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1148), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1168), .B1(new_n1161), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1167), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1164), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1163), .A2(new_n994), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1160), .A2(new_n762), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n868), .A2(new_n341), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n780), .A2(new_n217), .B1(new_n791), .B2(new_n470), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1115), .B1(new_n235), .B2(new_n796), .C1(new_n776), .C2(new_n784), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1176), .B(new_n1177), .C1(G87), .C2(new_n803), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1178), .B(new_n280), .C1(new_n505), .C2(new_n770), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(G283), .B2(new_n817), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n777), .A2(G125), .B1(G50), .B2(new_n800), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n798), .A2(new_n850), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT53), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n280), .B1(new_n816), .B2(G137), .ZN(new_n1184));
  INV_X1    g0984(.A(G128), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n787), .A2(new_n1185), .B1(new_n791), .B2(new_n857), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(new_n807), .B2(G159), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1181), .A2(new_n1183), .A3(new_n1184), .A4(new_n1187), .ZN(new_n1188));
  XOR2_X1   g0988(.A(KEYINPUT54), .B(G143), .Z(new_n1189));
  AOI21_X1  g0989(.A(new_n1188), .B1(new_n847), .B2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n761), .B1(new_n1180), .B2(new_n1190), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1174), .A2(new_n827), .A3(new_n1175), .A4(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1173), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1172), .A2(new_n1194), .ZN(G378));
  AOI22_X1  g0995(.A1(new_n1142), .A2(new_n1141), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1166), .B1(new_n1170), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n359), .A2(new_n360), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n352), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  XOR2_X1   g1000(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n350), .A2(new_n674), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1201), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n361), .A2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1202), .A2(new_n1203), .A3(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1204), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n352), .B(new_n1201), .C1(new_n359), .C2(new_n360), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n1207), .A2(new_n1208), .B1(new_n350), .B2(new_n674), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1206), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n931), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n958), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n918), .A2(new_n930), .A3(new_n1210), .A4(G330), .ZN(new_n1214));
  AND3_X1   g1014(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1213), .B1(new_n1212), .B2(new_n1214), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1197), .A2(KEYINPUT57), .A3(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT57), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1137), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1210), .B1(new_n938), .B2(G330), .ZN(new_n1221));
  AND4_X1   g1021(.A1(G330), .A2(new_n918), .A3(new_n930), .A4(new_n1210), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n958), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1219), .B1(new_n1220), .B2(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1218), .A2(new_n702), .A3(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1223), .A2(new_n994), .A3(new_n1224), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n770), .A2(new_n857), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n806), .A2(new_n850), .B1(new_n849), .B2(new_n780), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n1229), .B(new_n1230), .C1(G125), .C2(new_n817), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n803), .A2(new_n1189), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1231), .B(new_n1232), .C1(new_n1185), .C2(new_n791), .ZN(new_n1233));
  XOR2_X1   g1033(.A(KEYINPUT124), .B(KEYINPUT59), .Z(new_n1234));
  XNOR2_X1  g1034(.A(new_n1233), .B(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n982), .A2(G124), .ZN(new_n1236));
  AOI211_X1 g1036(.A(G33), .B(G41), .C1(new_n800), .C2(G159), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1235), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n223), .B1(G33), .B2(G41), .C1(new_n752), .C2(new_n259), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n974), .B1(new_n217), .B2(new_n770), .C1(new_n505), .C2(new_n791), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n796), .A2(new_n406), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n787), .A2(new_n470), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1074), .B1(new_n372), .B2(new_n780), .ZN(new_n1243));
  NOR4_X1   g1043(.A1(new_n1240), .A2(new_n1241), .A3(new_n1242), .A4(new_n1243), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n752), .A2(new_n259), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1244), .B(new_n1245), .C1(new_n794), .C2(new_n776), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT58), .ZN(new_n1247));
  OR2_X1    g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1238), .A2(new_n1239), .A3(new_n1248), .A4(new_n1249), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n1250), .A2(new_n761), .B1(new_n223), .B2(new_n868), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n827), .B(new_n1251), .C1(new_n1211), .C2(new_n763), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1228), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1227), .A2(new_n1254), .ZN(G375));
  OAI22_X1  g1055(.A1(new_n806), .A2(new_n223), .B1(new_n404), .B2(new_n798), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n1241), .B(new_n1256), .C1(G137), .C2(new_n792), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1062), .B1(new_n777), .B2(G128), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n817), .A2(G132), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n816), .A2(new_n1189), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1257), .A2(new_n1258), .A3(new_n1259), .A4(new_n1260), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n780), .A2(new_n850), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n777), .A2(G303), .B1(G77), .B2(new_n800), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n847), .A2(G107), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n322), .B1(new_n792), .B2(G283), .ZN(new_n1265));
  OAI22_X1  g1065(.A1(new_n787), .A2(new_n784), .B1(new_n770), .B2(new_n470), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1266), .B1(new_n807), .B2(new_n371), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1263), .A2(new_n1264), .A3(new_n1265), .A4(new_n1267), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n798), .A2(new_n217), .ZN(new_n1269));
  OAI22_X1  g1069(.A1(new_n1261), .A2(new_n1262), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n761), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n827), .B(new_n1271), .C1(new_n1158), .C2(new_n763), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(new_n235), .B2(new_n868), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1273), .B1(new_n1165), .B2(new_n994), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1143), .A2(new_n1151), .A3(new_n1137), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(new_n1029), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1274), .B1(new_n1276), .B2(new_n1152), .ZN(G381));
  NOR2_X1   g1077(.A1(G375), .A2(G378), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1105), .A2(new_n1135), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1029), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1280), .B1(new_n1104), .B2(new_n749), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1054), .B(new_n1049), .C1(new_n1281), .C2(new_n994), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1279), .A2(new_n1282), .A3(new_n993), .ZN(new_n1283));
  NOR3_X1   g1083(.A1(new_n1283), .A2(G396), .A3(G393), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(G381), .A2(G384), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1278), .A2(new_n1284), .A3(new_n1285), .ZN(G407));
  NAND2_X1  g1086(.A1(new_n1278), .A2(new_n675), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(G407), .A2(G213), .A3(new_n1287), .ZN(G409));
  INV_X1    g1088(.A(KEYINPUT125), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1220), .A2(new_n1225), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1253), .B1(new_n1290), .B2(new_n1029), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1289), .B1(new_n1291), .B2(G378), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1227), .A2(G378), .A3(new_n1254), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1193), .B1(new_n1171), .B2(new_n1164), .ZN(new_n1294));
  NOR3_X1   g1094(.A1(new_n1220), .A2(new_n1225), .A3(new_n1280), .ZN(new_n1295));
  OAI211_X1 g1095(.A(new_n1294), .B(KEYINPUT125), .C1(new_n1253), .C2(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1292), .A2(new_n1293), .A3(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT60), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1275), .A2(new_n1298), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1143), .A2(new_n1151), .A3(new_n1137), .A4(KEYINPUT60), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1299), .A2(new_n1167), .A3(new_n702), .A4(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n1274), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n870), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1301), .A2(G384), .A3(new_n1274), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n675), .A2(G213), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1297), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(KEYINPUT62), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1297), .A2(new_n1307), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n675), .A2(G213), .A3(G2897), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1304), .ZN(new_n1313));
  AOI21_X1  g1113(.A(G384), .B1(new_n1301), .B2(new_n1274), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1312), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1303), .A2(new_n1304), .A3(new_n1311), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1310), .A2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT61), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT62), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1297), .A2(new_n1321), .A3(new_n1306), .A4(new_n1307), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1309), .A2(new_n1319), .A3(new_n1320), .A4(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(G387), .A2(G390), .ZN(new_n1324));
  XNOR2_X1  g1124(.A(G393), .B(G396), .ZN(new_n1325));
  AND3_X1   g1125(.A1(new_n1324), .A2(new_n1283), .A3(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1325), .B1(new_n1324), .B2(new_n1283), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1323), .A2(new_n1329), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1317), .B1(new_n1307), .B2(new_n1297), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT63), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1308), .B1(new_n1331), .B2(new_n1332), .ZN(new_n1333));
  NAND4_X1  g1133(.A1(new_n1297), .A2(KEYINPUT63), .A3(new_n1306), .A4(new_n1307), .ZN(new_n1334));
  AND2_X1   g1134(.A1(new_n1334), .A2(new_n1328), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1333), .A2(new_n1335), .A3(new_n1320), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1330), .A2(new_n1336), .ZN(G405));
  NAND2_X1  g1137(.A1(G375), .A2(new_n1294), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1305), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT126), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1293), .A2(new_n1340), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1325), .ZN(new_n1342));
  NOR2_X1   g1142(.A1(G387), .A2(G390), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1279), .B1(new_n1282), .B2(new_n993), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1342), .B1(new_n1343), .B2(new_n1344), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1324), .A2(new_n1283), .A3(new_n1325), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1345), .A2(new_n1346), .A3(new_n1306), .ZN(new_n1347));
  AND3_X1   g1147(.A1(new_n1339), .A2(new_n1341), .A3(new_n1347), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1341), .B1(new_n1339), .B2(new_n1347), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1338), .B1(new_n1348), .B2(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1341), .ZN(new_n1351));
  NOR3_X1   g1151(.A1(new_n1326), .A2(new_n1327), .A3(new_n1305), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n1306), .B1(new_n1345), .B2(new_n1346), .ZN(new_n1353));
  OAI21_X1  g1153(.A(new_n1351), .B1(new_n1352), .B2(new_n1353), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1339), .A2(new_n1347), .A3(new_n1341), .ZN(new_n1355));
  NAND4_X1  g1155(.A1(new_n1354), .A2(new_n1294), .A3(G375), .A4(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1350), .A2(new_n1356), .ZN(G402));
endmodule


