

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782;

  NOR2_X1 U373 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U374 ( .A(n584), .B(n583), .ZN(n740) );
  BUF_X1 U375 ( .A(n579), .Z(n356) );
  NOR2_X1 U376 ( .A1(n416), .A2(n415), .ZN(n414) );
  AND2_X1 U377 ( .A1(n411), .A2(n410), .ZN(n409) );
  XNOR2_X1 U378 ( .A(n557), .B(KEYINPUT1), .ZN(n579) );
  AND2_X1 U379 ( .A1(n568), .A2(n365), .ZN(n359) );
  NAND2_X1 U380 ( .A1(n582), .A2(KEYINPUT105), .ZN(n426) );
  BUF_X1 U381 ( .A(n558), .Z(n728) );
  XNOR2_X1 U382 ( .A(n486), .B(n485), .ZN(n703) );
  XNOR2_X1 U383 ( .A(n446), .B(KEYINPUT64), .ZN(n447) );
  XNOR2_X1 U384 ( .A(n460), .B(n353), .ZN(n360) );
  XNOR2_X1 U385 ( .A(KEYINPUT70), .B(KEYINPUT77), .ZN(n353) );
  XNOR2_X2 U386 ( .A(n486), .B(n458), .ZN(n657) );
  XNOR2_X2 U387 ( .A(n564), .B(KEYINPUT6), .ZN(n582) );
  NAND2_X1 U388 ( .A1(n354), .A2(n409), .ZN(n415) );
  NAND2_X1 U389 ( .A1(n408), .A2(n419), .ZN(n354) );
  OR2_X2 U390 ( .A1(n657), .A2(G902), .ZN(n459) );
  NAND2_X1 U391 ( .A1(n355), .A2(n367), .ZN(n399) );
  NAND2_X1 U392 ( .A1(n395), .A2(n400), .ZN(n355) );
  XNOR2_X1 U393 ( .A(G146), .B(G125), .ZN(n494) );
  NAND2_X1 U394 ( .A1(n590), .A2(n589), .ZN(n594) );
  OR2_X1 U395 ( .A1(n541), .A2(n741), .ZN(n632) );
  XNOR2_X2 U396 ( .A(n641), .B(n640), .ZN(n645) );
  NOR2_X2 U397 ( .A1(n672), .A2(n434), .ZN(n593) );
  XNOR2_X2 U398 ( .A(n435), .B(KEYINPUT35), .ZN(n672) );
  XNOR2_X1 U399 ( .A(n548), .B(KEYINPUT0), .ZN(n572) );
  INV_X1 U400 ( .A(n742), .ZN(n746) );
  NAND2_X1 U401 ( .A1(n728), .A2(n480), .ZN(n568) );
  XNOR2_X1 U402 ( .A(G119), .B(G116), .ZN(n451) );
  INV_X2 U403 ( .A(G953), .ZN(n774) );
  NOR2_X1 U404 ( .A1(n670), .A2(n612), .ZN(n613) );
  NAND2_X1 U405 ( .A1(n414), .A2(n412), .ZN(n633) );
  AND2_X1 U406 ( .A1(n421), .A2(n419), .ZN(n416) );
  AND2_X1 U407 ( .A1(n439), .A2(n442), .ZN(n438) );
  XNOR2_X1 U408 ( .A(n444), .B(n443), .ZN(n442) );
  AND2_X1 U409 ( .A1(n588), .A2(n587), .ZN(n718) );
  BUF_X1 U410 ( .A(n541), .Z(n626) );
  XNOR2_X1 U411 ( .A(n505), .B(n504), .ZN(n541) );
  INV_X1 U412 ( .A(n702), .ZN(n358) );
  BUF_X1 U413 ( .A(n677), .Z(n764) );
  XNOR2_X2 U414 ( .A(n771), .B(G146), .ZN(n486) );
  XNOR2_X2 U415 ( .A(n499), .B(n449), .ZN(n771) );
  XNOR2_X2 U416 ( .A(n487), .B(n701), .ZN(n557) );
  NAND2_X1 U417 ( .A1(KEYINPUT47), .A2(n620), .ZN(n382) );
  XNOR2_X1 U418 ( .A(n388), .B(n538), .ZN(n769) );
  OR2_X1 U419 ( .A1(n742), .A2(n389), .ZN(n388) );
  AND2_X1 U420 ( .A1(n382), .A2(KEYINPUT79), .ZN(n378) );
  XNOR2_X1 U421 ( .A(n375), .B(n374), .ZN(n619) );
  INV_X1 U422 ( .A(KEYINPUT102), .ZN(n374) );
  OR2_X1 U423 ( .A1(n721), .A2(n718), .ZN(n375) );
  NAND2_X1 U424 ( .A1(n359), .A2(n718), .ZN(n411) );
  AND2_X1 U425 ( .A1(n718), .A2(n420), .ZN(n419) );
  INV_X1 U426 ( .A(KEYINPUT106), .ZN(n420) );
  INV_X1 U427 ( .A(KEYINPUT30), .ZN(n443) );
  XNOR2_X1 U428 ( .A(n470), .B(n469), .ZN(n558) );
  XNOR2_X1 U429 ( .A(KEYINPUT89), .B(KEYINPUT3), .ZN(n452) );
  XNOR2_X1 U430 ( .A(n392), .B(n391), .ZN(n390) );
  INV_X1 U431 ( .A(KEYINPUT28), .ZN(n391) );
  NAND2_X1 U432 ( .A1(n598), .A2(n417), .ZN(n392) );
  NOR2_X1 U433 ( .A1(n403), .A2(n635), .ZN(n402) );
  INV_X1 U434 ( .A(n589), .ZN(n403) );
  NAND2_X1 U435 ( .A1(n406), .A2(n405), .ZN(n386) );
  AND2_X1 U436 ( .A1(n768), .A2(n364), .ZN(n405) );
  NAND2_X1 U437 ( .A1(n767), .A2(n766), .ZN(n406) );
  AND2_X1 U438 ( .A1(n380), .A2(n623), .ZN(n379) );
  NAND2_X1 U439 ( .A1(G237), .A2(G234), .ZN(n473) );
  NOR2_X1 U440 ( .A1(G953), .A2(G237), .ZN(n513) );
  XNOR2_X1 U441 ( .A(G143), .B(G104), .ZN(n507) );
  XOR2_X1 U442 ( .A(G140), .B(G131), .Z(n508) );
  XNOR2_X1 U443 ( .A(G122), .B(G113), .ZN(n509) );
  XOR2_X1 U444 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n510) );
  XOR2_X1 U445 ( .A(G137), .B(G140), .Z(n481) );
  XNOR2_X1 U446 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n493) );
  INV_X1 U447 ( .A(KEYINPUT105), .ZN(n423) );
  OR2_X1 U448 ( .A1(n718), .A2(n420), .ZN(n410) );
  XNOR2_X1 U449 ( .A(n370), .B(n369), .ZN(n526) );
  INV_X1 U450 ( .A(KEYINPUT8), .ZN(n369) );
  NAND2_X1 U451 ( .A1(n774), .A2(G234), .ZN(n370) );
  XOR2_X1 U452 ( .A(KEYINPUT99), .B(KEYINPUT9), .Z(n523) );
  XNOR2_X1 U453 ( .A(KEYINPUT98), .B(KEYINPUT7), .ZN(n522) );
  XNOR2_X1 U454 ( .A(G134), .B(G107), .ZN(n520) );
  XOR2_X1 U455 ( .A(G122), .B(G116), .Z(n521) );
  NAND2_X1 U456 ( .A1(n373), .A2(n366), .ZN(n372) );
  NAND2_X1 U457 ( .A1(n438), .A2(n573), .ZN(n566) );
  NAND2_X1 U458 ( .A1(n591), .A2(KEYINPUT32), .ZN(n433) );
  INV_X1 U459 ( .A(n594), .ZN(n431) );
  BUF_X1 U460 ( .A(n564), .Z(n598) );
  XNOR2_X1 U461 ( .A(KEYINPUT72), .B(KEYINPUT16), .ZN(n488) );
  NOR2_X1 U462 ( .A1(n774), .A2(G952), .ZN(n707) );
  XNOR2_X1 U463 ( .A(n540), .B(n539), .ZN(n612) );
  NAND2_X1 U464 ( .A1(n363), .A2(n387), .ZN(n540) );
  INV_X1 U465 ( .A(n625), .ZN(n436) );
  XNOR2_X1 U466 ( .A(n586), .B(n437), .ZN(n428) );
  NAND2_X1 U467 ( .A1(n432), .A2(n429), .ZN(n671) );
  NAND2_X1 U468 ( .A1(n431), .A2(n430), .ZN(n429) );
  AND2_X1 U469 ( .A1(n427), .A2(n433), .ZN(n432) );
  NOR2_X1 U470 ( .A1(n591), .A2(KEYINPUT32), .ZN(n430) );
  XNOR2_X1 U471 ( .A(n376), .B(KEYINPUT101), .ZN(n721) );
  XNOR2_X1 U472 ( .A(n404), .B(KEYINPUT86), .ZN(n595) );
  INV_X1 U473 ( .A(KEYINPUT53), .ZN(n383) );
  XNOR2_X1 U474 ( .A(KEYINPUT15), .B(G902), .ZN(n648) );
  XOR2_X1 U475 ( .A(KEYINPUT24), .B(G119), .Z(n361) );
  INV_X1 U476 ( .A(n568), .ZN(n417) );
  NOR2_X1 U477 ( .A1(n441), .A2(n440), .ZN(n624) );
  AND2_X1 U478 ( .A1(n618), .A2(n382), .ZN(n362) );
  XNOR2_X1 U479 ( .A(n562), .B(n561), .ZN(n573) );
  AND2_X1 U480 ( .A1(n390), .A2(n560), .ZN(n363) );
  OR2_X1 U481 ( .A1(n770), .A2(n769), .ZN(n364) );
  AND2_X1 U482 ( .A1(n420), .A2(KEYINPUT105), .ZN(n365) );
  AND2_X1 U483 ( .A1(n763), .A2(KEYINPUT76), .ZN(n366) );
  AND2_X1 U484 ( .A1(n501), .A2(KEYINPUT2), .ZN(n367) );
  INV_X2 U485 ( .A(n700), .ZN(n689) );
  NAND2_X1 U486 ( .A1(n638), .A2(n639), .ZN(n641) );
  XNOR2_X2 U487 ( .A(n368), .B(KEYINPUT65), .ZN(n700) );
  NAND2_X1 U488 ( .A1(n397), .A2(n399), .ZN(n368) );
  INV_X1 U489 ( .A(n647), .ZN(n373) );
  NAND2_X2 U490 ( .A1(n645), .A2(n644), .ZN(n647) );
  NOR2_X1 U491 ( .A1(n677), .A2(n648), .ZN(n398) );
  NAND2_X1 U492 ( .A1(n372), .A2(n371), .ZN(n401) );
  NAND2_X1 U493 ( .A1(n647), .A2(n646), .ZN(n371) );
  NAND2_X1 U494 ( .A1(n377), .A2(n535), .ZN(n376) );
  INV_X1 U495 ( .A(n587), .ZN(n377) );
  NAND2_X1 U496 ( .A1(n618), .A2(n378), .ZN(n380) );
  NAND2_X1 U497 ( .A1(n381), .A2(n379), .ZN(n629) );
  NAND2_X1 U498 ( .A1(n615), .A2(n362), .ZN(n381) );
  XNOR2_X2 U499 ( .A(n459), .B(G472), .ZN(n564) );
  XNOR2_X1 U500 ( .A(n384), .B(n383), .ZN(G75) );
  NAND2_X1 U501 ( .A1(n385), .A2(n774), .ZN(n384) );
  XNOR2_X1 U502 ( .A(n386), .B(KEYINPUT121), .ZN(n385) );
  INV_X1 U503 ( .A(n647), .ZN(n400) );
  INV_X1 U504 ( .A(n769), .ZN(n387) );
  NAND2_X1 U505 ( .A1(n748), .A2(n745), .ZN(n389) );
  XNOR2_X2 U506 ( .A(n394), .B(n393), .ZN(n490) );
  XNOR2_X2 U507 ( .A(G110), .B(G107), .ZN(n393) );
  XNOR2_X2 U508 ( .A(G104), .B(G101), .ZN(n394) );
  INV_X1 U509 ( .A(n677), .ZN(n395) );
  NAND2_X1 U510 ( .A1(n401), .A2(n398), .ZN(n397) );
  NAND2_X1 U511 ( .A1(n590), .A2(n402), .ZN(n404) );
  XNOR2_X2 U512 ( .A(n554), .B(n553), .ZN(n590) );
  AND2_X1 U513 ( .A1(n631), .A2(n630), .ZN(n639) );
  INV_X1 U514 ( .A(n426), .ZN(n408) );
  NAND2_X1 U515 ( .A1(n568), .A2(KEYINPUT105), .ZN(n425) );
  NAND2_X1 U516 ( .A1(n413), .A2(n418), .ZN(n412) );
  INV_X1 U517 ( .A(n421), .ZN(n413) );
  NAND2_X1 U518 ( .A1(n426), .A2(n425), .ZN(n424) );
  NAND2_X1 U519 ( .A1(n417), .A2(n423), .ZN(n422) );
  NOR2_X1 U520 ( .A1(n424), .A2(n420), .ZN(n418) );
  NOR2_X1 U521 ( .A1(n582), .A2(n422), .ZN(n421) );
  NAND2_X1 U522 ( .A1(n594), .A2(KEYINPUT32), .ZN(n427) );
  NAND2_X1 U523 ( .A1(n428), .A2(n436), .ZN(n435) );
  NAND2_X1 U524 ( .A1(n671), .A2(n592), .ZN(n434) );
  INV_X1 U525 ( .A(KEYINPUT34), .ZN(n437) );
  NAND2_X1 U526 ( .A1(n573), .A2(n563), .ZN(n440) );
  INV_X1 U527 ( .A(n442), .ZN(n441) );
  AND2_X1 U528 ( .A1(n746), .A2(n563), .ZN(n439) );
  NAND2_X1 U529 ( .A1(n564), .A2(n745), .ZN(n444) );
  XOR2_X1 U530 ( .A(KEYINPUT87), .B(KEYINPUT36), .Z(n445) );
  INV_X1 U531 ( .A(KEYINPUT33), .ZN(n583) );
  BUF_X1 U532 ( .A(n663), .Z(n665) );
  XNOR2_X1 U533 ( .A(n649), .B(KEYINPUT59), .ZN(n650) );
  INV_X1 U534 ( .A(n356), .ZN(n635) );
  XNOR2_X2 U535 ( .A(KEYINPUT68), .B(KEYINPUT4), .ZN(n446) );
  XNOR2_X1 U536 ( .A(G143), .B(G128), .ZN(n528) );
  XNOR2_X2 U537 ( .A(n447), .B(n528), .ZN(n499) );
  INV_X1 U538 ( .A(G134), .ZN(n448) );
  XNOR2_X1 U539 ( .A(n448), .B(G131), .ZN(n449) );
  XNOR2_X1 U540 ( .A(G113), .B(KEYINPUT69), .ZN(n450) );
  XNOR2_X1 U541 ( .A(n451), .B(n450), .ZN(n453) );
  XNOR2_X1 U542 ( .A(n453), .B(n452), .ZN(n491) );
  NAND2_X1 U543 ( .A1(n513), .A2(G210), .ZN(n454) );
  XNOR2_X1 U544 ( .A(n454), .B(G137), .ZN(n456) );
  XNOR2_X1 U545 ( .A(G101), .B(KEYINPUT5), .ZN(n455) );
  XNOR2_X1 U546 ( .A(n456), .B(n455), .ZN(n457) );
  XOR2_X1 U547 ( .A(n491), .B(n457), .Z(n458) );
  XNOR2_X1 U548 ( .A(KEYINPUT95), .B(KEYINPUT23), .ZN(n460) );
  XNOR2_X1 U549 ( .A(G128), .B(G110), .ZN(n461) );
  XNOR2_X1 U550 ( .A(n361), .B(n461), .ZN(n462) );
  XNOR2_X1 U551 ( .A(n360), .B(n462), .ZN(n464) );
  NAND2_X1 U552 ( .A1(G221), .A2(n526), .ZN(n463) );
  XNOR2_X1 U553 ( .A(n464), .B(n463), .ZN(n466) );
  XNOR2_X1 U554 ( .A(n494), .B(KEYINPUT10), .ZN(n515) );
  INV_X1 U555 ( .A(n481), .ZN(n465) );
  XNOR2_X1 U556 ( .A(n515), .B(n465), .ZN(n772) );
  XNOR2_X1 U557 ( .A(n466), .B(n772), .ZN(n691) );
  INV_X1 U558 ( .A(G902), .ZN(n533) );
  NAND2_X1 U559 ( .A1(n691), .A2(n533), .ZN(n470) );
  NAND2_X1 U560 ( .A1(G234), .A2(n648), .ZN(n467) );
  XNOR2_X1 U561 ( .A(KEYINPUT20), .B(n467), .ZN(n471) );
  NAND2_X1 U562 ( .A1(G217), .A2(n471), .ZN(n468) );
  XNOR2_X1 U563 ( .A(n468), .B(KEYINPUT25), .ZN(n469) );
  NAND2_X1 U564 ( .A1(G221), .A2(n471), .ZN(n472) );
  XNOR2_X1 U565 ( .A(n472), .B(KEYINPUT21), .ZN(n727) );
  XOR2_X1 U566 ( .A(KEYINPUT73), .B(KEYINPUT14), .Z(n474) );
  XNOR2_X1 U567 ( .A(n474), .B(n473), .ZN(n477) );
  NAND2_X1 U568 ( .A1(n477), .A2(G902), .ZN(n475) );
  XNOR2_X1 U569 ( .A(n475), .B(KEYINPUT91), .ZN(n543) );
  NAND2_X1 U570 ( .A1(G953), .A2(n543), .ZN(n476) );
  OR2_X1 U571 ( .A1(n476), .A2(G900), .ZN(n478) );
  AND2_X1 U572 ( .A1(G952), .A2(n477), .ZN(n758) );
  NAND2_X1 U573 ( .A1(n758), .A2(n774), .ZN(n544) );
  NAND2_X1 U574 ( .A1(n478), .A2(n544), .ZN(n563) );
  INV_X1 U575 ( .A(n563), .ZN(n479) );
  NOR2_X1 U576 ( .A1(n727), .A2(n479), .ZN(n480) );
  NAND2_X1 U577 ( .A1(G227), .A2(n774), .ZN(n483) );
  XOR2_X1 U578 ( .A(n481), .B(KEYINPUT94), .Z(n482) );
  XNOR2_X1 U579 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U580 ( .A(n490), .B(n484), .ZN(n485) );
  OR2_X2 U581 ( .A1(n703), .A2(G902), .ZN(n487) );
  INV_X1 U582 ( .A(G469), .ZN(n701) );
  XNOR2_X1 U583 ( .A(n488), .B(G122), .ZN(n489) );
  XNOR2_X1 U584 ( .A(n490), .B(n489), .ZN(n492) );
  XNOR2_X1 U585 ( .A(n492), .B(n491), .ZN(n685) );
  XNOR2_X1 U586 ( .A(n494), .B(n493), .ZN(n497) );
  NAND2_X1 U587 ( .A1(n774), .A2(G224), .ZN(n495) );
  XNOR2_X1 U588 ( .A(n495), .B(KEYINPUT90), .ZN(n496) );
  XNOR2_X1 U589 ( .A(n496), .B(n497), .ZN(n498) );
  XNOR2_X1 U590 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U591 ( .A(n685), .B(n500), .ZN(n663) );
  INV_X1 U592 ( .A(n648), .ZN(n501) );
  OR2_X2 U593 ( .A1(n663), .A2(n501), .ZN(n505) );
  NOR2_X1 U594 ( .A1(G237), .A2(G902), .ZN(n502) );
  XNOR2_X1 U595 ( .A(KEYINPUT75), .B(n502), .ZN(n536) );
  NAND2_X1 U596 ( .A1(n536), .A2(G210), .ZN(n503) );
  XNOR2_X1 U597 ( .A(n503), .B(KEYINPUT78), .ZN(n504) );
  INV_X1 U598 ( .A(KEYINPUT38), .ZN(n506) );
  XNOR2_X1 U599 ( .A(n626), .B(n506), .ZN(n742) );
  XNOR2_X1 U600 ( .A(n508), .B(n507), .ZN(n512) );
  XNOR2_X1 U601 ( .A(n510), .B(n509), .ZN(n511) );
  XOR2_X1 U602 ( .A(n512), .B(n511), .Z(n517) );
  AND2_X1 U603 ( .A1(n513), .A2(G214), .ZN(n514) );
  XNOR2_X1 U604 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U605 ( .A(n517), .B(n516), .ZN(n649) );
  NAND2_X1 U606 ( .A1(n649), .A2(n533), .ZN(n519) );
  XOR2_X1 U607 ( .A(KEYINPUT13), .B(G475), .Z(n518) );
  XNOR2_X1 U608 ( .A(n519), .B(n518), .ZN(n588) );
  INV_X1 U609 ( .A(n588), .ZN(n535) );
  XNOR2_X1 U610 ( .A(n521), .B(n520), .ZN(n525) );
  XNOR2_X1 U611 ( .A(n523), .B(n522), .ZN(n524) );
  XOR2_X1 U612 ( .A(n525), .B(n524), .Z(n532) );
  NAND2_X1 U613 ( .A1(G217), .A2(n526), .ZN(n530) );
  INV_X1 U614 ( .A(KEYINPUT100), .ZN(n527) );
  XNOR2_X1 U615 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U616 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U617 ( .A(n532), .B(n531), .ZN(n696) );
  NAND2_X1 U618 ( .A1(n696), .A2(n533), .ZN(n534) );
  INV_X1 U619 ( .A(G478), .ZN(n695) );
  XNOR2_X1 U620 ( .A(n534), .B(n695), .ZN(n587) );
  AND2_X1 U621 ( .A1(n535), .A2(n587), .ZN(n748) );
  AND2_X1 U622 ( .A1(n536), .A2(G214), .ZN(n741) );
  INV_X1 U623 ( .A(n741), .ZN(n745) );
  INV_X1 U624 ( .A(KEYINPUT108), .ZN(n537) );
  XNOR2_X1 U625 ( .A(n537), .B(KEYINPUT41), .ZN(n538) );
  XNOR2_X1 U626 ( .A(KEYINPUT109), .B(KEYINPUT42), .ZN(n539) );
  XOR2_X1 U627 ( .A(G137), .B(n612), .Z(G39) );
  XNOR2_X1 U628 ( .A(KEYINPUT66), .B(KEYINPUT19), .ZN(n542) );
  XNOR2_X2 U629 ( .A(n632), .B(n542), .ZN(n616) );
  NOR2_X1 U630 ( .A1(G898), .A2(n774), .ZN(n686) );
  NAND2_X1 U631 ( .A1(n543), .A2(n686), .ZN(n545) );
  NAND2_X1 U632 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U633 ( .A(n546), .B(KEYINPUT92), .ZN(n547) );
  NAND2_X1 U634 ( .A1(n616), .A2(n547), .ZN(n548) );
  INV_X1 U635 ( .A(n727), .ZN(n549) );
  NAND2_X1 U636 ( .A1(n748), .A2(n549), .ZN(n551) );
  INV_X1 U637 ( .A(KEYINPUT103), .ZN(n550) );
  XNOR2_X1 U638 ( .A(n551), .B(n550), .ZN(n552) );
  OR2_X2 U639 ( .A1(n572), .A2(n552), .ZN(n554) );
  XNOR2_X1 U640 ( .A(KEYINPUT71), .B(KEYINPUT22), .ZN(n553) );
  INV_X1 U641 ( .A(n598), .ZN(n731) );
  NAND2_X1 U642 ( .A1(n731), .A2(n728), .ZN(n555) );
  NOR2_X1 U643 ( .A1(n635), .A2(n555), .ZN(n556) );
  NAND2_X1 U644 ( .A1(n590), .A2(n556), .ZN(n592) );
  XNOR2_X1 U645 ( .A(n592), .B(G110), .ZN(G12) );
  INV_X1 U646 ( .A(n557), .ZN(n560) );
  OR2_X1 U647 ( .A1(n558), .A2(n727), .ZN(n725) );
  INV_X1 U648 ( .A(n725), .ZN(n559) );
  NAND2_X1 U649 ( .A1(n560), .A2(n559), .ZN(n562) );
  INV_X1 U650 ( .A(KEYINPUT96), .ZN(n561) );
  XNOR2_X1 U651 ( .A(KEYINPUT85), .B(KEYINPUT39), .ZN(n565) );
  XNOR2_X1 U652 ( .A(n566), .B(n565), .ZN(n608) );
  INV_X1 U653 ( .A(n721), .ZN(n567) );
  OR2_X1 U654 ( .A1(n608), .A2(n567), .ZN(n642) );
  XNOR2_X1 U655 ( .A(n642), .B(G134), .ZN(G36) );
  NOR2_X1 U656 ( .A1(n633), .A2(n741), .ZN(n569) );
  NAND2_X1 U657 ( .A1(n569), .A2(n356), .ZN(n570) );
  XNOR2_X1 U658 ( .A(n570), .B(KEYINPUT43), .ZN(n571) );
  NAND2_X1 U659 ( .A1(n571), .A2(n626), .ZN(n643) );
  XNOR2_X1 U660 ( .A(n643), .B(G140), .ZN(G42) );
  XNOR2_X1 U661 ( .A(n572), .B(KEYINPUT93), .ZN(n585) );
  INV_X1 U662 ( .A(n585), .ZN(n575) );
  INV_X1 U663 ( .A(n573), .ZN(n574) );
  NOR2_X1 U664 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U665 ( .A(n576), .B(KEYINPUT97), .ZN(n577) );
  NOR2_X1 U666 ( .A1(n577), .A2(n598), .ZN(n709) );
  NAND2_X1 U667 ( .A1(n709), .A2(n718), .ZN(n578) );
  XNOR2_X1 U668 ( .A(n578), .B(G104), .ZN(G6) );
  NOR2_X1 U669 ( .A1(n579), .A2(n725), .ZN(n581) );
  INV_X1 U670 ( .A(KEYINPUT74), .ZN(n580) );
  XNOR2_X1 U671 ( .A(n581), .B(n580), .ZN(n597) );
  BUF_X1 U672 ( .A(n582), .Z(n589) );
  NOR2_X2 U673 ( .A1(n597), .A2(n589), .ZN(n584) );
  NAND2_X1 U674 ( .A1(n740), .A2(n585), .ZN(n586) );
  NAND2_X1 U675 ( .A1(n588), .A2(n377), .ZN(n625) );
  NAND2_X1 U676 ( .A1(n635), .A2(n728), .ZN(n591) );
  XNOR2_X1 U677 ( .A(n593), .B(KEYINPUT44), .ZN(n605) );
  NOR2_X1 U678 ( .A1(n595), .A2(n728), .ZN(n596) );
  XNOR2_X1 U679 ( .A(n596), .B(KEYINPUT104), .ZN(n656) );
  INV_X1 U680 ( .A(n597), .ZN(n599) );
  NAND2_X1 U681 ( .A1(n599), .A2(n598), .ZN(n736) );
  NOR2_X1 U682 ( .A1(n736), .A2(n572), .ZN(n600) );
  XOR2_X1 U683 ( .A(KEYINPUT31), .B(n600), .Z(n722) );
  NOR2_X1 U684 ( .A1(n709), .A2(n722), .ZN(n602) );
  XNOR2_X1 U685 ( .A(n619), .B(KEYINPUT80), .ZN(n601) );
  NOR2_X1 U686 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U687 ( .A1(n656), .A2(n603), .ZN(n604) );
  NAND2_X1 U688 ( .A1(n605), .A2(n604), .ZN(n607) );
  XNOR2_X1 U689 ( .A(KEYINPUT83), .B(KEYINPUT45), .ZN(n606) );
  XNOR2_X2 U690 ( .A(n607), .B(n606), .ZN(n677) );
  INV_X1 U691 ( .A(n608), .ZN(n609) );
  NAND2_X1 U692 ( .A1(n609), .A2(n718), .ZN(n611) );
  INV_X1 U693 ( .A(KEYINPUT40), .ZN(n610) );
  XNOR2_X1 U694 ( .A(n611), .B(n610), .ZN(n670) );
  XNOR2_X1 U695 ( .A(n613), .B(KEYINPUT46), .ZN(n631) );
  XOR2_X1 U696 ( .A(KEYINPUT80), .B(n619), .Z(n615) );
  INV_X1 U697 ( .A(KEYINPUT47), .ZN(n614) );
  INV_X1 U698 ( .A(KEYINPUT79), .ZN(n620) );
  NAND2_X1 U699 ( .A1(n363), .A2(n616), .ZN(n713) );
  NAND2_X1 U700 ( .A1(n614), .A2(KEYINPUT79), .ZN(n617) );
  NAND2_X1 U701 ( .A1(n713), .A2(n617), .ZN(n618) );
  INV_X1 U702 ( .A(n619), .ZN(n744) );
  NAND2_X1 U703 ( .A1(n713), .A2(n620), .ZN(n621) );
  NAND2_X1 U704 ( .A1(n744), .A2(n621), .ZN(n622) );
  NAND2_X1 U705 ( .A1(n622), .A2(KEYINPUT47), .ZN(n623) );
  NOR2_X1 U706 ( .A1(n626), .A2(n625), .ZN(n627) );
  NAND2_X1 U707 ( .A1(n624), .A2(n627), .ZN(n628) );
  XNOR2_X1 U708 ( .A(n628), .B(KEYINPUT107), .ZN(n781) );
  NOR2_X1 U709 ( .A1(n629), .A2(n781), .ZN(n630) );
  XNOR2_X1 U710 ( .A(n634), .B(n445), .ZN(n636) );
  NAND2_X1 U711 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X2 U712 ( .A(n637), .B(KEYINPUT110), .ZN(n675) );
  XNOR2_X1 U713 ( .A(n675), .B(KEYINPUT84), .ZN(n638) );
  INV_X1 U714 ( .A(KEYINPUT48), .ZN(n640) );
  AND2_X1 U715 ( .A1(n643), .A2(n642), .ZN(n644) );
  INV_X1 U716 ( .A(KEYINPUT2), .ZN(n763) );
  INV_X1 U717 ( .A(KEYINPUT76), .ZN(n646) );
  NAND2_X1 U718 ( .A1(n689), .A2(G475), .ZN(n651) );
  XNOR2_X1 U719 ( .A(n651), .B(n650), .ZN(n652) );
  NOR2_X1 U720 ( .A1(n652), .A2(n707), .ZN(n654) );
  XOR2_X1 U721 ( .A(KEYINPUT67), .B(KEYINPUT60), .Z(n653) );
  XNOR2_X1 U722 ( .A(n654), .B(n653), .ZN(G60) );
  XNOR2_X1 U723 ( .A(G101), .B(KEYINPUT111), .ZN(n655) );
  XNOR2_X1 U724 ( .A(n656), .B(n655), .ZN(G3) );
  NAND2_X1 U725 ( .A1(n689), .A2(G472), .ZN(n659) );
  XNOR2_X1 U726 ( .A(n657), .B(KEYINPUT62), .ZN(n658) );
  XNOR2_X1 U727 ( .A(n659), .B(n658), .ZN(n660) );
  NOR2_X1 U728 ( .A1(n660), .A2(n707), .ZN(n662) );
  XOR2_X1 U729 ( .A(KEYINPUT88), .B(KEYINPUT63), .Z(n661) );
  XNOR2_X1 U730 ( .A(n662), .B(n661), .ZN(G57) );
  NAND2_X1 U731 ( .A1(n689), .A2(G210), .ZN(n667) );
  XOR2_X1 U732 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n664) );
  XNOR2_X1 U733 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U734 ( .A(n667), .B(n666), .ZN(n668) );
  NOR2_X1 U735 ( .A1(n668), .A2(n707), .ZN(n669) );
  XNOR2_X1 U736 ( .A(n669), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U737 ( .A(n670), .B(G131), .Z(G33) );
  XNOR2_X1 U738 ( .A(n671), .B(G119), .ZN(G21) );
  XOR2_X1 U739 ( .A(n672), .B(G122), .Z(G24) );
  XOR2_X1 U740 ( .A(KEYINPUT115), .B(KEYINPUT37), .Z(n674) );
  XNOR2_X1 U741 ( .A(G125), .B(KEYINPUT116), .ZN(n673) );
  XNOR2_X1 U742 ( .A(n674), .B(n673), .ZN(n676) );
  XOR2_X1 U743 ( .A(n676), .B(n675), .Z(G27) );
  NOR2_X1 U744 ( .A1(n764), .A2(G953), .ZN(n678) );
  XOR2_X1 U745 ( .A(KEYINPUT126), .B(n678), .Z(n683) );
  XOR2_X1 U746 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n680) );
  NAND2_X1 U747 ( .A1(G224), .A2(G953), .ZN(n679) );
  XNOR2_X1 U748 ( .A(n680), .B(n679), .ZN(n681) );
  NAND2_X1 U749 ( .A1(n681), .A2(G898), .ZN(n682) );
  NAND2_X1 U750 ( .A1(n683), .A2(n682), .ZN(n684) );
  XOR2_X1 U751 ( .A(n684), .B(KEYINPUT127), .Z(n688) );
  NOR2_X1 U752 ( .A1(n685), .A2(n686), .ZN(n687) );
  XNOR2_X1 U753 ( .A(n688), .B(n687), .ZN(G69) );
  NAND2_X1 U754 ( .A1(n358), .A2(G217), .ZN(n693) );
  XNOR2_X1 U755 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n690) );
  XNOR2_X1 U756 ( .A(n691), .B(n690), .ZN(n692) );
  XNOR2_X1 U757 ( .A(n693), .B(n692), .ZN(n694) );
  NOR2_X1 U758 ( .A1(n694), .A2(n707), .ZN(G66) );
  NOR2_X1 U759 ( .A1(n700), .A2(n695), .ZN(n697) );
  XNOR2_X1 U760 ( .A(n697), .B(n696), .ZN(n698) );
  NOR2_X1 U761 ( .A1(n698), .A2(n707), .ZN(n699) );
  XNOR2_X1 U762 ( .A(n699), .B(KEYINPUT122), .ZN(G63) );
  BUF_X1 U763 ( .A(n700), .Z(n702) );
  NOR2_X1 U764 ( .A1(n702), .A2(n701), .ZN(n706) );
  XNOR2_X1 U765 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n704) );
  XNOR2_X1 U766 ( .A(n703), .B(n704), .ZN(n705) );
  XNOR2_X1 U767 ( .A(n706), .B(n705), .ZN(n708) );
  NOR2_X1 U768 ( .A1(n708), .A2(n707), .ZN(G54) );
  NAND2_X1 U769 ( .A1(n709), .A2(n721), .ZN(n711) );
  XOR2_X1 U770 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n710) );
  XNOR2_X1 U771 ( .A(n711), .B(n710), .ZN(n712) );
  XNOR2_X1 U772 ( .A(G107), .B(n712), .ZN(G9) );
  XOR2_X1 U773 ( .A(G128), .B(KEYINPUT29), .Z(n715) );
  INV_X1 U774 ( .A(n713), .ZN(n716) );
  NAND2_X1 U775 ( .A1(n716), .A2(n721), .ZN(n714) );
  XNOR2_X1 U776 ( .A(n715), .B(n714), .ZN(G30) );
  NAND2_X1 U777 ( .A1(n716), .A2(n718), .ZN(n717) );
  XNOR2_X1 U778 ( .A(n717), .B(G146), .ZN(G48) );
  XOR2_X1 U779 ( .A(G113), .B(KEYINPUT113), .Z(n720) );
  NAND2_X1 U780 ( .A1(n722), .A2(n718), .ZN(n719) );
  XNOR2_X1 U781 ( .A(n720), .B(n719), .ZN(G15) );
  NAND2_X1 U782 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U783 ( .A(n723), .B(KEYINPUT114), .ZN(n724) );
  XNOR2_X1 U784 ( .A(G116), .B(n724), .ZN(G18) );
  NAND2_X1 U785 ( .A1(n356), .A2(n725), .ZN(n726) );
  XOR2_X1 U786 ( .A(KEYINPUT50), .B(n726), .Z(n734) );
  NAND2_X1 U787 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U788 ( .A(n729), .B(KEYINPUT49), .ZN(n730) );
  XNOR2_X1 U789 ( .A(KEYINPUT117), .B(n730), .ZN(n732) );
  NAND2_X1 U790 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U791 ( .A1(n734), .A2(n733), .ZN(n735) );
  XOR2_X1 U792 ( .A(KEYINPUT118), .B(n735), .Z(n737) );
  NAND2_X1 U793 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U794 ( .A(n738), .B(KEYINPUT51), .ZN(n739) );
  NOR2_X1 U795 ( .A1(n739), .A2(n769), .ZN(n755) );
  INV_X1 U796 ( .A(n740), .ZN(n770) );
  NOR2_X1 U797 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U798 ( .A1(n744), .A2(n743), .ZN(n751) );
  NOR2_X1 U799 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U800 ( .A(n747), .B(KEYINPUT119), .ZN(n749) );
  NAND2_X1 U801 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U802 ( .A1(n751), .A2(n750), .ZN(n752) );
  XOR2_X1 U803 ( .A(KEYINPUT120), .B(n752), .Z(n753) );
  NOR2_X1 U804 ( .A1(n770), .A2(n753), .ZN(n754) );
  NOR2_X1 U805 ( .A1(n755), .A2(n754), .ZN(n756) );
  XOR2_X1 U806 ( .A(KEYINPUT52), .B(n756), .Z(n757) );
  NAND2_X1 U807 ( .A1(n758), .A2(n757), .ZN(n768) );
  NAND2_X1 U808 ( .A1(n647), .A2(n763), .ZN(n759) );
  XOR2_X1 U809 ( .A(KEYINPUT82), .B(n759), .Z(n762) );
  NAND2_X1 U810 ( .A1(n400), .A2(KEYINPUT2), .ZN(n760) );
  NOR2_X1 U811 ( .A1(n764), .A2(n760), .ZN(n761) );
  NOR2_X1 U812 ( .A1(n762), .A2(n761), .ZN(n767) );
  NAND2_X1 U813 ( .A1(n764), .A2(n763), .ZN(n765) );
  XOR2_X1 U814 ( .A(KEYINPUT81), .B(n765), .Z(n766) );
  XNOR2_X1 U815 ( .A(n772), .B(KEYINPUT94), .ZN(n773) );
  XNOR2_X1 U816 ( .A(n771), .B(n773), .ZN(n776) );
  XNOR2_X1 U817 ( .A(n647), .B(n776), .ZN(n775) );
  NAND2_X1 U818 ( .A1(n775), .A2(n774), .ZN(n780) );
  XNOR2_X1 U819 ( .A(G227), .B(n776), .ZN(n777) );
  NAND2_X1 U820 ( .A1(n777), .A2(G900), .ZN(n778) );
  NAND2_X1 U821 ( .A1(G953), .A2(n778), .ZN(n779) );
  NAND2_X1 U822 ( .A1(n780), .A2(n779), .ZN(G72) );
  XOR2_X1 U823 ( .A(G143), .B(n781), .Z(n782) );
  XNOR2_X1 U824 ( .A(KEYINPUT112), .B(n782), .ZN(G45) );
endmodule

