//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 0 0 0 1 0 0 0 0 1 0 1 1 1 0 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 1 1 1 1 1 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:09 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n558,
    new_n559, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n623, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1203;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT66), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n454), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n461), .A2(G101), .A3(G2104), .ZN(new_n462));
  XOR2_X1   g037(.A(new_n462), .B(KEYINPUT71), .Z(new_n463));
  INV_X1    g038(.A(KEYINPUT69), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  OAI211_X1 g040(.A(new_n464), .B(KEYINPUT3), .C1(new_n465), .C2(KEYINPUT70), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  OAI21_X1  g042(.A(KEYINPUT69), .B1(new_n467), .B2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT70), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n469), .A2(new_n467), .A3(G2104), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n466), .A2(new_n468), .A3(new_n470), .A4(new_n461), .ZN(new_n471));
  INV_X1    g046(.A(G137), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n463), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n467), .A2(G2104), .ZN(new_n475));
  AND3_X1   g050(.A1(new_n474), .A2(new_n475), .A3(KEYINPUT67), .ZN(new_n476));
  AOI21_X1  g051(.A(KEYINPUT67), .B1(new_n474), .B2(new_n475), .ZN(new_n477));
  OAI21_X1  g052(.A(G125), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(KEYINPUT68), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT67), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n467), .A2(G2104), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n474), .A2(new_n475), .A3(KEYINPUT67), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT68), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n485), .A2(new_n486), .A3(G125), .ZN(new_n487));
  NAND2_X1  g062(.A1(G113), .A2(G2104), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n479), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n473), .B1(new_n489), .B2(G2105), .ZN(G160));
  INV_X1    g065(.A(new_n471), .ZN(new_n491));
  AND2_X1   g066(.A1(new_n491), .A2(G136), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G112), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n493), .B1(new_n494), .B2(G2105), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n466), .A2(new_n468), .A3(new_n470), .A4(G2105), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT72), .ZN(new_n497));
  OR2_X1    g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n497), .ZN(new_n499));
  AND2_X1   g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI211_X1 g075(.A(new_n492), .B(new_n495), .C1(new_n500), .C2(G124), .ZN(G162));
  OR2_X1    g076(.A1(G102), .A2(G2105), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n502), .B(G2104), .C1(G114), .C2(new_n461), .ZN(new_n503));
  INV_X1    g078(.A(G126), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n503), .B1(new_n496), .B2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G138), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n506), .A2(G2105), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n466), .A2(new_n468), .A3(new_n470), .A4(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT4), .ZN(new_n509));
  NOR3_X1   g084(.A1(new_n506), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n510), .B1(new_n476), .B2(new_n477), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n505), .B1(new_n509), .B2(new_n511), .ZN(G164));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n517), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n517), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n521));
  OR2_X1    g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n521), .A2(new_n525), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n520), .A2(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  NAND3_X1  g103(.A1(new_n517), .A2(G63), .A3(G651), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(G89), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n524), .A2(new_n517), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT73), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n524), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n522), .A2(KEYINPUT73), .A3(new_n523), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n537), .A2(G543), .A3(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(G51), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n535), .A2(new_n541), .ZN(G168));
  AND3_X1   g117(.A1(new_n537), .A2(G543), .A3(new_n538), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G52), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(new_n519), .ZN(new_n546));
  INV_X1    g121(.A(new_n534), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G90), .ZN(new_n548));
  AND3_X1   g123(.A1(new_n544), .A2(new_n546), .A3(new_n548), .ZN(G171));
  NAND2_X1  g124(.A1(new_n543), .A2(G43), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n517), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n551), .A2(new_n519), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n547), .A2(G81), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n550), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  INV_X1    g136(.A(new_n517), .ZN(new_n562));
  INV_X1    g137(.A(G65), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G651), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n547), .A2(G91), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT9), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n543), .A2(new_n568), .A3(G53), .ZN(new_n569));
  INV_X1    g144(.A(G53), .ZN(new_n570));
  OAI21_X1  g145(.A(KEYINPUT9), .B1(new_n539), .B2(new_n570), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n567), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(G299));
  NAND3_X1  g148(.A1(new_n544), .A2(new_n546), .A3(new_n548), .ZN(G301));
  NAND2_X1  g149(.A1(G168), .A2(KEYINPUT74), .ZN(new_n575));
  OAI221_X1 g150(.A(new_n532), .B1(new_n533), .B2(new_n534), .C1(new_n540), .C2(new_n539), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT74), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(G286));
  OAI21_X1  g155(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n524), .A2(new_n517), .A3(G87), .ZN(new_n582));
  AND2_X1   g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n537), .A2(G49), .A3(G543), .A4(new_n538), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(KEYINPUT75), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT75), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n583), .A2(new_n587), .A3(new_n584), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G288));
  INV_X1    g165(.A(G61), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n591), .B1(new_n515), .B2(new_n516), .ZN(new_n592));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(G651), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n524), .A2(G48), .A3(G543), .ZN(new_n596));
  AND2_X1   g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n524), .A2(new_n517), .A3(G86), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(G305));
  NAND2_X1  g174(.A1(new_n547), .A2(G85), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G47), .ZN(new_n602));
  OAI221_X1 g177(.A(new_n600), .B1(new_n519), .B2(new_n601), .C1(new_n602), .C2(new_n539), .ZN(G290));
  NAND2_X1  g178(.A1(G301), .A2(G868), .ZN(new_n604));
  INV_X1    g179(.A(G54), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n605), .B1(new_n539), .B2(KEYINPUT76), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(KEYINPUT76), .B2(new_n539), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n547), .A2(KEYINPUT10), .A3(G92), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT10), .ZN(new_n609));
  INV_X1    g184(.A(G92), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n534), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(G79), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(G66), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n562), .B2(new_n613), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n608), .A2(new_n611), .B1(G651), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n607), .A2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n604), .B1(new_n617), .B2(G868), .ZN(G284));
  OAI21_X1  g193(.A(new_n604), .B1(new_n617), .B2(G868), .ZN(G321));
  NOR2_X1   g194(.A1(G299), .A2(G868), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n620), .B1(G868), .B2(new_n579), .ZN(G297));
  XNOR2_X1  g196(.A(G297), .B(KEYINPUT77), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n617), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n617), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G868), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G868), .B2(new_n555), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g203(.A1(new_n465), .A2(G2105), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n485), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT12), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT13), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(G2100), .Z(new_n633));
  NAND2_X1  g208(.A1(new_n500), .A2(G123), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n491), .A2(G135), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n461), .A2(G111), .ZN(new_n636));
  OAI21_X1  g211(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n637));
  OAI211_X1 g212(.A(new_n634), .B(new_n635), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(G2096), .Z(new_n639));
  NAND2_X1  g214(.A1(new_n633), .A2(new_n639), .ZN(G156));
  INV_X1    g215(.A(KEYINPUT14), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2427), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2430), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n641), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n645), .B1(new_n644), .B2(new_n643), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2451), .B(G2454), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT16), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n646), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(G14), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n651), .A2(new_n652), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(G401));
  XNOR2_X1  g231(.A(G2072), .B(G2078), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT17), .Z(new_n658));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2084), .B(G2090), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT78), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n663), .B1(new_n659), .B2(new_n657), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT80), .Z(new_n666));
  INV_X1    g241(.A(new_n663), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n667), .A2(new_n658), .A3(new_n660), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT81), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n667), .A2(new_n659), .A3(new_n657), .ZN(new_n670));
  XOR2_X1   g245(.A(KEYINPUT79), .B(KEYINPUT18), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n666), .A2(new_n669), .A3(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G2096), .B(G2100), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT82), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n673), .B(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(G227));
  XOR2_X1   g252(.A(G1971), .B(G1976), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT19), .ZN(new_n679));
  XOR2_X1   g254(.A(G1956), .B(G2474), .Z(new_n680));
  XOR2_X1   g255(.A(G1961), .B(G1966), .Z(new_n681));
  AND2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT20), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n680), .A2(new_n681), .ZN(new_n685));
  NOR3_X1   g260(.A1(new_n679), .A2(new_n682), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(new_n679), .B2(new_n685), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT83), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n688), .B(new_n690), .Z(new_n691));
  XOR2_X1   g266(.A(G1991), .B(G1996), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1981), .B(G1986), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n691), .A2(new_n692), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n691), .A2(new_n692), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n697), .A2(new_n694), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n696), .A2(new_n699), .ZN(G229));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NOR2_X1   g276(.A1(G168), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(new_n701), .B2(G21), .ZN(new_n703));
  INV_X1    g278(.A(G1966), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT89), .Z(new_n706));
  NOR2_X1   g281(.A1(G171), .A2(new_n701), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G5), .B2(new_n701), .ZN(new_n708));
  INV_X1    g283(.A(G1961), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(G29), .ZN(new_n711));
  OAI221_X1 g286(.A(new_n710), .B1(new_n711), .B2(new_n638), .C1(new_n703), .C2(new_n704), .ZN(new_n712));
  INV_X1    g287(.A(G28), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n713), .A2(KEYINPUT30), .ZN(new_n714));
  AOI21_X1  g289(.A(G29), .B1(new_n713), .B2(KEYINPUT30), .ZN(new_n715));
  OR2_X1    g290(.A1(KEYINPUT31), .A2(G11), .ZN(new_n716));
  NAND2_X1  g291(.A1(KEYINPUT31), .A2(G11), .ZN(new_n717));
  AOI22_X1  g292(.A1(new_n714), .A2(new_n715), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n711), .A2(G33), .ZN(new_n719));
  AOI22_X1  g294(.A1(new_n485), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n720), .A2(new_n461), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT25), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n491), .B2(G139), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n719), .B1(new_n725), .B2(G29), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  OAI221_X1 g302(.A(new_n718), .B1(new_n727), .B2(G2072), .C1(new_n709), .C2(new_n708), .ZN(new_n728));
  NOR3_X1   g303(.A1(new_n706), .A2(new_n712), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n711), .A2(G27), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G164), .B2(new_n711), .ZN(new_n731));
  INV_X1    g306(.A(G2078), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(G2072), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n733), .B1(new_n726), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(G160), .A2(new_n711), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n711), .B1(KEYINPUT24), .B2(G34), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(KEYINPUT24), .B2(G34), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(G2084), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT27), .B(G1996), .Z(new_n742));
  NAND2_X1  g317(.A1(new_n500), .A2(G129), .ZN(new_n743));
  NAND3_X1  g318(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT86), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT26), .ZN(new_n746));
  AOI22_X1  g321(.A1(new_n491), .A2(G141), .B1(G105), .B2(new_n629), .ZN(new_n747));
  AND2_X1   g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n743), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n749), .A2(new_n711), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(KEYINPUT87), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT87), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G29), .B2(G32), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n751), .B1(new_n750), .B2(new_n753), .ZN(new_n754));
  AOI211_X1 g329(.A(new_n735), .B(new_n741), .C1(new_n742), .C2(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n754), .A2(new_n742), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT88), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n729), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT90), .Z(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT84), .B(G16), .ZN(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n761), .A2(G22), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(G166), .B2(new_n761), .ZN(new_n763));
  INV_X1    g338(.A(G1971), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  MUX2_X1   g340(.A(G23), .B(new_n585), .S(G16), .Z(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT33), .B(G1976), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n701), .A2(G6), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G305), .B2(G16), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT32), .B(G1981), .Z(new_n771));
  OR2_X1    g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n770), .A2(new_n771), .ZN(new_n773));
  NAND4_X1  g348(.A1(new_n765), .A2(new_n768), .A3(new_n772), .A4(new_n773), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n774), .A2(KEYINPUT34), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(KEYINPUT34), .ZN(new_n776));
  NOR2_X1   g351(.A1(G25), .A2(G29), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n500), .A2(G119), .ZN(new_n778));
  OAI21_X1  g353(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n779));
  INV_X1    g354(.A(G107), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n779), .B1(new_n780), .B2(G2105), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n491), .B2(G131), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n778), .A2(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n777), .B1(new_n784), .B2(G29), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT35), .B(G1991), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  MUX2_X1   g362(.A(G24), .B(G290), .S(new_n761), .Z(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(G1986), .Z(new_n789));
  NAND4_X1  g364(.A1(new_n775), .A2(new_n776), .A3(new_n787), .A4(new_n789), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT36), .Z(new_n791));
  NOR2_X1   g366(.A1(new_n761), .A2(G19), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n555), .B2(new_n761), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G1341), .ZN(new_n794));
  INV_X1    g369(.A(G1348), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n617), .A2(G16), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G4), .B2(G16), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n794), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n797), .A2(new_n795), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n711), .A2(G26), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT28), .Z(new_n801));
  NAND2_X1  g376(.A1(new_n500), .A2(G128), .ZN(new_n802));
  OAI21_X1  g377(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n803));
  INV_X1    g378(.A(G116), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n803), .B1(new_n804), .B2(G2105), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n491), .B2(G140), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n802), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n801), .B1(new_n807), .B2(G29), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT85), .B(G2067), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n760), .A2(G20), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT23), .Z(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(G299), .B2(G16), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(G1956), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n798), .A2(new_n799), .A3(new_n810), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n711), .A2(G35), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G162), .B2(new_n711), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT91), .B(KEYINPUT29), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT92), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n817), .B(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(G2090), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NOR4_X1   g397(.A1(new_n759), .A2(new_n791), .A3(new_n815), .A4(new_n822), .ZN(G311));
  INV_X1    g398(.A(G311), .ZN(G150));
  XOR2_X1   g399(.A(KEYINPUT93), .B(G55), .Z(new_n825));
  NAND2_X1  g400(.A1(new_n543), .A2(new_n825), .ZN(new_n826));
  AOI22_X1  g401(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n827), .A2(new_n519), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n547), .A2(G93), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n826), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(KEYINPUT94), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT94), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n826), .A2(new_n832), .A3(new_n828), .A4(new_n829), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(G860), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT37), .Z(new_n836));
  NAND2_X1  g411(.A1(new_n617), .A2(G559), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT38), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n831), .A2(new_n554), .A3(new_n833), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n555), .A2(new_n830), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n838), .B(new_n841), .Z(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  AND2_X1   g418(.A1(new_n843), .A2(KEYINPUT39), .ZN(new_n844));
  INV_X1    g419(.A(G860), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(new_n843), .B2(KEYINPUT39), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n836), .B1(new_n844), .B2(new_n846), .ZN(G145));
  NAND2_X1  g422(.A1(new_n725), .A2(KEYINPUT96), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n749), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(new_n807), .ZN(new_n851));
  INV_X1    g426(.A(new_n807), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(new_n749), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n511), .A2(new_n509), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n496), .A2(new_n504), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n854), .A2(new_n855), .A3(new_n503), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT95), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n851), .A2(new_n853), .A3(new_n857), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n725), .A2(KEYINPUT96), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n857), .B1(new_n851), .B2(new_n853), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n849), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n861), .ZN(new_n863));
  NAND4_X1  g438(.A1(new_n863), .A2(new_n848), .A3(new_n859), .A4(new_n858), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n783), .B(new_n631), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n500), .A2(G130), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT97), .ZN(new_n867));
  OAI21_X1  g442(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n868));
  INV_X1    g443(.A(G118), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n868), .B1(new_n869), .B2(G2105), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n870), .B1(new_n491), .B2(G142), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n867), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n865), .B(new_n872), .ZN(new_n873));
  AND3_X1   g448(.A1(new_n862), .A2(new_n864), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n873), .B1(new_n862), .B2(new_n864), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n638), .B(G160), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(G162), .ZN(new_n878));
  AOI21_X1  g453(.A(G37), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT98), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n862), .A2(new_n864), .ZN(new_n881));
  INV_X1    g456(.A(new_n873), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n862), .A2(new_n864), .A3(new_n873), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n878), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n880), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  OAI211_X1 g462(.A(new_n880), .B(new_n886), .C1(new_n874), .C2(new_n875), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n879), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g466(.A(G290), .B(G305), .Z(new_n892));
  XOR2_X1   g467(.A(G303), .B(new_n585), .Z(new_n893));
  XNOR2_X1  g468(.A(new_n892), .B(new_n893), .ZN(new_n894));
  OR2_X1    g469(.A1(new_n894), .A2(KEYINPUT101), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(KEYINPUT42), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n841), .B(new_n625), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n616), .A2(new_n572), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(KEYINPUT99), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n617), .A2(G299), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT99), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n616), .A2(new_n572), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n900), .A2(new_n901), .A3(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n898), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT100), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n906), .B(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT41), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n904), .A2(KEYINPUT41), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n910), .A2(new_n898), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n897), .B(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(G868), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT102), .ZN(new_n916));
  INV_X1    g491(.A(new_n834), .ZN(new_n917));
  OAI211_X1 g492(.A(new_n915), .B(new_n916), .C1(G868), .C2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n913), .B(new_n896), .ZN(new_n919));
  INV_X1    g494(.A(G868), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n917), .A2(G868), .ZN(new_n922));
  OAI21_X1  g497(.A(KEYINPUT102), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n918), .A2(new_n923), .ZN(G295));
  INV_X1    g499(.A(KEYINPUT103), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n915), .B(new_n925), .C1(G868), .C2(new_n917), .ZN(new_n926));
  OAI21_X1  g501(.A(KEYINPUT103), .B1(new_n921), .B2(new_n922), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(G331));
  NAND3_X1  g503(.A1(new_n575), .A2(G171), .A3(new_n578), .ZN(new_n929));
  NAND3_X1  g504(.A1(G168), .A2(KEYINPUT104), .A3(G301), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT104), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n931), .B1(G171), .B2(new_n576), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n929), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(new_n841), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT105), .B1(new_n933), .B2(new_n841), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n932), .A2(new_n930), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n938), .A2(new_n840), .A3(new_n839), .A4(new_n929), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n934), .B1(new_n939), .B2(KEYINPUT105), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n904), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n933), .A2(new_n841), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n910), .B(new_n911), .C1(new_n942), .C2(new_n935), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n941), .A2(new_n894), .A3(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(G37), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n894), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n910), .A2(new_n911), .ZN(new_n948));
  NOR3_X1   g523(.A1(new_n948), .A2(new_n937), .A3(new_n940), .ZN(new_n949));
  NOR3_X1   g524(.A1(new_n935), .A2(new_n942), .A3(new_n905), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n947), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  AND3_X1   g526(.A1(new_n946), .A2(KEYINPUT43), .A3(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n935), .A2(new_n942), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n948), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n935), .A2(new_n936), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n939), .A2(KEYINPUT105), .A3(new_n934), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n905), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n947), .B1(new_n954), .B2(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n958), .A2(new_n944), .A3(new_n945), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT43), .ZN(new_n960));
  AND2_X1   g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT44), .B1(new_n952), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n951), .A2(new_n960), .A3(new_n945), .A4(new_n944), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n963), .A2(KEYINPUT106), .A3(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT106), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n946), .A2(new_n966), .A3(new_n960), .A4(new_n951), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n962), .B1(new_n968), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g544(.A(G2067), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n807), .B(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G1996), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n749), .B(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n783), .B(new_n786), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n971), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  XNOR2_X1  g550(.A(G290), .B(G1986), .ZN(new_n976));
  OR2_X1    g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n463), .B(G40), .C1(new_n472), .C2(new_n471), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n978), .B1(new_n489), .B2(G2105), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT45), .ZN(new_n981));
  XOR2_X1   g556(.A(KEYINPUT107), .B(G1384), .Z(new_n982));
  OAI21_X1  g557(.A(new_n981), .B1(G164), .B2(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n977), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(G303), .A2(G8), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT55), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n982), .ZN(new_n992));
  AOI22_X1  g567(.A1(new_n485), .A2(new_n510), .B1(KEYINPUT4), .B2(new_n508), .ZN(new_n993));
  OAI211_X1 g568(.A(KEYINPUT45), .B(new_n992), .C1(new_n993), .C2(new_n505), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT108), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n856), .A2(KEYINPUT108), .A3(KEYINPUT45), .A4(new_n992), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n981), .B1(G164), .B2(G1384), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n979), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n764), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT50), .ZN(new_n1002));
  INV_X1    g577(.A(G1384), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n856), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n979), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT109), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1006), .A2(new_n1007), .A3(new_n821), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n979), .A2(new_n1005), .A3(new_n1004), .A4(new_n821), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(KEYINPUT109), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1001), .A2(new_n1008), .A3(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n991), .B1(new_n1011), .B2(G8), .ZN(new_n1012));
  INV_X1    g587(.A(G8), .ZN(new_n1013));
  NOR2_X1   g588(.A1(G164), .A2(G1384), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1013), .B1(new_n979), .B2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n583), .A2(G1976), .A3(new_n584), .ZN(new_n1016));
  XOR2_X1   g591(.A(new_n1016), .B(KEYINPUT111), .Z(new_n1017));
  NAND2_X1  g592(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT52), .ZN(new_n1019));
  INV_X1    g594(.A(G1976), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT52), .B1(G288), .B2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1021), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1022));
  INV_X1    g597(.A(G1981), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n595), .A2(new_n1023), .A3(new_n598), .A4(new_n596), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT112), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n1024), .B(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g601(.A(KEYINPUT113), .B(G86), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n597), .B1(new_n534), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(G1981), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT49), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1026), .A2(new_n1029), .A3(KEYINPUT49), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1032), .A2(new_n1015), .A3(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1019), .A2(new_n1022), .A3(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(KEYINPUT115), .B1(new_n1012), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT115), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n1019), .A2(new_n1022), .A3(new_n1034), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n996), .A2(new_n997), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1039), .A2(new_n979), .A3(new_n999), .ZN(new_n1040));
  AOI22_X1  g615(.A1(new_n1040), .A2(new_n764), .B1(KEYINPUT109), .B2(new_n1009), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1013), .B1(new_n1041), .B2(new_n1008), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1037), .B(new_n1038), .C1(new_n1042), .C2(new_n991), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n856), .A2(KEYINPUT45), .A3(new_n1003), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n979), .A2(new_n999), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(new_n704), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n979), .A2(new_n1005), .A3(new_n1004), .A4(new_n740), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1013), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1048), .A2(KEYINPUT63), .A3(new_n579), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT110), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n991), .B(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1049), .B1(new_n1042), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1036), .A2(new_n1043), .A3(new_n1052), .ZN(new_n1053));
  AOI22_X1  g628(.A1(new_n1040), .A2(new_n764), .B1(new_n821), .B2(new_n1006), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n989), .B(new_n990), .C1(new_n1054), .C2(new_n1013), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1011), .A2(new_n1051), .A3(G8), .ZN(new_n1056));
  AOI22_X1  g631(.A1(new_n1006), .A2(new_n740), .B1(new_n1045), .B2(new_n704), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n1057), .A2(new_n1013), .A3(G286), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1055), .A2(new_n1056), .A3(new_n1038), .A4(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT63), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1053), .A2(new_n1061), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1056), .A2(new_n1035), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n589), .A2(new_n1020), .ZN(new_n1064));
  XOR2_X1   g639(.A(new_n1064), .B(KEYINPUT114), .Z(new_n1065));
  AND2_X1   g640(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1026), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1063), .B1(new_n1015), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1062), .A2(new_n1068), .ZN(new_n1069));
  AND2_X1   g644(.A1(new_n979), .A2(new_n999), .ZN(new_n1070));
  XNOR2_X1  g645(.A(KEYINPUT56), .B(G2072), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1070), .A2(new_n1039), .A3(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g647(.A(new_n572), .B(KEYINPUT57), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n979), .A2(new_n1005), .A3(new_n1004), .ZN(new_n1074));
  INV_X1    g649(.A(G1956), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1072), .A2(new_n1073), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1073), .B1(new_n1072), .B2(new_n1076), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1074), .A2(new_n795), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n979), .A2(new_n970), .A3(new_n1014), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n616), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1077), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1077), .ZN(new_n1083));
  OAI21_X1  g658(.A(KEYINPUT61), .B1(new_n1083), .B2(new_n1078), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1078), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT61), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1085), .A2(new_n1086), .A3(new_n1077), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1084), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT117), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n554), .B1(new_n1089), .B2(KEYINPUT59), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1070), .A2(new_n972), .A3(new_n1039), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT116), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n979), .A2(new_n1014), .ZN(new_n1093));
  XOR2_X1   g668(.A(KEYINPUT58), .B(G1341), .Z(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1091), .A2(new_n1092), .A3(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1092), .B1(new_n1091), .B2(new_n1095), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1090), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT59), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1098), .A2(KEYINPUT117), .A3(new_n1099), .ZN(new_n1100));
  OAI221_X1 g675(.A(new_n1090), .B1(new_n1089), .B2(KEYINPUT59), .C1(new_n1096), .C2(new_n1097), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1088), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT60), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT118), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(new_n617), .ZN(new_n1106));
  OAI211_X1 g681(.A(KEYINPUT118), .B(new_n616), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  OR3_X1    g683(.A1(new_n1103), .A2(KEYINPUT118), .A3(new_n1104), .ZN(new_n1109));
  AOI22_X1  g684(.A1(new_n1108), .A2(new_n1109), .B1(new_n1104), .B2(new_n1103), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1082), .B1(new_n1102), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT53), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1112), .A2(G2078), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n979), .A2(new_n983), .A3(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(KEYINPUT121), .B1(new_n998), .B2(new_n1114), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n979), .A2(new_n1113), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT121), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1116), .A2(new_n1117), .A3(new_n983), .A4(new_n1039), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1074), .A2(new_n709), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1115), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1070), .A2(new_n732), .A3(new_n1039), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(new_n1112), .ZN(new_n1122));
  AOI21_X1  g697(.A(G301), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n979), .A2(new_n999), .A3(new_n1044), .ZN(new_n1124));
  AOI22_X1  g699(.A1(new_n1124), .A2(new_n1113), .B1(new_n1074), .B2(new_n709), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1122), .A2(G301), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(KEYINPUT54), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n1128));
  NOR3_X1   g703(.A1(new_n1123), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  AND2_X1   g704(.A1(new_n1126), .A2(KEYINPUT54), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1122), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1115), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1132));
  OAI21_X1  g707(.A(G171), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(KEYINPUT122), .B1(new_n1130), .B2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1129), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT54), .ZN(new_n1136));
  NOR3_X1   g711(.A1(new_n1131), .A2(new_n1132), .A3(G171), .ZN(new_n1137));
  AOI21_X1  g712(.A(G301), .B1(new_n1122), .B2(new_n1125), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1136), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT120), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n576), .A2(G8), .ZN(new_n1141));
  XNOR2_X1  g716(.A(new_n1141), .B(KEYINPUT119), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1140), .B1(new_n1048), .B2(new_n1143), .ZN(new_n1144));
  OAI211_X1 g719(.A(KEYINPUT120), .B(new_n1142), .C1(new_n1057), .C2(new_n1013), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1144), .A2(new_n1145), .A3(KEYINPUT51), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT51), .ZN(new_n1147));
  OAI211_X1 g722(.A(new_n1140), .B(new_n1147), .C1(new_n1048), .C2(new_n1143), .ZN(new_n1148));
  OR2_X1    g723(.A1(new_n1057), .A2(new_n1142), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1146), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  AND3_X1   g725(.A1(new_n1055), .A2(new_n1056), .A3(new_n1038), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1139), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1135), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1069), .B1(new_n1111), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT123), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1150), .A2(KEYINPUT62), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT62), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1146), .A2(new_n1157), .A3(new_n1148), .A4(new_n1149), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1055), .A2(new_n1056), .A3(new_n1138), .A4(new_n1038), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1159), .ZN(new_n1160));
  AND4_X1   g735(.A1(new_n1155), .A2(new_n1156), .A3(new_n1158), .A4(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1159), .B1(new_n1150), .B2(KEYINPUT62), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1155), .B1(new_n1162), .B2(new_n1158), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n986), .B1(new_n1154), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n984), .A2(new_n972), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n1166), .B(KEYINPUT46), .ZN(new_n1167));
  AND2_X1   g742(.A1(new_n971), .A2(new_n850), .ZN(new_n1168));
  INV_X1    g743(.A(new_n984), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1167), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n1170), .B(KEYINPUT47), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n973), .A2(new_n971), .A3(new_n784), .A4(new_n786), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n852), .A2(new_n970), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1169), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NOR3_X1   g749(.A1(new_n1169), .A2(G1986), .A3(G290), .ZN(new_n1175));
  XOR2_X1   g750(.A(new_n1175), .B(KEYINPUT48), .Z(new_n1176));
  NAND2_X1  g751(.A1(new_n975), .A2(new_n984), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1174), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1171), .A2(new_n1178), .ZN(new_n1179));
  XOR2_X1   g754(.A(new_n1179), .B(KEYINPUT124), .Z(new_n1180));
  OAI21_X1  g755(.A(KEYINPUT125), .B1(new_n1165), .B2(new_n1180), .ZN(new_n1181));
  OR2_X1    g756(.A1(new_n1129), .A2(new_n1134), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1152), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1111), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1162), .A2(new_n1158), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1185), .A2(KEYINPUT123), .ZN(new_n1186));
  AND2_X1   g761(.A1(new_n1062), .A2(new_n1068), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1162), .A2(new_n1155), .A3(new_n1158), .ZN(new_n1188));
  NAND4_X1  g763(.A1(new_n1184), .A2(new_n1186), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1189), .A2(new_n985), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT125), .ZN(new_n1191));
  XNOR2_X1  g766(.A(new_n1179), .B(KEYINPUT124), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1181), .A2(new_n1193), .ZN(G329));
  assign    G231 = 1'b0;
  OAI211_X1 g769(.A(new_n676), .B(G319), .C1(new_n655), .C2(new_n654), .ZN(new_n1196));
  OAI21_X1  g770(.A(KEYINPUT126), .B1(G229), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g771(.A(new_n1196), .ZN(new_n1198));
  INV_X1    g772(.A(KEYINPUT126), .ZN(new_n1199));
  NAND4_X1  g773(.A1(new_n1198), .A2(new_n1199), .A3(new_n699), .A4(new_n696), .ZN(new_n1200));
  NAND2_X1  g774(.A1(new_n1197), .A2(new_n1200), .ZN(new_n1201));
  NAND4_X1  g775(.A1(new_n965), .A2(new_n890), .A3(new_n967), .A4(new_n1201), .ZN(G225));
  INV_X1    g776(.A(KEYINPUT127), .ZN(new_n1203));
  XNOR2_X1  g777(.A(G225), .B(new_n1203), .ZN(G308));
endmodule


