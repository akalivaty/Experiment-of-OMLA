//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 0 0 1 0 1 1 0 0 1 1 0 1 0 0 1 0 1 1 0 1 1 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 1 1 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:48 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n446, new_n448, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n555, new_n557,
    new_n558, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n612, new_n613, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1196, new_n1197,
    new_n1198;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT66), .Z(G173));
  XNOR2_X1  g022(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n448));
  AND2_X1   g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  NAND2_X1  g025(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n449), .A2(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(G101), .A2(G2104), .ZN(new_n471));
  INV_X1    g046(.A(G137), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n471), .B1(new_n466), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n470), .A2(new_n475), .ZN(G160));
  NOR2_X1   g051(.A1(new_n466), .A2(new_n474), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n466), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  NOR2_X1   g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI21_X1  g056(.A(G2104), .B1(new_n474), .B2(G112), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n478), .B(new_n480), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT68), .ZN(G162));
  INV_X1    g059(.A(KEYINPUT70), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(new_n474), .B2(G114), .ZN(new_n486));
  NOR2_X1   g061(.A1(G102), .A2(G2105), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OR2_X1    g063(.A1(G102), .A2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n489), .A2(new_n491), .A3(KEYINPUT70), .A4(G2104), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g068(.A(KEYINPUT3), .B(G2104), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT69), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n494), .A2(new_n495), .A3(G126), .A4(G2105), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n463), .A2(new_n465), .A3(G126), .A4(G2105), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT69), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n493), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n463), .A2(new_n465), .A3(G138), .A4(new_n474), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n494), .A2(KEYINPUT4), .A3(G138), .A4(new_n474), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n499), .A2(new_n504), .ZN(G164));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  XOR2_X1   g081(.A(KEYINPUT71), .B(KEYINPUT5), .Z(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT72), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT72), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n507), .A2(new_n510), .A3(G543), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT5), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n512), .A2(G62), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(G75), .A2(G543), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n506), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AND2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n520), .A2(new_n513), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G50), .ZN(new_n522));
  INV_X1    g097(.A(new_n520), .ZN(new_n523));
  NAND4_X1  g098(.A1(new_n509), .A2(new_n514), .A3(new_n511), .A4(new_n523), .ZN(new_n524));
  XOR2_X1   g099(.A(KEYINPUT73), .B(G88), .Z(new_n525));
  OAI21_X1  g100(.A(new_n522), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n517), .A2(new_n526), .ZN(G166));
  INV_X1    g102(.A(KEYINPUT7), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n521), .A2(G51), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  XOR2_X1   g105(.A(KEYINPUT74), .B(G89), .Z(new_n531));
  OAI21_X1  g106(.A(new_n530), .B1(new_n524), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n512), .A2(new_n514), .ZN(new_n534));
  INV_X1    g109(.A(G63), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n532), .B1(new_n536), .B2(G651), .ZN(G168));
  AND2_X1   g112(.A1(new_n512), .A2(new_n514), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G64), .ZN(new_n539));
  NAND2_X1  g114(.A1(G77), .A2(G543), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n506), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n521), .A2(G52), .ZN(new_n542));
  INV_X1    g117(.A(G90), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n524), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n541), .A2(new_n544), .ZN(G171));
  NAND2_X1  g120(.A1(new_n521), .A2(G43), .ZN(new_n546));
  INV_X1    g121(.A(G81), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n524), .B2(new_n547), .ZN(new_n548));
  NAND4_X1  g123(.A1(new_n509), .A2(G56), .A3(new_n514), .A4(new_n511), .ZN(new_n549));
  NAND2_X1  g124(.A1(G68), .A2(G543), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n506), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  AND3_X1   g129(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G36), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n555), .A2(new_n558), .ZN(G188));
  NAND4_X1  g134(.A1(new_n509), .A2(G65), .A3(new_n514), .A4(new_n511), .ZN(new_n560));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n506), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n524), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n562), .B1(G91), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n521), .A2(G53), .ZN(new_n565));
  XOR2_X1   g140(.A(new_n565), .B(KEYINPUT9), .Z(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n564), .A2(new_n567), .ZN(G299));
  INV_X1    g143(.A(G171), .ZN(G301));
  INV_X1    g144(.A(G168), .ZN(G286));
  INV_X1    g145(.A(G166), .ZN(G303));
  INV_X1    g146(.A(G74), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n534), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G651), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n563), .A2(G87), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n521), .A2(G49), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(G288));
  NAND3_X1  g152(.A1(new_n512), .A2(G61), .A3(new_n514), .ZN(new_n578));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n506), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n512), .A2(G86), .A3(new_n514), .ZN(new_n582));
  NAND2_X1  g157(.A1(G48), .A2(G543), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(new_n523), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n581), .A2(new_n585), .ZN(G305));
  NAND2_X1  g161(.A1(new_n538), .A2(G60), .ZN(new_n587));
  NAND2_X1  g162(.A1(G72), .A2(G543), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n506), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(G85), .ZN(new_n590));
  INV_X1    g165(.A(new_n521), .ZN(new_n591));
  XNOR2_X1  g166(.A(KEYINPUT75), .B(G47), .ZN(new_n592));
  OAI22_X1  g167(.A1(new_n524), .A2(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n589), .A2(new_n593), .ZN(G290));
  NAND3_X1  g169(.A1(new_n512), .A2(G66), .A3(new_n514), .ZN(new_n595));
  NAND2_X1  g170(.A1(G79), .A2(G543), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n563), .A2(KEYINPUT10), .A3(G92), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT10), .ZN(new_n599));
  INV_X1    g174(.A(G92), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n524), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n597), .A2(G651), .B1(new_n598), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n521), .A2(G54), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(new_n605), .B2(G171), .ZN(G284));
  OAI21_X1  g182(.A(new_n606), .B1(new_n605), .B2(G171), .ZN(G321));
  NAND2_X1  g183(.A1(G299), .A2(new_n605), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(new_n605), .B2(G168), .ZN(G297));
  OAI21_X1  g185(.A(new_n609), .B1(new_n605), .B2(G168), .ZN(G280));
  INV_X1    g186(.A(new_n604), .ZN(new_n612));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(G860), .ZN(G148));
  NAND2_X1  g189(.A1(new_n552), .A2(new_n605), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n604), .A2(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(new_n605), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g193(.A1(new_n479), .A2(G2104), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2100), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n477), .A2(G123), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n479), .A2(G135), .ZN(new_n624));
  NOR2_X1   g199(.A1(G99), .A2(G2105), .ZN(new_n625));
  OAI21_X1  g200(.A(G2104), .B1(new_n474), .B2(G111), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n623), .B(new_n624), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(G2096), .Z(new_n628));
  NAND2_X1  g203(.A1(new_n622), .A2(new_n628), .ZN(G156));
  XOR2_X1   g204(.A(KEYINPUT15), .B(G2435), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2438), .ZN(new_n631));
  XOR2_X1   g206(.A(G2427), .B(G2430), .Z(new_n632));
  OAI21_X1  g207(.A(KEYINPUT14), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT76), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n631), .A2(new_n632), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  XOR2_X1   g212(.A(G2443), .B(G2446), .Z(new_n638));
  XNOR2_X1  g213(.A(G2451), .B(G2454), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n637), .B(new_n640), .Z(new_n641));
  XOR2_X1   g216(.A(G1341), .B(G1348), .Z(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  INV_X1    g219(.A(KEYINPUT77), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n641), .A2(new_n643), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n641), .A2(KEYINPUT77), .A3(new_n643), .ZN(new_n648));
  NAND4_X1  g223(.A1(new_n646), .A2(new_n647), .A3(G14), .A4(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(G401));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2067), .B(G2678), .Z(new_n653));
  NOR2_X1   g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n652), .A2(new_n653), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(new_n656), .A3(KEYINPUT17), .ZN(new_n657));
  INV_X1    g232(.A(KEYINPUT18), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2072), .B(G2078), .ZN(new_n660));
  OAI211_X1 g235(.A(new_n659), .B(new_n660), .C1(new_n658), .C2(new_n654), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n661), .B1(new_n660), .B2(new_n659), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2096), .B(G2100), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(G227));
  XNOR2_X1  g239(.A(G1971), .B(G1976), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT19), .ZN(new_n666));
  XOR2_X1   g241(.A(G1956), .B(G2474), .Z(new_n667));
  XOR2_X1   g242(.A(G1961), .B(G1966), .Z(new_n668));
  NAND3_X1  g243(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n669), .B1(new_n667), .B2(new_n668), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n666), .A2(KEYINPUT78), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n667), .A2(new_n668), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n666), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT20), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G1986), .B(G1996), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(G1981), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(G1991), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n678), .B(new_n681), .ZN(G229));
  XNOR2_X1  g257(.A(KEYINPUT80), .B(G16), .ZN(new_n683));
  MUX2_X1   g258(.A(G19), .B(new_n552), .S(new_n683), .Z(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(G1341), .Z(new_n685));
  NOR2_X1   g260(.A1(new_n589), .A2(new_n593), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(new_n683), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(G24), .B2(new_n683), .ZN(new_n688));
  INV_X1    g263(.A(G1986), .ZN(new_n689));
  AOI22_X1  g264(.A1(new_n688), .A2(new_n689), .B1(KEYINPUT81), .B2(KEYINPUT36), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(new_n689), .B2(new_n688), .ZN(new_n691));
  INV_X1    g266(.A(G16), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n692), .A2(G23), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n693), .B1(G288), .B2(G16), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT33), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n695), .A2(G1976), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(G1976), .ZN(new_n697));
  MUX2_X1   g272(.A(G6), .B(G305), .S(G16), .Z(new_n698));
  XOR2_X1   g273(.A(KEYINPUT32), .B(G1981), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  MUX2_X1   g275(.A(G22), .B(G303), .S(new_n683), .Z(new_n701));
  INV_X1    g276(.A(G1971), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND4_X1  g278(.A1(new_n696), .A2(new_n697), .A3(new_n700), .A4(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n691), .B1(new_n704), .B2(KEYINPUT34), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n477), .A2(G119), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT79), .Z(new_n707));
  NAND2_X1  g282(.A1(new_n479), .A2(G131), .ZN(new_n708));
  NOR2_X1   g283(.A1(G95), .A2(G2105), .ZN(new_n709));
  OAI21_X1  g284(.A(G2104), .B1(new_n474), .B2(G107), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n707), .B(new_n708), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  MUX2_X1   g286(.A(G25), .B(new_n711), .S(G29), .Z(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT35), .B(G1991), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n712), .B(new_n713), .Z(new_n714));
  OAI211_X1 g289(.A(new_n705), .B(new_n714), .C1(KEYINPUT34), .C2(new_n704), .ZN(new_n715));
  NOR2_X1   g290(.A1(KEYINPUT81), .A2(KEYINPUT36), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n715), .A2(new_n716), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT31), .B(G11), .ZN(new_n719));
  INV_X1    g294(.A(G28), .ZN(new_n720));
  AOI21_X1  g295(.A(G29), .B1(new_n720), .B2(KEYINPUT30), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(KEYINPUT30), .B2(new_n720), .ZN(new_n722));
  INV_X1    g297(.A(G29), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n722), .B1(new_n627), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(G5), .A2(G16), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(G171), .B2(G16), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n724), .B1(new_n726), .B2(G1961), .ZN(new_n727));
  NAND2_X1  g302(.A1(G168), .A2(G16), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n728), .A2(KEYINPUT84), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT84), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G16), .B2(G21), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n729), .B1(new_n728), .B2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(G1966), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n732), .A2(new_n733), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n719), .B(new_n727), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT85), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT88), .ZN(new_n739));
  INV_X1    g314(.A(G35), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n739), .B1(new_n740), .B2(G29), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n723), .A2(KEYINPUT88), .A3(G35), .ZN(new_n742));
  OAI211_X1 g317(.A(new_n741), .B(new_n742), .C1(G162), .C2(new_n723), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT29), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G2090), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT90), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(G20), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n683), .A2(new_n748), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT91), .B(KEYINPUT23), .Z(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G299), .B2(G16), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(G1956), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n747), .A2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT92), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n744), .A2(G2090), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT89), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n692), .A2(G4), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(new_n612), .B2(new_n692), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G1348), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n758), .A2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(G26), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n763), .A2(G29), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n479), .A2(G140), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT82), .Z(new_n766));
  OR2_X1    g341(.A1(G104), .A2(G2105), .ZN(new_n767));
  OAI211_X1 g342(.A(new_n767), .B(G2104), .C1(G116), .C2(new_n474), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n477), .A2(G128), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n766), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n764), .B1(new_n770), .B2(G29), .ZN(new_n771));
  MUX2_X1   g346(.A(new_n764), .B(new_n771), .S(KEYINPUT28), .Z(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G2067), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n723), .A2(G33), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n494), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n775), .A2(new_n474), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G139), .B2(new_n479), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT83), .B(KEYINPUT25), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n474), .A2(G103), .A3(G2104), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  AND2_X1   g356(.A1(new_n777), .A2(new_n781), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n774), .B1(new_n782), .B2(new_n723), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n783), .A2(G2072), .ZN(new_n784));
  OR2_X1    g359(.A1(KEYINPUT24), .A2(G34), .ZN(new_n785));
  NAND2_X1  g360(.A1(KEYINPUT24), .A2(G34), .ZN(new_n786));
  AND3_X1   g361(.A1(new_n785), .A2(new_n723), .A3(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(new_n475), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n788), .A2(new_n469), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n787), .B1(new_n789), .B2(G29), .ZN(new_n790));
  INV_X1    g365(.A(G2084), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n792), .A2(KEYINPUT86), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n477), .A2(G129), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n479), .A2(G141), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n474), .A2(G105), .A3(G2104), .ZN(new_n796));
  NAND3_X1  g371(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT26), .Z(new_n798));
  NAND4_X1  g373(.A1(new_n794), .A2(new_n795), .A3(new_n796), .A4(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n800), .A2(G29), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G29), .B2(G32), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT27), .B(G1996), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n793), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n802), .A2(new_n803), .ZN(new_n805));
  OAI221_X1 g380(.A(new_n805), .B1(new_n791), .B2(new_n790), .C1(new_n783), .C2(G2072), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n792), .A2(KEYINPUT86), .ZN(new_n807));
  NOR3_X1   g382(.A1(new_n804), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n773), .A2(new_n784), .A3(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n726), .A2(G1961), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n723), .A2(G27), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(G164), .B2(new_n723), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT87), .ZN(new_n813));
  INV_X1    g388(.A(G2078), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NOR3_X1   g390(.A1(new_n809), .A2(new_n810), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n756), .A2(new_n762), .A3(new_n816), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n754), .A2(new_n755), .ZN(new_n818));
  NOR3_X1   g393(.A1(new_n738), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  AND4_X1   g394(.A1(new_n685), .A2(new_n717), .A3(new_n718), .A4(new_n819), .ZN(G311));
  NAND4_X1  g395(.A1(new_n717), .A2(new_n819), .A3(new_n685), .A4(new_n718), .ZN(G150));
  INV_X1    g396(.A(G93), .ZN(new_n822));
  INV_X1    g397(.A(G55), .ZN(new_n823));
  OAI22_X1  g398(.A1(new_n524), .A2(new_n822), .B1(new_n823), .B2(new_n591), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT93), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI221_X1 g401(.A(KEYINPUT93), .B1(new_n823), .B2(new_n591), .C1(new_n524), .C2(new_n822), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(G80), .A2(G543), .ZN(new_n829));
  INV_X1    g404(.A(G67), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n829), .B1(new_n534), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(G651), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n828), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(G860), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT37), .Z(new_n835));
  NAND2_X1  g410(.A1(new_n612), .A2(G559), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT38), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n833), .A2(new_n553), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n828), .A2(new_n832), .A3(new_n552), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT39), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n837), .B(new_n841), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n835), .B1(new_n842), .B2(G860), .ZN(G145));
  XNOR2_X1  g418(.A(new_n711), .B(new_n620), .ZN(new_n844));
  INV_X1    g419(.A(new_n479), .ZN(new_n845));
  INV_X1    g420(.A(G142), .ZN(new_n846));
  OR3_X1    g421(.A1(new_n845), .A2(KEYINPUT97), .A3(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(KEYINPUT97), .B1(new_n845), .B2(new_n846), .ZN(new_n848));
  OR2_X1    g423(.A1(G106), .A2(G2105), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n849), .B(G2104), .C1(G118), .C2(new_n474), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n477), .A2(G130), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n847), .A2(new_n848), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n844), .B(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT95), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n504), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n502), .A2(new_n503), .A3(KEYINPUT95), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n499), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(KEYINPUT96), .ZN(new_n858));
  AND3_X1   g433(.A1(new_n493), .A2(new_n496), .A3(new_n498), .ZN(new_n859));
  AND3_X1   g434(.A1(new_n502), .A2(new_n503), .A3(KEYINPUT95), .ZN(new_n860));
  AOI21_X1  g435(.A(KEYINPUT95), .B1(new_n502), .B2(new_n503), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT96), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n858), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(new_n770), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n866), .A2(new_n799), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n799), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n867), .A2(new_n782), .A3(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n782), .B1(new_n867), .B2(new_n868), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n853), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n871), .ZN(new_n873));
  INV_X1    g448(.A(new_n853), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n873), .A2(new_n874), .A3(new_n869), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n789), .B(KEYINPUT94), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(G162), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(new_n627), .ZN(new_n879));
  AOI21_X1  g454(.A(G37), .B1(new_n876), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n872), .A2(KEYINPUT98), .ZN(new_n881));
  INV_X1    g456(.A(new_n879), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT98), .ZN(new_n883));
  OAI211_X1 g458(.A(new_n883), .B(new_n853), .C1(new_n870), .C2(new_n871), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n881), .A2(new_n875), .A3(new_n882), .A4(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n880), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g462(.A(G305), .B(KEYINPUT100), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(G303), .ZN(new_n890));
  NAND2_X1  g465(.A1(G288), .A2(G166), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n890), .A2(G290), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(G290), .B1(new_n891), .B2(new_n890), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n888), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n890), .A2(new_n891), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(new_n686), .ZN(new_n896));
  XOR2_X1   g471(.A(G305), .B(KEYINPUT100), .Z(new_n897));
  NAND3_X1  g472(.A1(new_n890), .A2(G290), .A3(new_n891), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n894), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(KEYINPUT101), .B(KEYINPUT42), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(KEYINPUT101), .A2(KEYINPUT42), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n904), .B1(new_n894), .B2(new_n899), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n604), .A2(G299), .ZN(new_n906));
  AOI211_X1 g481(.A(new_n566), .B(new_n562), .C1(G91), .C2(new_n563), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n907), .A2(new_n603), .A3(new_n602), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n906), .A2(KEYINPUT99), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(KEYINPUT99), .B1(new_n906), .B2(new_n908), .ZN(new_n910));
  OR2_X1    g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n828), .A2(new_n832), .A3(new_n552), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n552), .B1(new_n828), .B2(new_n832), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n914), .A2(new_n616), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n914), .A2(new_n616), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n911), .A2(new_n917), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n906), .A2(KEYINPUT41), .A3(new_n908), .ZN(new_n919));
  AOI21_X1  g494(.A(KEYINPUT41), .B1(new_n906), .B2(new_n908), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n921), .B1(new_n915), .B2(new_n916), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT102), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n918), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n923), .B1(new_n918), .B2(new_n922), .ZN(new_n925));
  OAI22_X1  g500(.A1(new_n903), .A2(new_n905), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n918), .A2(new_n922), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(KEYINPUT102), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n905), .B1(new_n901), .B2(new_n902), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n918), .A2(new_n922), .A3(new_n923), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n926), .A2(new_n931), .A3(G868), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT103), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n833), .A2(new_n605), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n934), .B1(new_n936), .B2(new_n933), .ZN(G295));
  OAI21_X1  g512(.A(new_n934), .B1(new_n936), .B2(new_n933), .ZN(G331));
  XOR2_X1   g513(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n939));
  OAI21_X1  g514(.A(G168), .B1(new_n912), .B2(new_n913), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n838), .A2(G286), .A3(new_n839), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n940), .A2(new_n941), .A3(G171), .ZN(new_n942));
  AOI21_X1  g517(.A(G171), .B1(new_n940), .B2(new_n941), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n921), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n940), .A2(new_n941), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(G301), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n907), .B1(new_n603), .B2(new_n602), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n604), .A2(G299), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n940), .A2(new_n941), .A3(G171), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n946), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n944), .A2(new_n900), .A3(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(G37), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n900), .B1(new_n944), .B2(new_n951), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n939), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n909), .A2(new_n910), .ZN(new_n957));
  NOR3_X1   g532(.A1(new_n957), .A2(new_n942), .A3(new_n943), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT41), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n959), .B1(new_n947), .B2(new_n948), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n906), .A2(KEYINPUT41), .A3(new_n908), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n962), .B1(new_n950), .B2(new_n946), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n901), .B1(new_n958), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n939), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n964), .A2(new_n953), .A3(new_n952), .A4(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n956), .A2(new_n966), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n954), .A2(new_n939), .A3(new_n955), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n964), .A2(new_n953), .A3(new_n952), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n968), .B1(KEYINPUT43), .B2(new_n969), .ZN(new_n970));
  MUX2_X1   g545(.A(new_n967), .B(new_n970), .S(KEYINPUT44), .Z(G397));
  INV_X1    g546(.A(G1384), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n865), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT45), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(G160), .A2(G40), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n770), .B(G2067), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  XOR2_X1   g554(.A(new_n979), .B(KEYINPUT107), .Z(new_n980));
  NOR3_X1   g555(.A1(new_n975), .A2(G1996), .A3(new_n976), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(new_n800), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n982), .B(KEYINPUT105), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n977), .A2(G1996), .A3(new_n799), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n985), .B(KEYINPUT106), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n711), .A2(new_n713), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n711), .A2(new_n713), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n977), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n686), .B(new_n689), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n977), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n984), .A2(new_n986), .A3(new_n989), .A4(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT108), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n992), .B(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G1976), .ZN(new_n995));
  NOR2_X1   g570(.A1(G288), .A2(new_n995), .ZN(new_n996));
  OR2_X1    g571(.A1(new_n996), .A2(KEYINPUT111), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT109), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n998), .B1(new_n857), .B2(G1384), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n862), .A2(KEYINPUT109), .A3(new_n972), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AND2_X1   g576(.A1(G160), .A2(G40), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(G8), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n996), .A2(KEYINPUT111), .ZN(new_n1006));
  AND3_X1   g581(.A1(new_n997), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT113), .ZN(new_n1008));
  XOR2_X1   g583(.A(KEYINPUT112), .B(G1976), .Z(new_n1009));
  NOR2_X1   g584(.A1(new_n889), .A2(new_n1009), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1007), .B(new_n1008), .C1(KEYINPUT52), .C2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n997), .A2(new_n1008), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n997), .A2(new_n1005), .A3(new_n1006), .A4(new_n1010), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT52), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT114), .ZN(new_n1016));
  INV_X1    g591(.A(G1981), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1017), .B1(new_n581), .B2(new_n585), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n520), .B1(new_n582), .B2(new_n583), .ZN(new_n1019));
  NOR3_X1   g594(.A1(new_n580), .A2(new_n1019), .A3(G1981), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1016), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT49), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n581), .A2(new_n585), .A3(new_n1017), .ZN(new_n1023));
  OAI21_X1  g598(.A(G1981), .B1(new_n580), .B2(new_n1019), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1023), .A2(new_n1024), .A3(KEYINPUT114), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1021), .A2(new_n1022), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT115), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1021), .A2(KEYINPUT115), .A3(new_n1022), .A4(new_n1025), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1004), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1023), .A2(new_n1024), .A3(KEYINPUT49), .ZN(new_n1031));
  AOI22_X1  g606(.A1(new_n1011), .A2(new_n1015), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT110), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT50), .B1(new_n999), .B2(new_n1000), .ZN(new_n1034));
  NOR2_X1   g609(.A1(G164), .A2(G1384), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT50), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1002), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OR2_X1    g612(.A1(new_n1034), .A2(new_n1037), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1038), .A2(G2090), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1002), .B1(new_n1035), .B2(KEYINPUT45), .ZN(new_n1040));
  AOI21_X1  g615(.A(G1384), .B1(new_n858), .B2(new_n864), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1040), .B1(new_n1041), .B2(KEYINPUT45), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1042), .A2(G1971), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1033), .B1(new_n1039), .B2(new_n1043), .ZN(new_n1044));
  OAI221_X1 g619(.A(KEYINPUT110), .B1(new_n1042), .B2(G1971), .C1(G2090), .C2(new_n1038), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1044), .A2(new_n1045), .A3(G8), .ZN(new_n1046));
  NAND2_X1  g621(.A1(G303), .A2(G8), .ZN(new_n1047));
  XNOR2_X1  g622(.A(new_n1047), .B(KEYINPUT55), .ZN(new_n1048));
  OR2_X1    g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n999), .A2(KEYINPUT50), .A3(new_n1000), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1036), .B(new_n972), .C1(new_n499), .C2(new_n504), .ZN(new_n1051));
  XNOR2_X1  g626(.A(new_n1051), .B(KEYINPUT116), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1050), .A2(new_n1052), .A3(new_n1002), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1053), .A2(G2090), .ZN(new_n1054));
  OAI21_X1  g629(.A(G8), .B1(new_n1043), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1048), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1032), .A2(new_n1049), .A3(new_n1056), .ZN(new_n1057));
  XNOR2_X1  g632(.A(KEYINPUT56), .B(G2072), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1042), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G1956), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1053), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT57), .ZN(new_n1063));
  NAND2_X1  g638(.A1(G299), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n564), .A2(KEYINPUT57), .A3(new_n567), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1062), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G2067), .ZN(new_n1069));
  NOR3_X1   g644(.A1(new_n857), .A2(new_n998), .A3(G1384), .ZN(new_n1070));
  AOI21_X1  g645(.A(KEYINPUT109), .B1(new_n862), .B2(new_n972), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1069), .B(new_n1002), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT119), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G1348), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1075), .B1(new_n1034), .B2(new_n1037), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1001), .A2(KEYINPUT119), .A3(new_n1069), .A4(new_n1002), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1074), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(new_n612), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1068), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT118), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1081), .B1(new_n1062), .B2(new_n1067), .ZN(new_n1082));
  AOI22_X1  g657(.A1(new_n1042), .A2(new_n1058), .B1(new_n1053), .B2(new_n1060), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1083), .A2(KEYINPUT118), .A3(new_n1066), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1080), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT60), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1078), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(new_n612), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT120), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1078), .A2(new_n1086), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1087), .A2(KEYINPUT120), .A3(new_n612), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1091), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT120), .B1(new_n1087), .B2(new_n612), .ZN(new_n1095));
  AOI211_X1 g670(.A(new_n1089), .B(new_n604), .C1(new_n1078), .C2(new_n1086), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1094), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1093), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1082), .A2(new_n1084), .A3(new_n1068), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT61), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(G1996), .ZN(new_n1102));
  XOR2_X1   g677(.A(KEYINPUT58), .B(G1341), .Z(new_n1103));
  AOI22_X1  g678(.A1(new_n1042), .A2(new_n1102), .B1(new_n1003), .B2(new_n1103), .ZN(new_n1104));
  OR3_X1    g679(.A1(new_n1104), .A2(KEYINPUT59), .A3(new_n552), .ZN(new_n1105));
  OAI21_X1  g680(.A(KEYINPUT59), .B1(new_n1104), .B2(new_n552), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1100), .B1(new_n1083), .B2(new_n1066), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1105), .A2(new_n1106), .B1(new_n1107), .B2(new_n1068), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1101), .A2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1085), .B1(new_n1098), .B2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n976), .B1(KEYINPUT45), .B2(new_n1035), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1111), .B1(new_n1001), .B2(KEYINPUT45), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(new_n733), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1113), .B(G168), .C1(new_n1038), .C2(G2084), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(G8), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT121), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1115), .A2(new_n1116), .A3(KEYINPUT51), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1038), .A2(G2084), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1113), .ZN(new_n1119));
  OAI211_X1 g694(.A(G8), .B(G286), .C1(new_n1118), .C2(new_n1119), .ZN(new_n1120));
  OR2_X1    g695(.A1(new_n1116), .A2(KEYINPUT51), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1116), .A2(KEYINPUT51), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1114), .A2(G8), .A3(new_n1121), .A4(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1117), .A2(new_n1120), .A3(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(KEYINPUT53), .B1(new_n1042), .B2(new_n814), .ZN(new_n1125));
  INV_X1    g700(.A(G1961), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1125), .B1(new_n1126), .B2(new_n1038), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n788), .A2(KEYINPUT123), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n788), .A2(KEYINPUT123), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(G40), .ZN(new_n1130));
  AOI211_X1 g705(.A(new_n1128), .B(new_n1130), .C1(new_n1041), .C2(KEYINPUT45), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n469), .A2(KEYINPUT53), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1131), .A2(new_n814), .A3(new_n975), .A4(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1127), .A2(new_n1133), .ZN(new_n1134));
  XOR2_X1   g709(.A(G171), .B(KEYINPUT54), .Z(new_n1135));
  OR2_X1    g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT122), .ZN(new_n1137));
  NOR3_X1   g712(.A1(new_n1112), .A2(new_n1137), .A3(G2078), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1137), .B1(new_n1112), .B2(G2078), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(KEYINPUT53), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1127), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(new_n1135), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1124), .A2(new_n1136), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1110), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1124), .A2(KEYINPUT62), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT62), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1117), .A2(new_n1120), .A3(new_n1146), .A4(new_n1123), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1145), .A2(G171), .A3(new_n1141), .A4(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1057), .B1(new_n1144), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1150), .A2(new_n1031), .A3(new_n1005), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1151), .A2(new_n995), .A3(new_n889), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(new_n1023), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1154));
  INV_X1    g729(.A(G8), .ZN(new_n1155));
  NOR3_X1   g730(.A1(new_n1154), .A2(new_n1155), .A3(G286), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT63), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1156), .A2(new_n1157), .A3(new_n1056), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1049), .A2(new_n1158), .ZN(new_n1159));
  AOI22_X1  g734(.A1(new_n1153), .A2(new_n1005), .B1(new_n1032), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT117), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1046), .A2(new_n1161), .A3(new_n1048), .ZN(new_n1162));
  OR2_X1    g737(.A1(new_n1046), .A2(new_n1161), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1032), .A2(new_n1156), .A3(new_n1162), .A4(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(KEYINPUT63), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1160), .A2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n994), .B1(new_n1149), .B2(new_n1166), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n980), .A2(new_n983), .A3(new_n987), .A4(new_n986), .ZN(new_n1168));
  OR2_X1    g743(.A1(new_n770), .A2(G2067), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(new_n977), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n977), .A2(new_n689), .A3(new_n686), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n1172), .B(KEYINPUT48), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n984), .A2(new_n986), .A3(new_n989), .A4(new_n1173), .ZN(new_n1174));
  OR2_X1    g749(.A1(new_n981), .A2(KEYINPUT46), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n977), .B1(new_n799), .B2(new_n978), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n981), .A2(KEYINPUT46), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  XOR2_X1   g753(.A(KEYINPUT124), .B(KEYINPUT47), .Z(new_n1179));
  XNOR2_X1  g754(.A(new_n1178), .B(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1171), .A2(new_n1174), .A3(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT125), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND4_X1  g758(.A1(new_n1171), .A2(KEYINPUT125), .A3(new_n1174), .A4(new_n1180), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1167), .A2(new_n1185), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g761(.A(G229), .B1(new_n880), .B2(new_n885), .ZN(new_n1188));
  INV_X1    g762(.A(G319), .ZN(new_n1189));
  OR2_X1    g763(.A1(G227), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g764(.A(KEYINPUT126), .ZN(new_n1191));
  NAND2_X1  g765(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  OR2_X1    g766(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1193));
  AND3_X1   g767(.A1(new_n649), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  NAND3_X1  g768(.A1(new_n967), .A2(new_n1188), .A3(new_n1194), .ZN(G225));
  NAND2_X1  g769(.A1(G225), .A2(KEYINPUT127), .ZN(new_n1196));
  INV_X1    g770(.A(KEYINPUT127), .ZN(new_n1197));
  NAND4_X1  g771(.A1(new_n967), .A2(new_n1188), .A3(new_n1194), .A4(new_n1197), .ZN(new_n1198));
  NAND2_X1  g772(.A1(new_n1196), .A2(new_n1198), .ZN(G308));
endmodule


