

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585;

  NOR2_X1 U325 ( .A1(n517), .A2(n451), .ZN(n565) );
  NOR2_X1 U326 ( .A1(n535), .A2(n405), .ZN(n407) );
  INV_X1 U327 ( .A(KEYINPUT69), .ZN(n371) );
  XNOR2_X1 U328 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U329 ( .A(n374), .B(n373), .ZN(n378) );
  XNOR2_X1 U330 ( .A(n414), .B(KEYINPUT48), .ZN(n540) );
  XNOR2_X1 U331 ( .A(n384), .B(n383), .ZN(n576) );
  INV_X1 U332 ( .A(G190GAT), .ZN(n452) );
  XNOR2_X1 U333 ( .A(KEYINPUT41), .B(n576), .ZN(n545) );
  XNOR2_X1 U334 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U335 ( .A(n455), .B(n454), .ZN(G1351GAT) );
  XOR2_X1 U336 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n294) );
  XNOR2_X1 U337 ( .A(KEYINPUT18), .B(KEYINPUT85), .ZN(n293) );
  XNOR2_X1 U338 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U339 ( .A(G169GAT), .B(n295), .Z(n427) );
  XOR2_X1 U340 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n297) );
  XNOR2_X1 U341 ( .A(G183GAT), .B(KEYINPUT83), .ZN(n296) );
  XNOR2_X1 U342 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U343 ( .A(KEYINPUT86), .B(G71GAT), .Z(n299) );
  XNOR2_X1 U344 ( .A(G43GAT), .B(G134GAT), .ZN(n298) );
  XNOR2_X1 U345 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U346 ( .A(n301), .B(n300), .ZN(n311) );
  XOR2_X1 U347 ( .A(KEYINPUT81), .B(KEYINPUT0), .Z(n303) );
  XNOR2_X1 U348 ( .A(KEYINPUT82), .B(G120GAT), .ZN(n302) );
  XNOR2_X1 U349 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U350 ( .A(G113GAT), .B(n304), .Z(n446) );
  XOR2_X1 U351 ( .A(G190GAT), .B(G99GAT), .Z(n306) );
  XOR2_X1 U352 ( .A(G15GAT), .B(G127GAT), .Z(n399) );
  XNOR2_X1 U353 ( .A(n399), .B(G176GAT), .ZN(n305) );
  XNOR2_X1 U354 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U355 ( .A(n446), .B(n307), .Z(n309) );
  NAND2_X1 U356 ( .A1(G227GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U357 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U358 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U359 ( .A(n427), .B(n312), .Z(n527) );
  INV_X1 U360 ( .A(n527), .ZN(n517) );
  XOR2_X1 U361 ( .A(G204GAT), .B(KEYINPUT23), .Z(n314) );
  XNOR2_X1 U362 ( .A(KEYINPUT90), .B(G211GAT), .ZN(n313) );
  XNOR2_X1 U363 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U364 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n316) );
  XOR2_X1 U365 ( .A(G50GAT), .B(G162GAT), .Z(n337) );
  XOR2_X1 U366 ( .A(G22GAT), .B(G155GAT), .Z(n398) );
  XNOR2_X1 U367 ( .A(n337), .B(n398), .ZN(n315) );
  XNOR2_X1 U368 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U369 ( .A(n318), .B(n317), .Z(n320) );
  NAND2_X1 U370 ( .A1(G228GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U371 ( .A(n320), .B(n319), .ZN(n323) );
  XOR2_X1 U372 ( .A(G78GAT), .B(G148GAT), .Z(n322) );
  XNOR2_X1 U373 ( .A(G106GAT), .B(KEYINPUT70), .ZN(n321) );
  XNOR2_X1 U374 ( .A(n322), .B(n321), .ZN(n367) );
  XOR2_X1 U375 ( .A(n323), .B(n367), .Z(n330) );
  XOR2_X1 U376 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n325) );
  XNOR2_X1 U377 ( .A(KEYINPUT89), .B(KEYINPUT88), .ZN(n324) );
  XNOR2_X1 U378 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U379 ( .A(G141GAT), .B(n326), .Z(n445) );
  XOR2_X1 U380 ( .A(KEYINPUT87), .B(KEYINPUT21), .Z(n328) );
  XNOR2_X1 U381 ( .A(G197GAT), .B(G218GAT), .ZN(n327) );
  XNOR2_X1 U382 ( .A(n328), .B(n327), .ZN(n417) );
  XNOR2_X1 U383 ( .A(n445), .B(n417), .ZN(n329) );
  XNOR2_X1 U384 ( .A(n330), .B(n329), .ZN(n466) );
  XOR2_X1 U385 ( .A(KEYINPUT66), .B(KEYINPUT7), .Z(n332) );
  XNOR2_X1 U386 ( .A(G43GAT), .B(G29GAT), .ZN(n331) );
  XNOR2_X1 U387 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U388 ( .A(KEYINPUT8), .B(n333), .Z(n366) );
  INV_X1 U389 ( .A(n366), .ZN(n349) );
  XOR2_X1 U390 ( .A(G99GAT), .B(G85GAT), .Z(n370) );
  XOR2_X1 U391 ( .A(G36GAT), .B(G190GAT), .Z(n421) );
  XOR2_X1 U392 ( .A(n370), .B(n421), .Z(n335) );
  NAND2_X1 U393 ( .A1(G232GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U394 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U395 ( .A(G92GAT), .B(n336), .ZN(n347) );
  XOR2_X1 U396 ( .A(KEYINPUT74), .B(KEYINPUT11), .Z(n339) );
  XOR2_X1 U397 ( .A(G134GAT), .B(KEYINPUT75), .Z(n438) );
  XNOR2_X1 U398 ( .A(n337), .B(n438), .ZN(n338) );
  XNOR2_X1 U399 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U400 ( .A(n340), .B(KEYINPUT10), .Z(n345) );
  XOR2_X1 U401 ( .A(KEYINPUT73), .B(KEYINPUT76), .Z(n342) );
  XNOR2_X1 U402 ( .A(G106GAT), .B(KEYINPUT9), .ZN(n341) );
  XNOR2_X1 U403 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U404 ( .A(G218GAT), .B(n343), .ZN(n344) );
  XNOR2_X1 U405 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U406 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U407 ( .A(n349), .B(n348), .Z(n535) );
  XOR2_X1 U408 ( .A(G1GAT), .B(KEYINPUT64), .Z(n351) );
  XNOR2_X1 U409 ( .A(G8GAT), .B(KEYINPUT29), .ZN(n350) );
  XNOR2_X1 U410 ( .A(n351), .B(n350), .ZN(n364) );
  XOR2_X1 U411 ( .A(G113GAT), .B(G50GAT), .Z(n353) );
  XNOR2_X1 U412 ( .A(G169GAT), .B(G36GAT), .ZN(n352) );
  XNOR2_X1 U413 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U414 ( .A(G22GAT), .B(G141GAT), .Z(n355) );
  XNOR2_X1 U415 ( .A(G15GAT), .B(G197GAT), .ZN(n354) );
  XNOR2_X1 U416 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U417 ( .A(n357), .B(n356), .Z(n362) );
  XOR2_X1 U418 ( .A(KEYINPUT30), .B(KEYINPUT65), .Z(n359) );
  NAND2_X1 U419 ( .A1(G229GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U420 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U421 ( .A(KEYINPUT67), .B(n360), .ZN(n361) );
  XNOR2_X1 U422 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U423 ( .A(n364), .B(n363), .Z(n365) );
  XOR2_X1 U424 ( .A(n366), .B(n365), .Z(n571) );
  XNOR2_X1 U425 ( .A(n367), .B(KEYINPUT32), .ZN(n369) );
  AND2_X1 U426 ( .A1(G230GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U427 ( .A(n369), .B(n368), .ZN(n374) );
  XNOR2_X1 U428 ( .A(G120GAT), .B(n370), .ZN(n372) );
  XOR2_X1 U429 ( .A(KEYINPUT31), .B(KEYINPUT72), .Z(n376) );
  XNOR2_X1 U430 ( .A(KEYINPUT33), .B(KEYINPUT71), .ZN(n375) );
  XOR2_X1 U431 ( .A(n376), .B(n375), .Z(n377) );
  XNOR2_X1 U432 ( .A(n378), .B(n377), .ZN(n384) );
  XOR2_X1 U433 ( .A(G64GAT), .B(G92GAT), .Z(n380) );
  XNOR2_X1 U434 ( .A(G176GAT), .B(G204GAT), .ZN(n379) );
  XNOR2_X1 U435 ( .A(n380), .B(n379), .ZN(n416) );
  XOR2_X1 U436 ( .A(KEYINPUT13), .B(KEYINPUT68), .Z(n382) );
  XNOR2_X1 U437 ( .A(G71GAT), .B(G57GAT), .ZN(n381) );
  XNOR2_X1 U438 ( .A(n382), .B(n381), .ZN(n397) );
  XNOR2_X1 U439 ( .A(n416), .B(n397), .ZN(n383) );
  INV_X1 U440 ( .A(n545), .ZN(n562) );
  NAND2_X1 U441 ( .A1(n571), .A2(n562), .ZN(n385) );
  XNOR2_X1 U442 ( .A(n385), .B(KEYINPUT46), .ZN(n404) );
  XOR2_X1 U443 ( .A(KEYINPUT12), .B(G64GAT), .Z(n387) );
  XNOR2_X1 U444 ( .A(G1GAT), .B(G78GAT), .ZN(n386) );
  XNOR2_X1 U445 ( .A(n387), .B(n386), .ZN(n393) );
  XOR2_X1 U446 ( .A(KEYINPUT77), .B(G211GAT), .Z(n389) );
  XNOR2_X1 U447 ( .A(G8GAT), .B(G183GAT), .ZN(n388) );
  XNOR2_X1 U448 ( .A(n389), .B(n388), .ZN(n415) );
  XOR2_X1 U449 ( .A(KEYINPUT14), .B(n415), .Z(n391) );
  NAND2_X1 U450 ( .A1(G231GAT), .A2(G233GAT), .ZN(n390) );
  XNOR2_X1 U451 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U452 ( .A(n393), .B(n392), .ZN(n403) );
  XOR2_X1 U453 ( .A(KEYINPUT80), .B(KEYINPUT79), .Z(n395) );
  XNOR2_X1 U454 ( .A(KEYINPUT78), .B(KEYINPUT15), .ZN(n394) );
  XNOR2_X1 U455 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U456 ( .A(n397), .B(n396), .Z(n401) );
  XNOR2_X1 U457 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U458 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U459 ( .A(n403), .B(n402), .ZN(n580) );
  XNOR2_X1 U460 ( .A(KEYINPUT114), .B(n580), .ZN(n567) );
  NAND2_X1 U461 ( .A1(n404), .A2(n567), .ZN(n405) );
  XNOR2_X1 U462 ( .A(KEYINPUT47), .B(KEYINPUT115), .ZN(n406) );
  XNOR2_X1 U463 ( .A(n407), .B(n406), .ZN(n413) );
  XNOR2_X1 U464 ( .A(n535), .B(KEYINPUT99), .ZN(n408) );
  XNOR2_X1 U465 ( .A(KEYINPUT36), .B(n408), .ZN(n583) );
  NOR2_X1 U466 ( .A1(n580), .A2(n583), .ZN(n409) );
  XNOR2_X1 U467 ( .A(n409), .B(KEYINPUT45), .ZN(n410) );
  INV_X1 U468 ( .A(n571), .ZN(n543) );
  NAND2_X1 U469 ( .A1(n410), .A2(n543), .ZN(n411) );
  NOR2_X1 U470 ( .A1(n576), .A2(n411), .ZN(n412) );
  NOR2_X1 U471 ( .A1(n413), .A2(n412), .ZN(n414) );
  XNOR2_X1 U472 ( .A(n416), .B(n415), .ZN(n425) );
  XOR2_X1 U473 ( .A(n417), .B(KEYINPUT94), .Z(n419) );
  NAND2_X1 U474 ( .A1(G226GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U475 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U476 ( .A(n420), .B(KEYINPUT95), .Z(n423) );
  XNOR2_X1 U477 ( .A(n421), .B(KEYINPUT93), .ZN(n422) );
  XNOR2_X1 U478 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U479 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U480 ( .A(n427), .B(n426), .ZN(n515) );
  NOR2_X1 U481 ( .A1(n540), .A2(n515), .ZN(n428) );
  XNOR2_X1 U482 ( .A(KEYINPUT54), .B(n428), .ZN(n449) );
  XOR2_X1 U483 ( .A(G85GAT), .B(G162GAT), .Z(n430) );
  XNOR2_X1 U484 ( .A(G29GAT), .B(G127GAT), .ZN(n429) );
  XNOR2_X1 U485 ( .A(n430), .B(n429), .ZN(n434) );
  XOR2_X1 U486 ( .A(G57GAT), .B(G155GAT), .Z(n432) );
  XNOR2_X1 U487 ( .A(G1GAT), .B(G148GAT), .ZN(n431) );
  XNOR2_X1 U488 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U489 ( .A(n434), .B(n433), .Z(n440) );
  XOR2_X1 U490 ( .A(KEYINPUT92), .B(KEYINPUT91), .Z(n436) );
  NAND2_X1 U491 ( .A1(G225GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U492 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U493 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U494 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U495 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n442) );
  XNOR2_X1 U496 ( .A(KEYINPUT4), .B(KEYINPUT5), .ZN(n441) );
  XNOR2_X1 U497 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U498 ( .A(n444), .B(n443), .Z(n448) );
  XNOR2_X1 U499 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U500 ( .A(n448), .B(n447), .Z(n464) );
  INV_X1 U501 ( .A(n464), .ZN(n512) );
  NAND2_X1 U502 ( .A1(n449), .A2(n512), .ZN(n569) );
  NOR2_X1 U503 ( .A1(n466), .A2(n569), .ZN(n450) );
  XNOR2_X1 U504 ( .A(n450), .B(KEYINPUT55), .ZN(n451) );
  NAND2_X1 U505 ( .A1(n565), .A2(n535), .ZN(n455) );
  XOR2_X1 U506 ( .A(KEYINPUT126), .B(KEYINPUT58), .Z(n453) );
  XOR2_X1 U507 ( .A(KEYINPUT96), .B(KEYINPUT34), .Z(n457) );
  XNOR2_X1 U508 ( .A(G1GAT), .B(KEYINPUT97), .ZN(n456) );
  XNOR2_X1 U509 ( .A(n457), .B(n456), .ZN(n472) );
  NOR2_X1 U510 ( .A1(n576), .A2(n543), .ZN(n483) );
  NOR2_X1 U511 ( .A1(n517), .A2(n515), .ZN(n458) );
  NOR2_X1 U512 ( .A1(n466), .A2(n458), .ZN(n459) );
  XOR2_X1 U513 ( .A(KEYINPUT25), .B(n459), .Z(n462) );
  XNOR2_X1 U514 ( .A(KEYINPUT27), .B(n515), .ZN(n465) );
  NAND2_X1 U515 ( .A1(n517), .A2(n466), .ZN(n460) );
  XNOR2_X1 U516 ( .A(n460), .B(KEYINPUT26), .ZN(n570) );
  NOR2_X1 U517 ( .A1(n465), .A2(n570), .ZN(n461) );
  NOR2_X1 U518 ( .A1(n462), .A2(n461), .ZN(n463) );
  NOR2_X1 U519 ( .A1(n464), .A2(n463), .ZN(n468) );
  NOR2_X1 U520 ( .A1(n512), .A2(n465), .ZN(n542) );
  XOR2_X1 U521 ( .A(n466), .B(KEYINPUT28), .Z(n521) );
  NAND2_X1 U522 ( .A1(n542), .A2(n521), .ZN(n525) );
  NOR2_X1 U523 ( .A1(n527), .A2(n525), .ZN(n467) );
  NOR2_X1 U524 ( .A1(n468), .A2(n467), .ZN(n479) );
  NOR2_X1 U525 ( .A1(n580), .A2(n535), .ZN(n469) );
  XOR2_X1 U526 ( .A(KEYINPUT16), .B(n469), .Z(n470) );
  NOR2_X1 U527 ( .A1(n479), .A2(n470), .ZN(n498) );
  NAND2_X1 U528 ( .A1(n483), .A2(n498), .ZN(n477) );
  NOR2_X1 U529 ( .A1(n512), .A2(n477), .ZN(n471) );
  XOR2_X1 U530 ( .A(n472), .B(n471), .Z(G1324GAT) );
  NOR2_X1 U531 ( .A1(n515), .A2(n477), .ZN(n473) );
  XOR2_X1 U532 ( .A(G8GAT), .B(n473), .Z(G1325GAT) );
  NOR2_X1 U533 ( .A1(n517), .A2(n477), .ZN(n475) );
  XNOR2_X1 U534 ( .A(KEYINPUT98), .B(KEYINPUT35), .ZN(n474) );
  XNOR2_X1 U535 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U536 ( .A(G15GAT), .B(n476), .ZN(G1326GAT) );
  NOR2_X1 U537 ( .A1(n521), .A2(n477), .ZN(n478) );
  XOR2_X1 U538 ( .A(G22GAT), .B(n478), .Z(G1327GAT) );
  NOR2_X1 U539 ( .A1(n479), .A2(n583), .ZN(n480) );
  NAND2_X1 U540 ( .A1(n580), .A2(n480), .ZN(n482) );
  XNOR2_X1 U541 ( .A(KEYINPUT100), .B(KEYINPUT37), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n482), .B(n481), .ZN(n510) );
  NAND2_X1 U543 ( .A1(n510), .A2(n483), .ZN(n484) );
  XOR2_X1 U544 ( .A(KEYINPUT38), .B(n484), .Z(n485) );
  XNOR2_X1 U545 ( .A(KEYINPUT101), .B(n485), .ZN(n495) );
  NOR2_X1 U546 ( .A1(n495), .A2(n512), .ZN(n489) );
  XOR2_X1 U547 ( .A(KEYINPUT102), .B(KEYINPUT39), .Z(n487) );
  XNOR2_X1 U548 ( .A(G29GAT), .B(KEYINPUT103), .ZN(n486) );
  XNOR2_X1 U549 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U550 ( .A(n489), .B(n488), .ZN(G1328GAT) );
  NOR2_X1 U551 ( .A1(n495), .A2(n515), .ZN(n490) );
  XOR2_X1 U552 ( .A(KEYINPUT104), .B(n490), .Z(n491) );
  XNOR2_X1 U553 ( .A(G36GAT), .B(n491), .ZN(G1329GAT) );
  NOR2_X1 U554 ( .A1(n495), .A2(n517), .ZN(n493) );
  XNOR2_X1 U555 ( .A(KEYINPUT105), .B(KEYINPUT40), .ZN(n492) );
  XNOR2_X1 U556 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U557 ( .A(G43GAT), .B(n494), .ZN(G1330GAT) );
  NOR2_X1 U558 ( .A1(n521), .A2(n495), .ZN(n496) );
  XOR2_X1 U559 ( .A(KEYINPUT106), .B(n496), .Z(n497) );
  XNOR2_X1 U560 ( .A(G50GAT), .B(n497), .ZN(G1331GAT) );
  NOR2_X1 U561 ( .A1(n571), .A2(n545), .ZN(n511) );
  NAND2_X1 U562 ( .A1(n511), .A2(n498), .ZN(n505) );
  NOR2_X1 U563 ( .A1(n512), .A2(n505), .ZN(n499) );
  XOR2_X1 U564 ( .A(G57GAT), .B(n499), .Z(n500) );
  XNOR2_X1 U565 ( .A(KEYINPUT42), .B(n500), .ZN(G1332GAT) );
  NOR2_X1 U566 ( .A1(n515), .A2(n505), .ZN(n501) );
  XOR2_X1 U567 ( .A(G64GAT), .B(n501), .Z(G1333GAT) );
  NOR2_X1 U568 ( .A1(n517), .A2(n505), .ZN(n503) );
  XNOR2_X1 U569 ( .A(KEYINPUT107), .B(KEYINPUT108), .ZN(n502) );
  XNOR2_X1 U570 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U571 ( .A(G71GAT), .B(n504), .ZN(G1334GAT) );
  NOR2_X1 U572 ( .A1(n505), .A2(n521), .ZN(n509) );
  XOR2_X1 U573 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n507) );
  XNOR2_X1 U574 ( .A(G78GAT), .B(KEYINPUT110), .ZN(n506) );
  XNOR2_X1 U575 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U576 ( .A(n509), .B(n508), .ZN(G1335GAT) );
  NAND2_X1 U577 ( .A1(n511), .A2(n510), .ZN(n520) );
  NOR2_X1 U578 ( .A1(n512), .A2(n520), .ZN(n514) );
  XNOR2_X1 U579 ( .A(G85GAT), .B(KEYINPUT111), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n514), .B(n513), .ZN(G1336GAT) );
  NOR2_X1 U581 ( .A1(n515), .A2(n520), .ZN(n516) );
  XOR2_X1 U582 ( .A(G92GAT), .B(n516), .Z(G1337GAT) );
  NOR2_X1 U583 ( .A1(n517), .A2(n520), .ZN(n518) );
  XOR2_X1 U584 ( .A(KEYINPUT112), .B(n518), .Z(n519) );
  XNOR2_X1 U585 ( .A(G99GAT), .B(n519), .ZN(G1338GAT) );
  NOR2_X1 U586 ( .A1(n521), .A2(n520), .ZN(n523) );
  XNOR2_X1 U587 ( .A(KEYINPUT44), .B(KEYINPUT113), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(n524), .ZN(G1339GAT) );
  NOR2_X1 U590 ( .A1(n540), .A2(n525), .ZN(n526) );
  NAND2_X1 U591 ( .A1(n527), .A2(n526), .ZN(n536) );
  NOR2_X1 U592 ( .A1(n543), .A2(n536), .ZN(n528) );
  XOR2_X1 U593 ( .A(G113GAT), .B(n528), .Z(G1340GAT) );
  NOR2_X1 U594 ( .A1(n545), .A2(n536), .ZN(n530) );
  XNOR2_X1 U595 ( .A(KEYINPUT49), .B(KEYINPUT116), .ZN(n529) );
  XNOR2_X1 U596 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U597 ( .A(G120GAT), .B(n531), .ZN(G1341GAT) );
  NOR2_X1 U598 ( .A1(n567), .A2(n536), .ZN(n533) );
  XNOR2_X1 U599 ( .A(KEYINPUT50), .B(KEYINPUT117), .ZN(n532) );
  XNOR2_X1 U600 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(n534), .ZN(G1342GAT) );
  INV_X1 U602 ( .A(n535), .ZN(n554) );
  NOR2_X1 U603 ( .A1(n554), .A2(n536), .ZN(n538) );
  XNOR2_X1 U604 ( .A(KEYINPUT118), .B(KEYINPUT51), .ZN(n537) );
  XNOR2_X1 U605 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U606 ( .A(G134GAT), .B(n539), .ZN(G1343GAT) );
  NOR2_X1 U607 ( .A1(n570), .A2(n540), .ZN(n541) );
  NAND2_X1 U608 ( .A1(n542), .A2(n541), .ZN(n553) );
  NOR2_X1 U609 ( .A1(n543), .A2(n553), .ZN(n544) );
  XOR2_X1 U610 ( .A(G141GAT), .B(n544), .Z(G1344GAT) );
  NOR2_X1 U611 ( .A1(n553), .A2(n545), .ZN(n549) );
  XOR2_X1 U612 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n547) );
  XNOR2_X1 U613 ( .A(G148GAT), .B(KEYINPUT119), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(G1345GAT) );
  NOR2_X1 U616 ( .A1(n580), .A2(n553), .ZN(n551) );
  XNOR2_X1 U617 ( .A(KEYINPUT120), .B(KEYINPUT121), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U619 ( .A(G155GAT), .B(n552), .ZN(G1346GAT) );
  NOR2_X1 U620 ( .A1(n554), .A2(n553), .ZN(n556) );
  XNOR2_X1 U621 ( .A(KEYINPUT122), .B(KEYINPUT123), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U623 ( .A(G162GAT), .B(n557), .ZN(G1347GAT) );
  NAND2_X1 U624 ( .A1(n571), .A2(n565), .ZN(n558) );
  XNOR2_X1 U625 ( .A(G169GAT), .B(n558), .ZN(G1348GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT57), .B(KEYINPUT125), .Z(n560) );
  XNOR2_X1 U627 ( .A(G176GAT), .B(KEYINPUT124), .ZN(n559) );
  XNOR2_X1 U628 ( .A(n560), .B(n559), .ZN(n561) );
  XOR2_X1 U629 ( .A(KEYINPUT56), .B(n561), .Z(n564) );
  NAND2_X1 U630 ( .A1(n565), .A2(n562), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(G1349GAT) );
  INV_X1 U632 ( .A(n565), .ZN(n566) );
  NOR2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U634 ( .A(G183GAT), .B(n568), .Z(G1350GAT) );
  XOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT59), .Z(n573) );
  NOR2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n579) );
  NAND2_X1 U637 ( .A1(n579), .A2(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n575) );
  XOR2_X1 U639 ( .A(KEYINPUT60), .B(KEYINPUT127), .Z(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1352GAT) );
  XOR2_X1 U641 ( .A(G204GAT), .B(KEYINPUT61), .Z(n578) );
  NAND2_X1 U642 ( .A1(n579), .A2(n576), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1353GAT) );
  INV_X1 U644 ( .A(n579), .ZN(n582) );
  OR2_X1 U645 ( .A1(n582), .A2(n580), .ZN(n581) );
  XNOR2_X1 U646 ( .A(G211GAT), .B(n581), .ZN(G1354GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U648 ( .A(KEYINPUT62), .B(n584), .Z(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

