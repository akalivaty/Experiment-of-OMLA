//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 1 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 0 1 0 0 1 0 0 0 1 1 1 1 0 1 1 0 1 1 1 0 0 1 0 1 1 1 1 1 1 0 1 1 1 0 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:38 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  INV_X1    g0011(.A(G58), .ZN(new_n212));
  INV_X1    g0012(.A(G68), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n206), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g0019(.A(KEYINPUT64), .B(G77), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G68), .A2(G238), .B1(G97), .B2(G257), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G58), .B2(G232), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G107), .A2(G264), .ZN(new_n226));
  NAND4_X1  g0026(.A1(new_n223), .A2(new_n224), .A3(new_n225), .A4(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n208), .B1(new_n222), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n211), .B(new_n219), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n235), .B(new_n238), .Z(G358));
  XOR2_X1   g0039(.A(G68), .B(G77), .Z(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G58), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(new_n220), .ZN(new_n247));
  AND2_X1   g0047(.A1(KEYINPUT3), .A2(G33), .ZN(new_n248));
  NOR2_X1   g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G1698), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT3), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n252), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G223), .ZN(new_n258));
  AOI21_X1  g0058(.A(G1698), .B1(new_n255), .B2(new_n256), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(KEYINPUT66), .A3(G222), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(KEYINPUT66), .B1(new_n259), .B2(G222), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n251), .B(new_n258), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G41), .ZN(new_n266));
  INV_X1    g0066(.A(G45), .ZN(new_n267));
  AOI21_X1  g0067(.A(G1), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G226), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT65), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(KEYINPUT65), .ZN(new_n274));
  OAI211_X1 g0074(.A(G1), .B(G13), .C1(new_n254), .C2(new_n266), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n272), .A2(G274), .A3(new_n274), .A4(new_n275), .ZN(new_n276));
  AND2_X1   g0076(.A1(new_n270), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n265), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G169), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n217), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G50), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n286), .B1(new_n205), .B2(G20), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n285), .A2(new_n287), .B1(new_n286), .B2(new_n282), .ZN(new_n288));
  NOR2_X1   g0088(.A1(G50), .A2(G58), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n206), .B1(new_n289), .B2(new_n213), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n206), .A2(new_n254), .ZN(new_n291));
  INV_X1    g0091(.A(G150), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  XOR2_X1   g0093(.A(KEYINPUT8), .B(G58), .Z(new_n294));
  NOR2_X1   g0094(.A1(new_n254), .A2(G20), .ZN(new_n295));
  AOI211_X1 g0095(.A(new_n290), .B(new_n293), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n284), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n288), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n270), .A2(new_n276), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n299), .B1(new_n263), .B2(new_n264), .ZN(new_n300));
  INV_X1    g0100(.A(G179), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AND3_X1   g0102(.A1(new_n280), .A2(new_n298), .A3(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT68), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n300), .A2(new_n304), .A3(G190), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n304), .B1(new_n300), .B2(G190), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n278), .A2(G200), .ZN(new_n309));
  INV_X1    g0109(.A(new_n298), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT9), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT9), .ZN(new_n312));
  AOI21_X1  g0112(.A(KEYINPUT67), .B1(new_n298), .B2(new_n312), .ZN(new_n313));
  AND3_X1   g0113(.A1(new_n298), .A2(KEYINPUT67), .A3(new_n312), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n309), .B(new_n311), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(KEYINPUT10), .B1(new_n308), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n307), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(new_n305), .ZN(new_n318));
  AND2_X1   g0118(.A1(new_n309), .A2(new_n311), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT10), .ZN(new_n320));
  OR2_X1    g0120(.A1(new_n314), .A2(new_n313), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n318), .A2(new_n319), .A3(new_n320), .A4(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n303), .B1(new_n316), .B2(new_n322), .ZN(new_n323));
  NOR2_X1   g0123(.A1(G20), .A2(G33), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n324), .A2(G50), .B1(G20), .B2(new_n213), .ZN(new_n325));
  INV_X1    g0125(.A(new_n295), .ZN(new_n326));
  INV_X1    g0126(.A(G77), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n325), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n284), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT11), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n328), .A2(KEYINPUT11), .A3(new_n284), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n205), .A2(G20), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n297), .A2(G68), .A3(new_n281), .A4(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT12), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n336), .B1(new_n282), .B2(new_n213), .ZN(new_n337));
  NOR3_X1   g0137(.A1(new_n281), .A2(KEYINPUT12), .A3(G68), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n335), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT71), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n335), .B(KEYINPUT71), .C1(new_n337), .C2(new_n338), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n333), .A2(KEYINPUT72), .A3(new_n341), .A4(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT72), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n331), .A2(new_n342), .A3(new_n332), .ZN(new_n345));
  AND2_X1   g0145(.A1(new_n339), .A2(new_n340), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n344), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n343), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n269), .A2(G238), .ZN(new_n350));
  NOR2_X1   g0150(.A1(G226), .A2(G1698), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n351), .B1(new_n232), .B2(G1698), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n255), .A2(new_n256), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n352), .A2(new_n353), .B1(G33), .B2(G97), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n350), .B(new_n276), .C1(new_n354), .C2(new_n275), .ZN(new_n355));
  XNOR2_X1  g0155(.A(KEYINPUT69), .B(KEYINPUT13), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(G33), .A2(G97), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n232), .A2(G1698), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(G226), .B2(G1698), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n359), .B1(new_n361), .B2(new_n250), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n264), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n363), .A2(new_n276), .A3(new_n356), .A4(new_n350), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n358), .A2(KEYINPUT70), .A3(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT70), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n355), .A2(new_n366), .A3(new_n357), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n365), .A2(G169), .A3(new_n367), .ZN(new_n368));
  AND2_X1   g0168(.A1(new_n368), .A2(KEYINPUT14), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT14), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n365), .A2(new_n370), .A3(G169), .A4(new_n367), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n355), .A2(KEYINPUT13), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n372), .A2(G179), .A3(new_n364), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n349), .B1(new_n369), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n365), .A2(G200), .A3(new_n367), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n372), .A2(G190), .A3(new_n364), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n348), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(G232), .A2(G1698), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n252), .A2(G238), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n353), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n381), .B(new_n264), .C1(G107), .C2(new_n353), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n269), .A2(G244), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n382), .A2(new_n276), .A3(new_n383), .ZN(new_n384));
  OR2_X1    g0184(.A1(new_n384), .A2(G179), .ZN(new_n385));
  AND2_X1   g0185(.A1(new_n294), .A2(new_n324), .ZN(new_n386));
  XNOR2_X1  g0186(.A(KEYINPUT15), .B(G87), .ZN(new_n387));
  OAI22_X1  g0187(.A1(new_n326), .A2(new_n387), .B1(new_n220), .B2(new_n206), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n284), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n327), .B1(new_n205), .B2(G20), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n285), .A2(new_n390), .B1(new_n220), .B2(new_n282), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n384), .A2(new_n279), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n385), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n392), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n384), .A2(G200), .ZN(new_n396));
  INV_X1    g0196(.A(G190), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n395), .B(new_n396), .C1(new_n397), .C2(new_n384), .ZN(new_n398));
  AND2_X1   g0198(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n323), .A2(new_n375), .A3(new_n378), .A4(new_n399), .ZN(new_n400));
  OAI211_X1 g0200(.A(G226), .B(G1698), .C1(new_n248), .C2(new_n249), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT75), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n353), .A2(KEYINPUT75), .A3(G226), .A4(G1698), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n259), .A2(G223), .B1(G33), .B2(G87), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n275), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n269), .A2(G232), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n276), .ZN(new_n409));
  OAI21_X1  g0209(.A(G200), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  AND2_X1   g0210(.A1(new_n408), .A2(new_n276), .ZN(new_n411));
  OAI211_X1 g0211(.A(G223), .B(new_n252), .C1(new_n248), .C2(new_n249), .ZN(new_n412));
  INV_X1    g0212(.A(G87), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n412), .B1(new_n254), .B2(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n414), .B1(new_n403), .B2(new_n404), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n411), .B(G190), .C1(new_n415), .C2(new_n275), .ZN(new_n416));
  AND2_X1   g0216(.A1(new_n410), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(KEYINPUT7), .B1(new_n250), .B2(new_n206), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n255), .A2(KEYINPUT7), .A3(new_n206), .A4(new_n256), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(G68), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(G58), .A2(G68), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NOR2_X1   g0223(.A1(G58), .A2(G68), .ZN(new_n424));
  OAI21_X1  g0224(.A(G20), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n324), .A2(G159), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n421), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT16), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n297), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT74), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n255), .A2(new_n206), .A3(new_n256), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT7), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n419), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n206), .B1(new_n214), .B2(new_n422), .ZN(new_n435));
  INV_X1    g0235(.A(G159), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n291), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(KEYINPUT73), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT73), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n425), .A2(new_n439), .A3(new_n426), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n434), .A2(G68), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n430), .B1(new_n441), .B2(KEYINPUT16), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n438), .A2(new_n440), .ZN(new_n443));
  AND4_X1   g0243(.A1(new_n430), .A2(new_n443), .A3(new_n421), .A4(KEYINPUT16), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n429), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n285), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n294), .A2(new_n334), .ZN(new_n447));
  OAI22_X1  g0247(.A1(new_n446), .A2(new_n447), .B1(new_n281), .B2(new_n294), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n417), .A2(new_n445), .A3(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT77), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT17), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n443), .A2(new_n421), .A3(KEYINPUT16), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT74), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n441), .A2(new_n430), .A3(KEYINPUT16), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n448), .B1(new_n457), .B2(new_n429), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n451), .A2(new_n452), .ZN(new_n459));
  NAND2_X1  g0259(.A1(KEYINPUT77), .A2(KEYINPUT17), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n458), .A2(new_n459), .A3(new_n460), .A4(new_n417), .ZN(new_n461));
  AND2_X1   g0261(.A1(new_n453), .A2(new_n461), .ZN(new_n462));
  OAI21_X1  g0262(.A(G169), .B1(new_n407), .B2(new_n409), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n411), .B(G179), .C1(new_n415), .C2(new_n275), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  OAI21_X1  g0266(.A(KEYINPUT18), .B1(new_n458), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT76), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT18), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n213), .B1(new_n433), .B2(new_n419), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n425), .A2(new_n426), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n428), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n284), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n473), .B1(new_n455), .B2(new_n456), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n469), .B(new_n465), .C1(new_n474), .C2(new_n448), .ZN(new_n475));
  AND3_X1   g0275(.A1(new_n467), .A2(new_n468), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n468), .B1(new_n467), .B2(new_n475), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n462), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n205), .B(G45), .C1(new_n266), .C2(KEYINPUT5), .ZN(new_n479));
  INV_X1    g0279(.A(G274), .ZN(new_n480));
  NOR3_X1   g0280(.A1(new_n264), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT5), .ZN(new_n482));
  OAI21_X1  g0282(.A(KEYINPUT80), .B1(new_n482), .B2(G41), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT80), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n484), .A2(new_n266), .A3(KEYINPUT5), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT81), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n483), .A2(new_n485), .A3(KEYINPUT81), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n481), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT82), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n481), .A2(new_n488), .A3(KEYINPUT82), .A4(new_n489), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n353), .A2(KEYINPUT4), .A3(G244), .A4(new_n252), .ZN(new_n495));
  NAND2_X1  g0295(.A1(G33), .A2(G283), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n250), .A2(new_n221), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n495), .B(new_n496), .C1(new_n497), .C2(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n353), .A2(G250), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n252), .B1(new_n499), .B2(KEYINPUT4), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n264), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(G257), .ZN(new_n502));
  AND2_X1   g0302(.A1(new_n483), .A2(new_n485), .ZN(new_n503));
  INV_X1    g0303(.A(new_n479), .ZN(new_n504));
  AOI211_X1 g0304(.A(new_n502), .B(new_n264), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n494), .A2(new_n501), .A3(G190), .A4(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT83), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n494), .A2(new_n501), .A3(new_n506), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(G200), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n434), .A2(G107), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT78), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n434), .A2(KEYINPUT78), .A3(G107), .ZN(new_n515));
  INV_X1    g0315(.A(G107), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n516), .A2(KEYINPUT6), .A3(G97), .ZN(new_n517));
  INV_X1    g0317(.A(G97), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n518), .A2(new_n516), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n519), .A2(new_n202), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n517), .B1(new_n520), .B2(KEYINPUT6), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n521), .A2(G20), .B1(G77), .B2(new_n324), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n514), .A2(new_n515), .A3(new_n522), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n282), .A2(G97), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n205), .A2(G33), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n281), .A2(new_n525), .A3(new_n217), .A4(new_n283), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n524), .B1(G97), .B2(new_n526), .ZN(new_n527));
  OR2_X1    g0327(.A1(new_n527), .A2(KEYINPUT79), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(KEYINPUT79), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n523), .A2(new_n284), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n505), .B1(new_n492), .B2(new_n493), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n531), .A2(KEYINPUT83), .A3(G190), .A4(new_n501), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n509), .A2(new_n511), .A3(new_n530), .A4(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT23), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(new_n206), .B2(G107), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n516), .A2(KEYINPUT23), .A3(G20), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n206), .A2(G33), .A3(G116), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n206), .B(G87), .C1(new_n248), .C2(new_n249), .ZN(new_n541));
  XOR2_X1   g0341(.A(KEYINPUT86), .B(KEYINPUT22), .Z(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n541), .A2(new_n542), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n540), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT24), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n546), .A2(KEYINPUT87), .A3(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(KEYINPUT24), .B1(new_n546), .B2(KEYINPUT87), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT87), .ZN(new_n550));
  OR2_X1    g0350(.A1(new_n541), .A2(new_n542), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n543), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n550), .B1(new_n552), .B2(new_n540), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n284), .B(new_n548), .C1(new_n549), .C2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n282), .A2(new_n516), .ZN(new_n555));
  NOR2_X1   g0355(.A1(KEYINPUT88), .A2(KEYINPUT25), .ZN(new_n556));
  OR2_X1    g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AND2_X1   g0357(.A1(KEYINPUT88), .A2(KEYINPUT25), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n558), .B1(new_n555), .B2(new_n556), .ZN(new_n559));
  INV_X1    g0359(.A(new_n526), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n557), .A2(new_n559), .B1(G107), .B2(new_n560), .ZN(new_n561));
  OAI211_X1 g0361(.A(G250), .B(new_n252), .C1(new_n248), .C2(new_n249), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(KEYINPUT89), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT89), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n353), .A2(new_n564), .A3(G250), .A4(new_n252), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n353), .A2(G257), .A3(G1698), .ZN(new_n566));
  NAND2_X1  g0366(.A1(G33), .A2(G294), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n563), .A2(new_n565), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n264), .B1(new_n503), .B2(new_n504), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n568), .A2(new_n264), .B1(G264), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n494), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n571), .A2(G190), .ZN(new_n572));
  AOI21_X1  g0372(.A(G200), .B1(new_n494), .B2(new_n570), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n554), .B(new_n561), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n523), .A2(new_n284), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n528), .A2(new_n529), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n510), .A2(new_n279), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n531), .A2(new_n301), .A3(new_n501), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(G200), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n205), .A2(new_n480), .A3(G45), .ZN(new_n582));
  INV_X1    g0382(.A(G250), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(new_n267), .B2(G1), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n275), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(KEYINPUT84), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT84), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n275), .A2(new_n587), .A3(new_n582), .A4(new_n584), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n221), .A2(G1698), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n590), .B1(G238), .B2(G1698), .ZN(new_n591));
  INV_X1    g0391(.A(G116), .ZN(new_n592));
  OAI22_X1  g0392(.A1(new_n591), .A2(new_n250), .B1(new_n254), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n264), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n581), .B1(new_n589), .B2(new_n594), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n589), .A2(new_n594), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n595), .B1(G190), .B2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT19), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n598), .B1(new_n326), .B2(new_n518), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n353), .A2(new_n206), .A3(G68), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n206), .B1(new_n359), .B2(new_n598), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(G87), .B2(new_n203), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n599), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n603), .A2(new_n284), .B1(new_n282), .B2(new_n387), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n560), .A2(G87), .ZN(new_n605));
  AND2_X1   g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n597), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n533), .A2(new_n574), .A3(new_n580), .A4(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n589), .A2(G179), .A3(new_n594), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(new_n596), .B2(new_n279), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n604), .B1(new_n387), .B2(new_n526), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(G169), .B1(new_n494), .B2(new_n570), .ZN(new_n614));
  INV_X1    g0414(.A(new_n571), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n614), .B1(new_n615), .B2(new_n301), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n554), .A2(new_n561), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n613), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n257), .A2(G264), .B1(new_n250), .B2(G303), .ZN(new_n619));
  AND3_X1   g0419(.A1(new_n259), .A2(KEYINPUT85), .A3(G257), .ZN(new_n620));
  AOI21_X1  g0420(.A(KEYINPUT85), .B1(new_n259), .B2(G257), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n264), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n569), .A2(G270), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n494), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n496), .B(new_n206), .C1(G33), .C2(new_n518), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n626), .B(new_n284), .C1(new_n206), .C2(G116), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT20), .ZN(new_n628));
  XNOR2_X1  g0428(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n281), .A2(G116), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n630), .B1(new_n560), .B2(G116), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  NOR3_X1   g0433(.A1(new_n625), .A2(new_n633), .A3(new_n301), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n279), .B1(new_n629), .B2(new_n631), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n625), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(KEYINPUT21), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT21), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n625), .A2(new_n638), .A3(new_n635), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n634), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n632), .B1(new_n625), .B2(G200), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n641), .B1(new_n397), .B2(new_n625), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n618), .A2(new_n640), .A3(new_n642), .ZN(new_n643));
  NOR4_X1   g0443(.A1(new_n400), .A2(new_n478), .A3(new_n608), .A4(new_n643), .ZN(G372));
  INV_X1    g0444(.A(new_n303), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n445), .A2(new_n449), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n469), .B1(new_n646), .B2(new_n465), .ZN(new_n647));
  INV_X1    g0447(.A(new_n475), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n368), .A2(KEYINPUT14), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n650), .A2(new_n373), .A3(new_n371), .ZN(new_n651));
  INV_X1    g0451(.A(new_n394), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n651), .A2(new_n349), .B1(new_n378), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n453), .A2(new_n461), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n649), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT90), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n316), .A2(new_n322), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n658), .B1(new_n655), .B2(new_n656), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n645), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n400), .A2(new_n478), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n616), .A2(new_n617), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n640), .A2(new_n663), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n533), .A2(new_n580), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n574), .A2(new_n607), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT26), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n607), .A2(new_n612), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n668), .B1(new_n580), .B2(new_n669), .ZN(new_n670));
  AOI22_X1  g0470(.A1(new_n606), .A2(new_n597), .B1(new_n610), .B2(new_n611), .ZN(new_n671));
  AOI22_X1  g0471(.A1(new_n575), .A2(new_n576), .B1(new_n510), .B2(new_n279), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n671), .A2(new_n672), .A3(KEYINPUT26), .A4(new_n579), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n613), .B1(new_n670), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n667), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n662), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n661), .A2(new_n676), .ZN(G369));
  NAND3_X1  g0477(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(new_n680), .A3(G213), .ZN(new_n681));
  INV_X1    g0481(.A(G343), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n617), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(KEYINPUT92), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n574), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n684), .A2(KEYINPUT92), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n663), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n663), .A2(new_n683), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g0491(.A(KEYINPUT91), .B(G330), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n637), .A2(new_n639), .ZN(new_n693));
  INV_X1    g0493(.A(new_n634), .ZN(new_n694));
  AND3_X1   g0494(.A1(new_n693), .A2(new_n642), .A3(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n683), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n695), .B1(new_n633), .B2(new_n696), .ZN(new_n697));
  OR3_X1    g0497(.A1(new_n640), .A2(new_n633), .A3(new_n696), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n692), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n691), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT93), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n640), .A2(new_n683), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n689), .B1(new_n688), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n702), .A2(new_n704), .ZN(G399));
  INV_X1    g0505(.A(new_n209), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(G41), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n203), .A2(G87), .A3(G116), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n708), .A2(G1), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(new_n215), .B2(new_n708), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT28), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n683), .B1(new_n667), .B2(new_n674), .ZN(new_n713));
  XNOR2_X1  g0513(.A(KEYINPUT95), .B(KEYINPUT29), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n625), .ZN(new_n717));
  INV_X1    g0517(.A(new_n510), .ZN(new_n718));
  INV_X1    g0518(.A(new_n609), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n719), .A2(new_n570), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n717), .A2(new_n718), .A3(KEYINPUT30), .A4(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT30), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n531), .A2(new_n719), .A3(new_n501), .A4(new_n570), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n722), .B1(new_n723), .B2(new_n625), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n596), .A2(G179), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n625), .A2(new_n510), .A3(new_n571), .A4(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n721), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(KEYINPUT31), .B1(new_n727), .B2(new_n683), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n724), .A2(new_n726), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(KEYINPUT94), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT94), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n724), .A2(new_n731), .A3(new_n726), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n730), .A2(new_n732), .A3(new_n721), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT31), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n696), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n728), .B1(new_n733), .B2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n608), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n737), .A2(new_n695), .A3(new_n618), .A4(new_n696), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n692), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  AOI211_X1 g0539(.A(KEYINPUT29), .B(new_n683), .C1(new_n667), .C2(new_n674), .ZN(new_n740));
  NOR3_X1   g0540(.A1(new_n716), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n741), .B(KEYINPUT96), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n712), .B1(new_n742), .B2(G1), .ZN(G364));
  INV_X1    g0543(.A(G13), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(G20), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n205), .B1(new_n745), .B2(G45), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n707), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G13), .A2(G33), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(G20), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n217), .B1(G20), .B2(new_n279), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g0556(.A(new_n756), .B(KEYINPUT97), .ZN(new_n757));
  XOR2_X1   g0557(.A(new_n757), .B(KEYINPUT98), .Z(new_n758));
  NOR2_X1   g0558(.A1(new_n706), .A2(new_n353), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n760), .B1(new_n267), .B2(new_n216), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n761), .B1(new_n242), .B2(new_n267), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n706), .A2(new_n250), .ZN(new_n763));
  AOI22_X1  g0563(.A1(new_n763), .A2(G355), .B1(new_n592), .B2(new_n706), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n758), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(G20), .A2(G179), .ZN(new_n766));
  XOR2_X1   g0566(.A(new_n766), .B(KEYINPUT99), .Z(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G190), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(G200), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G58), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n767), .A2(new_n397), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n581), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G68), .ZN(new_n773));
  AND2_X1   g0573(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n768), .A2(new_n581), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n771), .A2(G200), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  OAI221_X1 g0578(.A(new_n774), .B1(new_n286), .B2(new_n776), .C1(new_n220), .C2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n581), .A2(G179), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n780), .A2(G20), .A3(new_n397), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT100), .Z(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n516), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G179), .A2(G200), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n785), .A2(G20), .A3(new_n397), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n436), .ZN(new_n787));
  XOR2_X1   g0587(.A(new_n787), .B(KEYINPUT32), .Z(new_n788));
  NAND3_X1  g0588(.A1(new_n780), .A2(G20), .A3(G190), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n785), .A2(G190), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G20), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n353), .B1(new_n789), .B2(new_n413), .C1(new_n792), .C2(new_n518), .ZN(new_n793));
  OR3_X1    g0593(.A1(new_n784), .A2(new_n788), .A3(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n779), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  OR2_X1    g0596(.A1(new_n796), .A2(KEYINPUT101), .ZN(new_n797));
  AOI22_X1  g0597(.A1(G311), .A2(new_n777), .B1(new_n775), .B2(G326), .ZN(new_n798));
  XNOR2_X1  g0598(.A(KEYINPUT33), .B(G317), .ZN(new_n799));
  AOI22_X1  g0599(.A1(G322), .A2(new_n769), .B1(new_n772), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n782), .A2(G283), .ZN(new_n801));
  INV_X1    g0601(.A(new_n786), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n353), .B1(new_n802), .B2(G329), .ZN(new_n803));
  INV_X1    g0603(.A(G303), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n803), .B1(new_n804), .B2(new_n789), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n805), .B1(G294), .B2(new_n791), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n798), .A2(new_n800), .A3(new_n801), .A4(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n796), .A2(KEYINPUT101), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n797), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n765), .B1(new_n809), .B2(new_n754), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n697), .A2(new_n698), .A3(new_n752), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n749), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n699), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n697), .A2(new_n692), .A3(new_n698), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n748), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT102), .ZN(G396));
  OAI21_X1  g0617(.A(new_n398), .B1(new_n395), .B2(new_n696), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(new_n394), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n652), .A2(new_n696), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n713), .B(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n739), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n748), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(new_n824), .B2(new_n823), .ZN(new_n826));
  AOI22_X1  g0626(.A1(G137), .A2(new_n775), .B1(new_n772), .B2(G150), .ZN(new_n827));
  INV_X1    g0627(.A(G143), .ZN(new_n828));
  INV_X1    g0628(.A(new_n769), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n827), .B1(new_n828), .B2(new_n829), .C1(new_n436), .C2(new_n778), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n830), .B(KEYINPUT34), .Z(new_n831));
  NOR2_X1   g0631(.A1(new_n783), .A2(new_n213), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n792), .A2(new_n212), .ZN(new_n833));
  INV_X1    g0633(.A(G132), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n353), .B1(new_n786), .B2(new_n834), .C1(new_n789), .C2(new_n286), .ZN(new_n835));
  NOR4_X1   g0635(.A1(new_n831), .A2(new_n832), .A3(new_n833), .A4(new_n835), .ZN(new_n836));
  AOI22_X1  g0636(.A1(G311), .A2(new_n802), .B1(new_n791), .B2(G97), .ZN(new_n837));
  INV_X1    g0637(.A(G283), .ZN(new_n838));
  INV_X1    g0638(.A(new_n772), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n837), .B1(new_n783), .B2(new_n413), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n250), .B1(new_n789), .B2(new_n516), .ZN(new_n841));
  XOR2_X1   g0641(.A(new_n841), .B(KEYINPUT103), .Z(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n592), .B2(new_n778), .ZN(new_n843));
  INV_X1    g0643(.A(G294), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n844), .A2(new_n829), .B1(new_n776), .B2(new_n804), .ZN(new_n845));
  NOR3_X1   g0645(.A1(new_n840), .A2(new_n843), .A3(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n754), .B1(new_n836), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n754), .A2(new_n750), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n749), .B1(new_n327), .B2(new_n848), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n847), .B(new_n849), .C1(new_n751), .C2(new_n822), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n826), .A2(new_n850), .ZN(new_n851));
  XOR2_X1   g0651(.A(new_n851), .B(KEYINPUT104), .Z(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(G384));
  NOR2_X1   g0653(.A1(new_n745), .A2(new_n205), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n349), .A2(new_n683), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n375), .A2(new_n378), .A3(new_n855), .ZN(new_n856));
  AND3_X1   g0656(.A1(new_n348), .A2(new_n376), .A3(new_n377), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n349), .B(new_n683), .C1(new_n651), .C2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n821), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  NOR3_X1   g0659(.A1(new_n643), .A2(new_n608), .A3(new_n683), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n727), .A2(new_n683), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n734), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n727), .A2(KEYINPUT31), .A3(new_n683), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n859), .B(KEYINPUT40), .C1(new_n860), .C2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT105), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n458), .B2(new_n466), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n646), .A2(KEYINPUT105), .A3(new_n465), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n681), .B(KEYINPUT106), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n474), .B2(new_n448), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT37), .ZN(new_n872));
  AND3_X1   g0672(.A1(new_n871), .A2(new_n450), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n284), .B1(new_n441), .B2(KEYINPUT16), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n875), .B1(new_n456), .B2(new_n455), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n465), .B1(new_n876), .B2(new_n448), .ZN(new_n877));
  INV_X1    g0677(.A(new_n681), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n878), .B1(new_n876), .B2(new_n448), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n877), .A2(new_n879), .A3(new_n450), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(KEYINPUT37), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n874), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT76), .B1(new_n647), .B2(new_n648), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n467), .A2(new_n468), .A3(new_n475), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n654), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI211_X1 g0685(.A(KEYINPUT38), .B(new_n882), .C1(new_n885), .C2(new_n879), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT38), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n871), .B1(new_n462), .B2(new_n649), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n871), .B(new_n450), .C1(new_n458), .C2(new_n466), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n869), .A2(new_n873), .B1(new_n889), .B2(KEYINPUT37), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n887), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n865), .B1(new_n886), .B2(new_n891), .ZN(new_n892));
  AND3_X1   g0692(.A1(new_n727), .A2(KEYINPUT31), .A3(new_n683), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n893), .A2(new_n728), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n738), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n895), .A2(new_n859), .ZN(new_n896));
  INV_X1    g0696(.A(new_n879), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n478), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT38), .B1(new_n898), .B2(new_n882), .ZN(new_n899));
  AOI22_X1  g0699(.A1(new_n869), .A2(new_n873), .B1(new_n880), .B2(KEYINPUT37), .ZN(new_n900));
  AOI211_X1 g0700(.A(new_n887), .B(new_n900), .C1(new_n478), .C2(new_n897), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n896), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT40), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n892), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(new_n662), .B2(new_n895), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n905), .A2(new_n692), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n904), .A2(new_n662), .A3(new_n895), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n882), .B1(new_n885), .B2(new_n879), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n887), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n910), .A2(KEYINPUT39), .A3(new_n886), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n886), .A2(new_n891), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT39), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n375), .A2(new_n683), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n911), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n649), .A2(new_n870), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n910), .A2(new_n886), .ZN(new_n918));
  INV_X1    g0718(.A(new_n820), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n919), .B1(new_n713), .B2(new_n819), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n856), .A2(new_n858), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n917), .B1(new_n918), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n916), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n662), .B1(new_n716), .B2(new_n740), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n661), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n925), .B(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n854), .B1(new_n908), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n928), .B2(new_n908), .ZN(new_n930));
  OR2_X1    g0730(.A1(new_n521), .A2(KEYINPUT35), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n521), .A2(KEYINPUT35), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n931), .A2(G116), .A3(new_n218), .A4(new_n932), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT36), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n216), .A2(new_n247), .A3(new_n422), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(G50), .B2(new_n213), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n936), .A2(G1), .A3(new_n744), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n930), .A2(new_n934), .A3(new_n937), .ZN(G367));
  OAI21_X1  g0738(.A(new_n665), .B1(new_n530), .B2(new_n696), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n580), .B2(new_n696), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n691), .A2(new_n703), .A3(new_n940), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n941), .A2(KEYINPUT42), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n580), .B1(new_n939), .B2(new_n663), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n941), .A2(KEYINPUT42), .B1(new_n696), .B2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT107), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n606), .A2(new_n696), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n945), .B1(new_n947), .B2(new_n612), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n613), .A2(KEYINPUT107), .A3(new_n946), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n948), .B(new_n949), .C1(new_n669), .C2(new_n946), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n942), .A2(new_n944), .B1(KEYINPUT43), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n950), .A2(KEYINPUT43), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n951), .A2(new_n953), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n701), .A2(new_n940), .ZN(new_n956));
  OR3_X1    g0756(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n956), .B1(new_n954), .B2(new_n955), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n707), .B(KEYINPUT41), .Z(new_n959));
  NOR2_X1   g0759(.A1(new_n704), .A2(new_n940), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(KEYINPUT108), .B2(KEYINPUT44), .ZN(new_n961));
  NAND2_X1  g0761(.A1(KEYINPUT108), .A2(KEYINPUT44), .ZN(new_n962));
  NOR2_X1   g0762(.A1(KEYINPUT108), .A2(KEYINPUT44), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n704), .B2(new_n940), .ZN(new_n964));
  AND3_X1   g0764(.A1(new_n961), .A2(new_n962), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n704), .A2(new_n940), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT45), .ZN(new_n967));
  OR3_X1    g0767(.A1(new_n965), .A2(new_n701), .A3(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n691), .A2(new_n703), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT109), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n699), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n813), .B(KEYINPUT109), .C1(new_n691), .C2(new_n703), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n691), .A2(new_n703), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n973), .B(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n701), .B1(new_n965), .B2(new_n967), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n968), .A2(new_n975), .A3(new_n742), .A4(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n959), .B1(new_n977), .B2(new_n742), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n957), .B(new_n958), .C1(new_n978), .C2(new_n747), .ZN(new_n979));
  INV_X1    g0779(.A(new_n387), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n757), .B1(new_n706), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n759), .A2(new_n238), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n749), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n792), .A2(new_n213), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n353), .B1(new_n781), .B2(new_n220), .ZN(new_n985));
  INV_X1    g0785(.A(G137), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n789), .A2(new_n212), .B1(new_n786), .B2(new_n986), .ZN(new_n987));
  NOR3_X1   g0787(.A1(new_n984), .A2(new_n985), .A3(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n839), .B2(new_n436), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n286), .A2(new_n778), .B1(new_n829), .B2(new_n292), .ZN(new_n990));
  AOI211_X1 g0790(.A(new_n989), .B(new_n990), .C1(G143), .C2(new_n775), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n991), .B(KEYINPUT111), .Z(new_n992));
  INV_X1    g0792(.A(KEYINPUT46), .ZN(new_n993));
  NOR3_X1   g0793(.A1(new_n789), .A2(new_n993), .A3(new_n592), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n993), .B1(new_n789), .B2(new_n592), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n516), .B2(new_n792), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n994), .B(new_n996), .C1(new_n769), .C2(G303), .ZN(new_n997));
  INV_X1    g0797(.A(G317), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n250), .B1(new_n786), .B2(new_n998), .C1(new_n781), .C2(new_n518), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n999), .A2(KEYINPUT110), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n775), .A2(G311), .B1(new_n999), .B2(KEYINPUT110), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(G283), .A2(new_n777), .B1(new_n772), .B2(G294), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n997), .A2(new_n1000), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n992), .A2(new_n1003), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT112), .Z(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT47), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n983), .B1(new_n753), .B2(new_n950), .C1(new_n1006), .C2(new_n755), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n979), .A2(new_n1007), .ZN(G387));
  AOI21_X1  g0808(.A(new_n708), .B1(new_n975), .B2(new_n742), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n742), .B2(new_n975), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n709), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n763), .A2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(G107), .B2(new_n209), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n235), .A2(new_n267), .ZN(new_n1014));
  AOI211_X1 g0814(.A(G45), .B(new_n1011), .C1(G68), .C2(G77), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n294), .A2(new_n286), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT50), .Z(new_n1017));
  AOI21_X1  g0817(.A(new_n760), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1013), .B1(new_n1014), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n748), .B1(new_n1019), .B2(new_n758), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n691), .A2(new_n753), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n789), .A2(new_n220), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1022), .A2(new_n250), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1023), .B1(new_n292), .B2(new_n786), .C1(new_n783), .C2(new_n518), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT113), .Z(new_n1025));
  AOI22_X1  g0825(.A1(G68), .A2(new_n777), .B1(new_n772), .B2(new_n294), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT114), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n792), .A2(new_n387), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n829), .A2(new_n286), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n1028), .B(new_n1029), .C1(G159), .C2(new_n775), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1025), .A2(new_n1027), .A3(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n353), .B1(new_n802), .B2(G326), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n792), .A2(new_n838), .B1(new_n789), .B2(new_n844), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(G311), .A2(new_n772), .B1(new_n775), .B2(G322), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1034), .B1(new_n804), .B2(new_n778), .C1(new_n998), .C2(new_n829), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT48), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1033), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n1036), .B2(new_n1035), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT49), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1032), .B1(new_n592), .B2(new_n781), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1031), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  OR2_X1    g0842(.A1(new_n1042), .A2(KEYINPUT115), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n755), .B1(new_n1042), .B2(KEYINPUT115), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1020), .B(new_n1021), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(new_n975), .B2(new_n747), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1010), .A2(new_n1046), .ZN(G393));
  NAND3_X1  g0847(.A1(new_n968), .A2(new_n747), .A3(new_n976), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(G311), .A2(new_n769), .B1(new_n775), .B2(G317), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT52), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n353), .B1(new_n802), .B2(G322), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1051), .B1(new_n838), .B2(new_n789), .C1(new_n592), .C2(new_n792), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n844), .A2(new_n778), .B1(new_n839), .B2(new_n804), .ZN(new_n1053));
  OR4_X1    g0853(.A1(new_n784), .A2(new_n1050), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(G150), .A2(new_n775), .B1(new_n769), .B2(G159), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT51), .Z(new_n1056));
  NOR2_X1   g0856(.A1(new_n792), .A2(new_n327), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n353), .B1(new_n786), .B2(new_n828), .C1(new_n789), .C2(new_n213), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n1057), .B(new_n1058), .C1(new_n782), .C2(G87), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(G50), .A2(new_n772), .B1(new_n777), .B2(new_n294), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1056), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n755), .B1(new_n1054), .B2(new_n1061), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n760), .A2(new_n245), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n757), .B1(G97), .B2(new_n706), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n749), .B(new_n1062), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n940), .B2(new_n753), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1048), .A2(new_n1066), .ZN(new_n1067));
  AND2_X1   g0867(.A1(new_n977), .A2(new_n707), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n968), .A2(new_n976), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n975), .A2(new_n742), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1067), .B1(new_n1068), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(G390));
  INV_X1    g0873(.A(new_n920), .ZN(new_n1074));
  OAI21_X1  g0874(.A(G330), .B1(new_n864), .B2(new_n860), .ZN(new_n1075));
  NOR3_X1   g0875(.A1(new_n1075), .A2(new_n922), .A3(new_n821), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n921), .B1(new_n739), .B2(new_n822), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1074), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n922), .B1(new_n1075), .B2(new_n821), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n739), .A2(new_n859), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1079), .A2(new_n920), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1078), .A2(new_n1081), .ZN(new_n1082));
  OR2_X1    g0882(.A1(new_n657), .A2(new_n659), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n662), .A2(G330), .A3(new_n895), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1083), .A2(new_n926), .A3(new_n1084), .A4(new_n645), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1082), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n915), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n920), .B2(new_n922), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n911), .A2(new_n914), .A3(new_n1089), .ZN(new_n1090));
  AND2_X1   g0890(.A1(new_n886), .A2(new_n891), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1091), .B(new_n1088), .C1(new_n922), .C2(new_n920), .ZN(new_n1092));
  AND3_X1   g0892(.A1(new_n1090), .A2(new_n1092), .A3(new_n1076), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n1090), .A2(new_n1092), .B1(new_n739), .B2(new_n859), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1087), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n1080), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1090), .A2(new_n1092), .A3(new_n1076), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1085), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1097), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1095), .A2(new_n1100), .A3(new_n707), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n848), .ZN(new_n1102));
  INV_X1    g0902(.A(G128), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n1103), .A2(new_n776), .B1(new_n839), .B2(new_n986), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(KEYINPUT54), .B(G143), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n834), .A2(new_n829), .B1(new_n778), .B2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n789), .A2(new_n292), .ZN(new_n1107));
  XOR2_X1   g0907(.A(new_n1107), .B(KEYINPUT53), .Z(new_n1108));
  INV_X1    g0908(.A(new_n781), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n250), .B1(new_n1109), .B2(G50), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n802), .A2(G125), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1110), .B(new_n1111), .C1(new_n436), .C2(new_n792), .ZN(new_n1112));
  NOR4_X1   g0912(.A1(new_n1104), .A2(new_n1106), .A3(new_n1108), .A4(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT116), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(G107), .A2(new_n772), .B1(new_n775), .B2(G283), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n1115), .B1(new_n518), .B2(new_n778), .C1(new_n592), .C2(new_n829), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n250), .B1(new_n786), .B2(new_n844), .C1(new_n789), .C2(new_n413), .ZN(new_n1117));
  NOR4_X1   g0917(.A1(new_n1116), .A2(new_n832), .A3(new_n1057), .A4(new_n1117), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1114), .A2(new_n1118), .ZN(new_n1119));
  AND2_X1   g0919(.A1(new_n1119), .A2(KEYINPUT117), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n754), .B1(new_n1119), .B2(KEYINPUT117), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n748), .B1(new_n294), .B2(new_n1102), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n911), .A2(new_n914), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1122), .B1(new_n1123), .B2(new_n750), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1124), .B1(new_n1125), .B2(new_n747), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1101), .A2(new_n1126), .ZN(G378));
  NAND2_X1  g0927(.A1(new_n1100), .A2(new_n1086), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(KEYINPUT57), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n310), .A2(new_n681), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1130), .B(KEYINPUT55), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  OR2_X1    g0932(.A1(new_n323), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n323), .A2(new_n1132), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  XOR2_X1   g0935(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1133), .A2(new_n1136), .A3(new_n1134), .ZN(new_n1139));
  AND2_X1   g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(new_n904), .B2(G330), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n865), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(new_n912), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n895), .A2(new_n859), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(new_n910), .B2(new_n886), .ZN(new_n1145));
  OAI211_X1 g0945(.A(G330), .B(new_n1143), .C1(new_n1145), .C2(KEYINPUT40), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1140), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n925), .B1(new_n1141), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n916), .A2(new_n924), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n902), .A2(new_n903), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1152), .A2(G330), .A3(new_n1143), .A4(new_n1140), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1150), .A2(new_n1151), .A3(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1149), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT120), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1154), .A2(KEYINPUT120), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1129), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n1149), .A2(new_n1154), .B1(new_n1100), .B2(new_n1086), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n707), .B1(new_n1160), .B2(KEYINPUT57), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n746), .B1(new_n1149), .B2(new_n1154), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n792), .A2(new_n292), .B1(new_n1105), .B2(new_n789), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n775), .A2(G125), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n1164), .B1(new_n829), .B2(new_n1103), .C1(new_n986), .C2(new_n778), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n1163), .B(new_n1165), .C1(G132), .C2(new_n772), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT59), .ZN(new_n1167));
  OR2_X1    g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1109), .A2(G159), .ZN(new_n1170));
  AOI211_X1 g0970(.A(G33), .B(G41), .C1(new_n802), .C2(G124), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .A4(new_n1171), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n516), .A2(new_n829), .B1(new_n778), .B2(new_n387), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n781), .A2(new_n212), .B1(new_n838), .B2(new_n786), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n250), .A2(new_n266), .ZN(new_n1175));
  NOR4_X1   g0975(.A1(new_n984), .A2(new_n1174), .A3(new_n1022), .A4(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n839), .B2(new_n518), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1173), .B(new_n1177), .C1(G116), .C2(new_n775), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(KEYINPUT58), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1175), .B(new_n286), .C1(G33), .C2(G41), .ZN(new_n1180));
  OR2_X1    g0980(.A1(new_n1178), .A2(KEYINPUT58), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1172), .A2(new_n1179), .A3(new_n1180), .A4(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(new_n754), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n749), .B1(new_n286), .B2(new_n848), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1183), .B(new_n1184), .C1(new_n1140), .C2(new_n751), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NOR3_X1   g0986(.A1(new_n1162), .A2(KEYINPUT119), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT119), .ZN(new_n1188));
  AND3_X1   g0988(.A1(new_n1150), .A2(new_n1151), .A3(new_n1153), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n1150), .A2(new_n1153), .B1(new_n916), .B2(new_n924), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n747), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1188), .B1(new_n1191), .B2(new_n1185), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n1159), .A2(new_n1161), .B1(new_n1187), .B2(new_n1192), .ZN(G375));
  NAND3_X1  g0993(.A1(new_n1085), .A2(new_n1078), .A3(new_n1081), .ZN(new_n1194));
  XOR2_X1   g0994(.A(new_n959), .B(KEYINPUT121), .Z(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1087), .A2(new_n1194), .A3(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1082), .A2(new_n747), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n748), .B1(G68), .B2(new_n1102), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(G107), .A2(new_n777), .B1(new_n772), .B2(G116), .ZN(new_n1200));
  XOR2_X1   g1000(.A(new_n1200), .B(KEYINPUT122), .Z(new_n1201));
  OAI221_X1 g1001(.A(new_n250), .B1(new_n786), .B2(new_n804), .C1(new_n789), .C2(new_n518), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1028), .B(new_n1202), .C1(new_n782), .C2(G77), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(G283), .A2(new_n769), .B1(new_n775), .B2(G294), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1201), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n777), .A2(G150), .B1(G50), .B2(new_n791), .ZN(new_n1206));
  XOR2_X1   g1006(.A(new_n1206), .B(KEYINPUT124), .Z(new_n1207));
  OAI21_X1  g1007(.A(new_n353), .B1(new_n781), .B2(new_n212), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n789), .A2(new_n436), .B1(new_n786), .B2(new_n1103), .ZN(new_n1209));
  OR3_X1    g1009(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(G132), .A2(new_n775), .B1(new_n769), .B2(G137), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1211), .B1(new_n839), .B2(new_n1105), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1212), .B(KEYINPUT123), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1205), .B1(new_n1210), .B2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1199), .B1(new_n1214), .B2(new_n754), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n751), .B2(new_n921), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1197), .A2(new_n1198), .A3(new_n1216), .ZN(G381));
  INV_X1    g1017(.A(KEYINPUT57), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n1100), .B2(new_n1086), .ZN(new_n1219));
  AOI21_X1  g1019(.A(KEYINPUT120), .B1(new_n1149), .B2(new_n1154), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1158), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1219), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1085), .B1(new_n1125), .B2(new_n1082), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1218), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1222), .A2(new_n707), .A3(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(G378), .ZN(new_n1227));
  OAI21_X1  g1027(.A(KEYINPUT119), .B1(new_n1162), .B2(new_n1186), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1191), .A2(new_n1188), .A3(new_n1185), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n1226), .A2(new_n1227), .A3(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n979), .A2(new_n1072), .A3(new_n1007), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  NOR4_X1   g1033(.A1(G393), .A2(G384), .A3(G396), .A4(G381), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1231), .A2(new_n1233), .A3(new_n1234), .ZN(G407));
  NAND3_X1  g1035(.A1(new_n1226), .A2(new_n1230), .A3(new_n1227), .ZN(new_n1236));
  INV_X1    g1036(.A(G213), .ZN(new_n1237));
  OR3_X1    g1037(.A1(new_n1237), .A2(KEYINPUT125), .A3(G343), .ZN(new_n1238));
  OAI21_X1  g1038(.A(KEYINPUT125), .B1(new_n1237), .B2(G343), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  OAI211_X1 g1040(.A(G407), .B(G213), .C1(new_n1236), .C2(new_n1240), .ZN(G409));
  INV_X1    g1041(.A(new_n1240), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1101), .A2(new_n1126), .A3(new_n1185), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(new_n1160), .B2(new_n1196), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n747), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1242), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1155), .A2(new_n1128), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n708), .B1(new_n1247), .B2(new_n1218), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n1248), .A2(new_n1222), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1246), .B1(new_n1227), .B2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1198), .A2(new_n1216), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1194), .B(KEYINPUT60), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1099), .A2(new_n708), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1251), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1254), .A2(new_n852), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1254), .A2(new_n852), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1242), .A2(G2897), .ZN(new_n1258));
  XOR2_X1   g1058(.A(new_n1258), .B(KEYINPUT126), .Z(new_n1259));
  NAND3_X1  g1059(.A1(new_n1256), .A2(new_n1257), .A3(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1257), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1261), .A2(new_n1255), .ZN(new_n1262));
  OR2_X1    g1062(.A1(new_n1258), .A2(KEYINPUT126), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1260), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(KEYINPUT61), .B1(new_n1250), .B2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(G375), .A2(G378), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1262), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1266), .A2(new_n1267), .A3(new_n1246), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(KEYINPUT62), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT62), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1266), .A2(new_n1270), .A3(new_n1267), .A4(new_n1246), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1265), .A2(new_n1269), .A3(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1072), .B1(new_n979), .B2(new_n1007), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(G393), .A2(G396), .ZN(new_n1274));
  AND2_X1   g1074(.A1(G393), .A2(G396), .ZN(new_n1275));
  OAI22_X1  g1075(.A1(new_n1233), .A2(new_n1273), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1273), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1275), .A2(new_n1274), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1277), .A2(new_n1278), .A3(new_n1232), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1276), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1272), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT63), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1268), .A2(new_n1283), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1266), .A2(KEYINPUT63), .A3(new_n1267), .A4(new_n1246), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1280), .A2(new_n1265), .A3(new_n1284), .A4(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1282), .A2(new_n1286), .ZN(G405));
  AOI21_X1  g1087(.A(new_n1227), .B1(new_n1226), .B2(new_n1230), .ZN(new_n1288));
  OAI21_X1  g1088(.A(KEYINPUT127), .B1(new_n1231), .B2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT127), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1266), .A2(new_n1290), .A3(new_n1236), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1289), .A2(new_n1291), .A3(new_n1267), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1266), .A2(new_n1290), .A3(new_n1236), .A4(new_n1262), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n1280), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1281), .A2(new_n1292), .A3(new_n1293), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(G402));
endmodule


