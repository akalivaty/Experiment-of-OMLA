//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 0 0 0 0 0 0 1 1 1 1 0 1 1 0 0 1 1 0 0 1 1 1 1 1 1 0 0 0 1 1 1 1 1 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:49 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n770, new_n771,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041;
  AND2_X1   g000(.A1(KEYINPUT72), .A2(G953), .ZN(new_n187));
  NOR2_X1   g001(.A1(KEYINPUT72), .A2(G953), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT22), .B(G137), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n190), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT23), .ZN(new_n194));
  INV_X1    g008(.A(G119), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n194), .B1(new_n195), .B2(G128), .ZN(new_n196));
  INV_X1    g010(.A(G128), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(KEYINPUT23), .A3(G119), .ZN(new_n198));
  OAI211_X1 g012(.A(new_n196), .B(new_n198), .C1(G119), .C2(new_n197), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G110), .ZN(new_n200));
  XNOR2_X1  g014(.A(KEYINPUT24), .B(G110), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT78), .ZN(new_n202));
  OR2_X1    g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n202), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g019(.A(G119), .B(G128), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n200), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT16), .ZN(new_n209));
  INV_X1    g023(.A(G140), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(G125), .ZN(new_n211));
  INV_X1    g025(.A(G125), .ZN(new_n212));
  OR2_X1    g026(.A1(KEYINPUT79), .A2(G140), .ZN(new_n213));
  NAND2_X1  g027(.A1(KEYINPUT79), .A2(G140), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT80), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n211), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  AND2_X1   g031(.A1(KEYINPUT79), .A2(G140), .ZN(new_n218));
  NOR2_X1   g032(.A1(KEYINPUT79), .A2(G140), .ZN(new_n219));
  OAI21_X1  g033(.A(G125), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT80), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n209), .B1(new_n217), .B2(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(KEYINPUT16), .B1(new_n210), .B2(G125), .ZN(new_n223));
  OAI21_X1  g037(.A(G146), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n211), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n216), .B(G125), .C1(new_n218), .C2(new_n219), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n221), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(KEYINPUT16), .ZN(new_n228));
  INV_X1    g042(.A(G146), .ZN(new_n229));
  INV_X1    g043(.A(new_n223), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n208), .B1(new_n224), .B2(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n223), .B1(new_n227), .B2(KEYINPUT16), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n233), .A2(new_n229), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n210), .A2(G125), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n225), .A2(new_n235), .A3(new_n229), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n206), .B1(new_n203), .B2(new_n204), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n199), .A2(G110), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n234), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n193), .B1(new_n232), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n208), .ZN(new_n242));
  NOR3_X1   g056(.A1(new_n222), .A2(G146), .A3(new_n223), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n242), .B1(new_n234), .B2(new_n243), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n224), .B(new_n236), .C1(new_n238), .C2(new_n237), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n244), .A2(new_n245), .A3(new_n192), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n241), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT76), .B(G217), .ZN(new_n248));
  INV_X1    g062(.A(G902), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n248), .B1(G234), .B2(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n250), .A2(G902), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n241), .A2(new_n246), .A3(new_n249), .ZN(new_n253));
  NAND2_X1  g067(.A1(KEYINPUT82), .A2(KEYINPUT25), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT81), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  XOR2_X1   g071(.A(new_n250), .B(KEYINPUT77), .Z(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n241), .A2(new_n246), .A3(new_n255), .A4(new_n249), .ZN(new_n261));
  AOI21_X1  g075(.A(KEYINPUT25), .B1(new_n261), .B2(KEYINPUT82), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n252), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  NOR2_X1   g077(.A1(G472), .A2(G902), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT71), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n266), .B1(new_n195), .B2(G116), .ZN(new_n267));
  INV_X1    g081(.A(G116), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n268), .A2(KEYINPUT70), .A3(G119), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n195), .A2(G116), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT2), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n273), .A2(G113), .ZN(new_n274));
  INV_X1    g088(.A(G113), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n275), .A2(KEYINPUT2), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n272), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n265), .B1(new_n271), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n275), .A2(KEYINPUT2), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n273), .A2(G113), .ZN(new_n280));
  AOI22_X1  g094(.A1(new_n279), .A2(new_n280), .B1(G116), .B2(new_n195), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n281), .A2(KEYINPUT71), .A3(new_n270), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n270), .A2(new_n272), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n274), .A2(new_n276), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n278), .A2(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(KEYINPUT64), .B1(new_n229), .B2(G143), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT64), .ZN(new_n287));
  INV_X1    g101(.A(G143), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n287), .A2(new_n288), .A3(G146), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n288), .A2(G146), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT65), .ZN(new_n294));
  XNOR2_X1  g108(.A(KEYINPUT0), .B(G128), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n293), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT11), .ZN(new_n298));
  INV_X1    g112(.A(G134), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n298), .B1(new_n299), .B2(G137), .ZN(new_n300));
  INV_X1    g114(.A(G137), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n301), .A2(KEYINPUT11), .A3(G134), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n299), .A2(G137), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n300), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G131), .ZN(new_n305));
  INV_X1    g119(.A(G131), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n300), .A2(new_n302), .A3(new_n306), .A4(new_n303), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n291), .B1(new_n286), .B2(new_n289), .ZN(new_n309));
  OAI21_X1  g123(.A(KEYINPUT65), .B1(new_n309), .B2(new_n295), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT66), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n311), .B1(new_n288), .B2(G146), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n229), .A2(KEYINPUT66), .A3(G143), .ZN(new_n313));
  AOI22_X1  g127(.A1(new_n312), .A2(new_n313), .B1(new_n288), .B2(G146), .ZN(new_n314));
  AND2_X1   g128(.A1(KEYINPUT0), .A2(G128), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n297), .A2(new_n308), .A3(new_n310), .A4(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n288), .A2(G146), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n229), .A2(KEYINPUT66), .A3(G143), .ZN(new_n319));
  AOI21_X1  g133(.A(KEYINPUT66), .B1(new_n229), .B2(G143), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  XNOR2_X1  g135(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G128), .ZN(new_n323));
  OAI21_X1  g137(.A(KEYINPUT69), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT1), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT68), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT68), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(KEYINPUT1), .ZN(new_n328));
  AND3_X1   g142(.A1(new_n326), .A2(new_n328), .A3(G128), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT69), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n314), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(G128), .B1(new_n322), .B2(new_n291), .ZN(new_n332));
  AOI22_X1  g146(.A1(new_n324), .A2(new_n331), .B1(new_n332), .B2(new_n293), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT67), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n334), .B1(new_n299), .B2(G137), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n301), .A2(KEYINPUT67), .A3(G134), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n335), .A2(new_n303), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G131), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n307), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n285), .B(new_n317), .C1(new_n333), .C2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n332), .A2(new_n293), .ZN(new_n342));
  AND3_X1   g156(.A1(new_n314), .A2(new_n330), .A3(new_n329), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n330), .B1(new_n314), .B2(new_n329), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n339), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n285), .B1(new_n347), .B2(new_n317), .ZN(new_n348));
  OAI21_X1  g162(.A(KEYINPUT28), .B1(new_n341), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT28), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n340), .A2(KEYINPUT74), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(KEYINPUT74), .B1(new_n340), .B2(new_n350), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n349), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G237), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n189), .A2(G210), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(KEYINPUT27), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT27), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n189), .A2(new_n358), .A3(G210), .A4(new_n355), .ZN(new_n359));
  XNOR2_X1  g173(.A(KEYINPUT26), .B(G101), .ZN(new_n360));
  AND3_X1   g174(.A1(new_n357), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n360), .B1(new_n357), .B2(new_n359), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n354), .A2(KEYINPUT75), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n324), .A2(new_n331), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n339), .B1(new_n366), .B2(new_n342), .ZN(new_n367));
  AND4_X1   g181(.A1(new_n308), .A2(new_n297), .A3(new_n310), .A4(new_n316), .ZN(new_n368));
  OAI21_X1  g182(.A(KEYINPUT30), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT30), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n370), .B(new_n317), .C1(new_n333), .C2(new_n339), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n285), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT73), .ZN(new_n373));
  AND3_X1   g187(.A1(new_n340), .A2(new_n373), .A3(new_n363), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n373), .B1(new_n340), .B2(new_n363), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(KEYINPUT31), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT31), .ZN(new_n379));
  NOR4_X1   g193(.A1(new_n372), .A2(new_n374), .A3(new_n376), .A4(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n365), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT75), .ZN(new_n382));
  INV_X1    g196(.A(new_n285), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n383), .B1(new_n367), .B2(new_n368), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n350), .B1(new_n384), .B2(new_n340), .ZN(new_n385));
  AND3_X1   g199(.A1(new_n340), .A2(KEYINPUT74), .A3(new_n350), .ZN(new_n386));
  NOR3_X1   g200(.A1(new_n385), .A2(new_n386), .A3(new_n352), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n382), .B1(new_n387), .B2(new_n363), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n264), .B1(new_n381), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT32), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n371), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n370), .B1(new_n347), .B2(new_n317), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n383), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n340), .A2(new_n373), .A3(new_n363), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n395), .A2(new_n377), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n379), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n375), .A2(KEYINPUT31), .A3(new_n377), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n400), .A2(new_n388), .A3(new_n365), .ZN(new_n401));
  INV_X1    g215(.A(new_n264), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n402), .A2(new_n391), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n385), .A2(new_n352), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n404), .A2(KEYINPUT29), .A3(new_n363), .A4(new_n351), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n364), .B1(new_n372), .B2(new_n341), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT29), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NOR4_X1   g222(.A1(new_n385), .A2(new_n386), .A3(new_n352), .A4(new_n364), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n405), .B(new_n249), .C1(new_n408), .C2(new_n409), .ZN(new_n410));
  AOI22_X1  g224(.A1(new_n401), .A2(new_n403), .B1(new_n410), .B2(G472), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n263), .B1(new_n392), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(G214), .B1(G237), .B2(G902), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(G475), .A2(G902), .ZN(new_n415));
  OR2_X1    g229(.A1(KEYINPUT72), .A2(G953), .ZN(new_n416));
  NAND2_X1  g230(.A1(KEYINPUT72), .A2(G953), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n416), .A2(G214), .A3(new_n355), .A4(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(KEYINPUT89), .B(G143), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  OR2_X1    g234(.A1(KEYINPUT89), .A2(G143), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n189), .A2(G214), .A3(new_n355), .A4(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(G131), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT17), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n420), .A2(new_n422), .A3(new_n306), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n306), .B1(new_n420), .B2(new_n422), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(KEYINPUT17), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n224), .A2(new_n427), .A3(new_n231), .A4(new_n429), .ZN(new_n430));
  XNOR2_X1  g244(.A(G113), .B(G122), .ZN(new_n431));
  INV_X1    g245(.A(G104), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n431), .B(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n227), .A2(G146), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n236), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n428), .A2(KEYINPUT18), .ZN(new_n436));
  NAND2_X1  g250(.A1(KEYINPUT18), .A2(G131), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n420), .A2(new_n422), .A3(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n435), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  AND3_X1   g253(.A1(new_n430), .A2(new_n433), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n424), .A2(new_n426), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n227), .A2(KEYINPUT19), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n225), .A2(new_n235), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n442), .B1(KEYINPUT19), .B2(new_n443), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n224), .B(new_n441), .C1(new_n444), .C2(G146), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n433), .B1(new_n445), .B2(new_n439), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n415), .B1(new_n440), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(KEYINPUT20), .ZN(new_n448));
  AND3_X1   g262(.A1(new_n420), .A2(new_n422), .A3(new_n306), .ZN(new_n449));
  OAI22_X1  g263(.A1(new_n233), .A2(new_n229), .B1(new_n428), .B2(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n443), .A2(KEYINPUT19), .ZN(new_n451));
  AOI211_X1 g265(.A(G146), .B(new_n451), .C1(new_n227), .C2(KEYINPUT19), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n439), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n433), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n430), .A2(new_n433), .A3(new_n439), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT20), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n457), .A2(new_n458), .A3(new_n415), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n448), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(G234), .A2(G237), .ZN(new_n461));
  INV_X1    g275(.A(G953), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n461), .A2(G952), .A3(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n463), .B(KEYINPUT93), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n189), .ZN(new_n466));
  AND3_X1   g280(.A1(new_n466), .A2(G902), .A3(new_n461), .ZN(new_n467));
  XNOR2_X1  g281(.A(KEYINPUT21), .B(G898), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n433), .B1(new_n430), .B2(new_n439), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n249), .B1(new_n440), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(G475), .ZN(new_n473));
  INV_X1    g287(.A(G478), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n474), .A2(KEYINPUT15), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n288), .A2(KEYINPUT13), .A3(G128), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(KEYINPUT90), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n288), .A2(G128), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT13), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT90), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n481), .A2(new_n288), .A3(KEYINPUT13), .A4(G128), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n197), .A2(G143), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n477), .A2(new_n480), .A3(new_n482), .A4(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(G134), .ZN(new_n485));
  XNOR2_X1  g299(.A(G116), .B(G122), .ZN(new_n486));
  INV_X1    g300(.A(G107), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n486), .B(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n478), .A2(new_n483), .A3(new_n299), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n485), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n268), .A2(KEYINPUT14), .A3(G122), .ZN(new_n491));
  INV_X1    g305(.A(new_n486), .ZN(new_n492));
  OAI211_X1 g306(.A(G107), .B(new_n491), .C1(new_n492), .C2(KEYINPUT14), .ZN(new_n493));
  OAI21_X1  g307(.A(KEYINPUT91), .B1(new_n492), .B2(G107), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n478), .A2(new_n483), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(G134), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n489), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT91), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n486), .A2(new_n498), .A3(new_n487), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n493), .A2(new_n494), .A3(new_n497), .A4(new_n499), .ZN(new_n500));
  XNOR2_X1  g314(.A(KEYINPUT9), .B(G234), .ZN(new_n501));
  NOR3_X1   g315(.A1(new_n248), .A2(new_n501), .A3(G953), .ZN(new_n502));
  AND3_X1   g316(.A1(new_n490), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n502), .B1(new_n490), .B2(new_n500), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n249), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT92), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n475), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n505), .A2(new_n506), .ZN(new_n508));
  OAI211_X1 g322(.A(KEYINPUT92), .B(new_n249), .C1(new_n503), .C2(new_n504), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n507), .B1(new_n510), .B2(new_n475), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n460), .A2(new_n470), .A3(new_n473), .A4(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n270), .A2(KEYINPUT5), .A3(new_n272), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n272), .A2(KEYINPUT5), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n514), .A2(new_n275), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(G101), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n487), .A2(G104), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n432), .A2(G107), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n487), .A2(KEYINPUT83), .A3(G104), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT3), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n487), .A2(KEYINPUT83), .A3(KEYINPUT3), .A4(G104), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n519), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n526), .A2(G101), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n520), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n281), .A2(KEYINPUT71), .A3(new_n270), .ZN(new_n529));
  AOI21_X1  g343(.A(KEYINPUT71), .B1(new_n281), .B2(new_n270), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n516), .B(new_n528), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n432), .A2(G107), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT3), .B1(new_n532), .B2(KEYINPUT83), .ZN(new_n533));
  INV_X1    g347(.A(new_n524), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n519), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT4), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n535), .A2(new_n536), .A3(G101), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n525), .A2(new_n527), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(KEYINPUT4), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n526), .B1(new_n523), .B2(new_n524), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n540), .A2(new_n517), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n537), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n531), .B1(new_n542), .B2(new_n285), .ZN(new_n543));
  XNOR2_X1  g357(.A(G110), .B(G122), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n531), .B(new_n544), .C1(new_n542), .C2(new_n285), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(KEYINPUT6), .A3(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT6), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n543), .A2(new_n549), .A3(new_n545), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n297), .A2(new_n310), .A3(new_n316), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(G125), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n212), .B(new_n342), .C1(new_n343), .C2(new_n344), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(G224), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n555), .A2(G953), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n556), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n552), .A2(new_n553), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n548), .A2(new_n550), .A3(new_n560), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n561), .A2(new_n249), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT7), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n556), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n552), .A2(new_n553), .A3(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n564), .B1(new_n552), .B2(new_n553), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n531), .A2(KEYINPUT86), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n278), .A2(new_n282), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n528), .B1(new_n570), .B2(new_n516), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n516), .B1(new_n529), .B2(new_n530), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT86), .ZN(new_n574));
  INV_X1    g388(.A(new_n528), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n544), .B(KEYINPUT8), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT87), .ZN(new_n579));
  NOR3_X1   g393(.A1(new_n572), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n577), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n581), .B1(new_n571), .B2(new_n574), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n573), .A2(new_n575), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n583), .A2(KEYINPUT86), .A3(new_n531), .ZN(new_n584));
  AOI21_X1  g398(.A(KEYINPUT87), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  OAI211_X1 g399(.A(KEYINPUT88), .B(new_n568), .C1(new_n580), .C2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n547), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n579), .B1(new_n572), .B2(new_n578), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n582), .A2(KEYINPUT87), .A3(new_n584), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(KEYINPUT88), .B1(new_n590), .B2(new_n568), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n562), .B1(new_n587), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(G210), .B1(G237), .B2(G902), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n547), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n558), .A2(KEYINPUT7), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n554), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n565), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n599), .B1(new_n588), .B2(new_n589), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n596), .B1(new_n600), .B2(KEYINPUT88), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n590), .A2(new_n568), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT88), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n605), .A2(new_n562), .A3(new_n593), .ZN(new_n606));
  AOI211_X1 g420(.A(new_n414), .B(new_n512), .C1(new_n595), .C2(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(G221), .B1(new_n501), .B2(G902), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(G469), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n189), .A2(G227), .ZN(new_n611));
  XOR2_X1   g425(.A(G110), .B(G140), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g428(.A(KEYINPUT10), .B1(new_n333), .B2(new_n575), .ZN(new_n615));
  OAI21_X1  g429(.A(G128), .B1(new_n291), .B2(new_n325), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n321), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n617), .B1(new_n343), .B2(new_n344), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT10), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n618), .A2(new_n619), .A3(new_n528), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n615), .A2(new_n620), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n540), .A2(KEYINPUT4), .A3(new_n517), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n535), .A2(G101), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n536), .B1(new_n525), .B2(new_n527), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n297), .A2(new_n310), .A3(new_n316), .ZN(new_n626));
  AOI21_X1  g440(.A(KEYINPUT84), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT84), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n542), .A2(new_n628), .A3(new_n551), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n621), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT85), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n630), .A2(new_n631), .A3(new_n308), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n628), .B1(new_n542), .B2(new_n551), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n623), .A2(new_n624), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n626), .A2(KEYINPUT84), .A3(new_n634), .A4(new_n537), .ZN(new_n635));
  AOI22_X1  g449(.A1(new_n633), .A2(new_n635), .B1(new_n615), .B2(new_n620), .ZN(new_n636));
  INV_X1    g450(.A(new_n308), .ZN(new_n637));
  OAI21_X1  g451(.A(KEYINPUT85), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n632), .A2(new_n638), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n621), .B(new_n637), .C1(new_n627), .C2(new_n629), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n614), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n618), .A2(new_n528), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n642), .B1(new_n345), .B2(new_n528), .ZN(new_n643));
  AND3_X1   g457(.A1(new_n643), .A2(KEYINPUT12), .A3(new_n308), .ZN(new_n644));
  AOI21_X1  g458(.A(KEYINPUT12), .B1(new_n643), .B2(new_n308), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n640), .A2(new_n614), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  OAI211_X1 g462(.A(new_n610), .B(new_n249), .C1(new_n641), .C2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n647), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n640), .B1(new_n644), .B2(new_n645), .ZN(new_n651));
  AOI22_X1  g465(.A1(new_n639), .A2(new_n650), .B1(new_n651), .B2(new_n613), .ZN(new_n652));
  OAI21_X1  g466(.A(G469), .B1(new_n652), .B2(G902), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n609), .B1(new_n649), .B2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n412), .A2(new_n607), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G101), .ZN(G3));
  AOI211_X1 g470(.A(new_n263), .B(new_n609), .C1(new_n649), .C2(new_n653), .ZN(new_n657));
  AOI211_X1 g471(.A(new_n414), .B(new_n469), .C1(new_n595), .C2(new_n606), .ZN(new_n658));
  INV_X1    g472(.A(G472), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n659), .B1(new_n401), .B2(new_n249), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n363), .B1(new_n404), .B2(new_n351), .ZN(new_n661));
  AOI22_X1  g475(.A1(KEYINPUT75), .A2(new_n661), .B1(new_n398), .B2(new_n399), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n402), .B1(new_n662), .B2(new_n388), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  AND3_X1   g478(.A1(new_n657), .A2(new_n658), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n460), .A2(new_n473), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n503), .A2(new_n504), .ZN(new_n667));
  OAI21_X1  g481(.A(KEYINPUT33), .B1(new_n502), .B2(KEYINPUT94), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n669), .A2(G478), .A3(new_n249), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT95), .B(G478), .Z(new_n671));
  NAND2_X1  g485(.A1(new_n505), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n666), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(new_n674), .B(KEYINPUT96), .Z(new_n675));
  NAND2_X1  g489(.A1(new_n665), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT34), .B(G104), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G6));
  INV_X1    g492(.A(new_n666), .ZN(new_n679));
  INV_X1    g493(.A(new_n511), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n665), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(KEYINPUT35), .B(G107), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(KEYINPUT97), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n683), .B(new_n685), .ZN(G9));
  NAND2_X1  g500(.A1(new_n244), .A2(new_n245), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n193), .A2(KEYINPUT36), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n251), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n690), .B1(new_n260), .B2(new_n262), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n660), .A2(new_n663), .A3(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n693), .A2(new_n607), .A3(new_n654), .ZN(new_n694));
  XOR2_X1   g508(.A(KEYINPUT37), .B(G110), .Z(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT98), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n694), .B(new_n696), .ZN(G12));
  AOI21_X1  g511(.A(new_n692), .B1(new_n392), .B2(new_n411), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n414), .B1(new_n595), .B2(new_n606), .ZN(new_n699));
  INV_X1    g513(.A(new_n467), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n464), .B1(new_n700), .B2(G900), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n681), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n698), .A2(new_n654), .A3(new_n699), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G128), .ZN(G30));
  XNOR2_X1  g519(.A(KEYINPUT101), .B(KEYINPUT39), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n701), .B(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n654), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(KEYINPUT102), .ZN(new_n710));
  OR2_X1    g524(.A1(new_n710), .A2(KEYINPUT40), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(KEYINPUT40), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n595), .A2(new_n606), .ZN(new_n713));
  XOR2_X1   g527(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(KEYINPUT100), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n713), .B(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n401), .A2(new_n403), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n364), .B1(new_n341), .B2(new_n348), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n397), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g533(.A(G472), .B1(new_n719), .B2(G902), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n392), .A2(new_n717), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n511), .B1(new_n460), .B2(new_n473), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n723), .A2(new_n414), .A3(new_n691), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n716), .A2(new_n721), .A3(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n711), .A2(new_n712), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G143), .ZN(G45));
  NOR2_X1   g541(.A1(new_n674), .A2(new_n702), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n698), .A2(new_n654), .A3(new_n699), .A4(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G146), .ZN(G48));
  AOI21_X1  g544(.A(new_n631), .B1(new_n630), .B2(new_n308), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n636), .A2(KEYINPUT85), .A3(new_n637), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n640), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n648), .B1(new_n733), .B2(new_n613), .ZN(new_n734));
  OAI21_X1  g548(.A(G469), .B1(new_n734), .B2(G902), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n735), .A2(new_n608), .A3(new_n649), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT103), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(new_n738));
  AND2_X1   g552(.A1(new_n412), .A2(new_n658), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n738), .A2(new_n739), .A3(new_n675), .ZN(new_n740));
  XNOR2_X1  g554(.A(KEYINPUT41), .B(G113), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G15));
  NAND3_X1  g556(.A1(new_n738), .A2(new_n739), .A3(new_n682), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G116), .ZN(G18));
  INV_X1    g558(.A(KEYINPUT104), .ZN(new_n745));
  INV_X1    g559(.A(new_n512), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n410), .A2(G472), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n717), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(KEYINPUT32), .B1(new_n401), .B2(new_n264), .ZN(new_n749));
  OAI211_X1 g563(.A(new_n746), .B(new_n691), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n699), .A2(new_n608), .A3(new_n649), .A4(new_n735), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n745), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n592), .A2(new_n594), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n593), .B1(new_n605), .B2(new_n562), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n413), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n736), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n756), .A2(KEYINPUT104), .A3(new_n746), .A4(new_n698), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n752), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G119), .ZN(G21));
  OAI21_X1  g573(.A(KEYINPUT105), .B1(new_n755), .B2(new_n723), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT105), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n699), .A2(new_n761), .A3(new_n722), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n661), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n402), .B1(new_n400), .B2(new_n764), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n660), .A2(new_n263), .A3(new_n765), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n766), .A2(new_n470), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n738), .A2(new_n763), .A3(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G122), .ZN(G24));
  NOR3_X1   g583(.A1(new_n660), .A2(new_n692), .A3(new_n765), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n756), .A2(new_n728), .A3(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G125), .ZN(G27));
  NOR2_X1   g586(.A1(new_n713), .A2(new_n414), .ZN(new_n773));
  NOR2_X1   g587(.A1(KEYINPUT106), .A2(KEYINPUT42), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n674), .A2(new_n702), .A3(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n412), .A2(new_n654), .A3(new_n773), .A4(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(KEYINPUT106), .A2(KEYINPUT42), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n753), .A2(new_n754), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n654), .A2(new_n780), .A3(new_n413), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n781), .A2(new_n412), .A3(new_n775), .A4(new_n777), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(new_n306), .ZN(G33));
  NAND4_X1  g598(.A1(new_n412), .A2(new_n654), .A3(new_n703), .A4(new_n773), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G134), .ZN(G36));
  OR2_X1    g600(.A1(new_n652), .A2(KEYINPUT45), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n652), .A2(KEYINPUT45), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n787), .A2(G469), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(G469), .A2(G902), .ZN(new_n790));
  AOI21_X1  g604(.A(KEYINPUT46), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n649), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n789), .A2(KEYINPUT46), .A3(new_n790), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n609), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n708), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n679), .A2(new_n673), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT43), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n691), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT44), .ZN(new_n802));
  OR3_X1    g616(.A1(new_n801), .A2(new_n802), .A3(new_n664), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n802), .B1(new_n801), .B2(new_n664), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n797), .A2(new_n773), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(KEYINPUT107), .B(G137), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n805), .B(new_n806), .ZN(G39));
  NAND3_X1  g621(.A1(new_n773), .A2(new_n263), .A3(new_n728), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n808), .A2(new_n749), .A3(new_n748), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n795), .A2(KEYINPUT47), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n795), .A2(KEYINPUT47), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G140), .ZN(G42));
  INV_X1    g627(.A(KEYINPUT51), .ZN(new_n814));
  AOI22_X1  g628(.A1(new_n632), .A2(new_n638), .B1(new_n637), .B2(new_n636), .ZN(new_n815));
  OAI22_X1  g629(.A1(new_n815), .A2(new_n614), .B1(new_n646), .B2(new_n647), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n610), .B1(new_n816), .B2(new_n249), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n792), .A2(new_n817), .A3(new_n608), .ZN(new_n818));
  OR3_X1    g632(.A1(new_n810), .A2(new_n811), .A3(new_n818), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n800), .A2(new_n465), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(new_n766), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n819), .A2(new_n773), .A3(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n821), .A2(new_n716), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n736), .A2(new_n413), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(KEYINPUT116), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT50), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n825), .A2(KEYINPUT50), .A3(new_n827), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n721), .A2(new_n263), .A3(new_n464), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n736), .A2(new_n414), .A3(new_n713), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AND4_X1   g649(.A1(new_n679), .A2(new_n835), .A3(new_n672), .A4(new_n670), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n820), .A2(new_n834), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n836), .B1(new_n770), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n832), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n814), .B1(new_n824), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n835), .A2(new_n675), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n841), .A2(G952), .A3(new_n462), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n837), .A2(new_n412), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT48), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n843), .A2(KEYINPUT118), .A3(new_n844), .ZN(new_n845));
  XOR2_X1   g659(.A(KEYINPUT118), .B(KEYINPUT48), .Z(new_n846));
  OAI21_X1  g660(.A(new_n845), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  AOI211_X1 g661(.A(new_n842), .B(new_n847), .C1(new_n756), .C2(new_n822), .ZN(new_n848));
  INV_X1    g662(.A(new_n839), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n849), .A2(KEYINPUT51), .A3(new_n823), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n850), .A2(KEYINPUT117), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n850), .A2(KEYINPUT117), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n840), .B(new_n848), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n771), .A2(new_n704), .A3(new_n729), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n690), .B(new_n701), .C1(new_n260), .C2(new_n262), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n855), .B(KEYINPUT113), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n721), .A2(new_n654), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n857), .B1(new_n762), .B2(new_n760), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT52), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n854), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n859), .B1(new_n854), .B2(new_n858), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n738), .B(new_n739), .C1(new_n675), .C2(new_n682), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n864), .A2(new_n758), .A3(new_n768), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n681), .A2(new_n674), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n657), .A2(new_n658), .A3(new_n664), .A4(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n655), .A2(new_n694), .A3(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT110), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n458), .B1(new_n457), .B2(new_n415), .ZN(new_n871));
  INV_X1    g685(.A(new_n415), .ZN(new_n872));
  AOI211_X1 g686(.A(KEYINPUT20), .B(new_n872), .C1(new_n455), .C2(new_n456), .ZN(new_n873));
  OAI211_X1 g687(.A(new_n473), .B(new_n511), .C1(new_n871), .C2(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n874), .A2(new_n702), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n780), .A2(new_n870), .A3(new_n413), .A4(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n875), .A2(new_n595), .A3(new_n413), .A4(new_n606), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(KEYINPUT110), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n876), .A2(new_n698), .A3(new_n878), .A4(new_n654), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n770), .A2(new_n654), .A3(new_n728), .A4(new_n773), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n879), .A2(new_n785), .A3(new_n880), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n783), .A2(new_n869), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(KEYINPUT111), .B1(new_n866), .B2(new_n882), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n879), .A2(new_n785), .A3(new_n880), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n655), .A2(new_n694), .A3(new_n868), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n884), .A2(new_n885), .A3(new_n779), .A4(new_n782), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT111), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n886), .A2(new_n865), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n863), .B1(new_n883), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(KEYINPUT53), .B1(new_n863), .B2(KEYINPUT112), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n771), .A2(new_n704), .A3(new_n729), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n763), .A2(new_n654), .A3(new_n721), .A4(new_n856), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT52), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n894), .A2(new_n860), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n866), .A2(new_n882), .A3(KEYINPUT111), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n887), .B1(new_n886), .B2(new_n865), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT53), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT112), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n899), .B1(new_n895), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(KEYINPUT54), .B1(new_n891), .B2(new_n902), .ZN(new_n903));
  XNOR2_X1  g717(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n886), .A2(new_n865), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n863), .A2(KEYINPUT53), .A3(new_n905), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n904), .B(new_n906), .C1(new_n898), .C2(KEYINPUT53), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT115), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n889), .A2(new_n899), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n910), .A2(KEYINPUT115), .A3(new_n904), .A4(new_n906), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n903), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  OAI22_X1  g726(.A1(new_n853), .A2(new_n912), .B1(G952), .B2(G953), .ZN(new_n913));
  OR3_X1    g727(.A1(new_n263), .A2(new_n609), .A3(new_n414), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n914), .B(KEYINPUT108), .Z(new_n915));
  NOR2_X1   g729(.A1(new_n716), .A2(new_n798), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n792), .A2(new_n817), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT49), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n917), .A2(new_n918), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n920), .A2(new_n721), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n915), .A2(new_n916), .A3(new_n919), .A4(new_n921), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT109), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n913), .A2(new_n923), .ZN(G75));
  NOR2_X1   g738(.A1(new_n189), .A2(G952), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n898), .A2(KEYINPUT53), .ZN(new_n927));
  INV_X1    g741(.A(new_n906), .ZN(new_n928));
  OAI211_X1 g742(.A(G210), .B(G902), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT56), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n548), .A2(new_n550), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(new_n560), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT55), .Z(new_n934));
  OAI21_X1  g748(.A(new_n926), .B1(new_n931), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n931), .A2(new_n934), .ZN(new_n936));
  OR2_X1    g750(.A1(new_n936), .A2(KEYINPUT119), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(KEYINPUT119), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n935), .B1(new_n937), .B2(new_n938), .ZN(G51));
  NAND2_X1  g753(.A1(new_n910), .A2(new_n906), .ZN(new_n940));
  INV_X1    g754(.A(new_n904), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n907), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n790), .B(KEYINPUT57), .Z(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n816), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n940), .A2(G902), .ZN(new_n947));
  OR2_X1    g761(.A1(new_n947), .A2(new_n789), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n925), .B1(new_n946), .B2(new_n948), .ZN(G54));
  INV_X1    g763(.A(new_n457), .ZN(new_n950));
  NAND2_X1  g764(.A1(KEYINPUT58), .A2(G475), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n950), .B1(new_n947), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n926), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n947), .A2(new_n950), .A3(new_n951), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n953), .A2(new_n954), .ZN(G60));
  NAND2_X1  g769(.A1(G478), .A2(G902), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT59), .Z(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n669), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n925), .B1(new_n943), .B2(new_n959), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n907), .A2(new_n908), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT54), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n889), .A2(new_n890), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n898), .A2(new_n901), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n962), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n961), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n957), .B1(new_n966), .B2(new_n909), .ZN(new_n967));
  OAI211_X1 g781(.A(KEYINPUT120), .B(new_n960), .C1(new_n967), .C2(new_n669), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT120), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n669), .B1(new_n912), .B2(new_n958), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n904), .B1(new_n910), .B2(new_n906), .ZN(new_n971));
  INV_X1    g785(.A(new_n907), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n959), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n926), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n969), .B1(new_n970), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n968), .A2(new_n975), .ZN(G63));
  NAND2_X1  g790(.A1(G217), .A2(G902), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT121), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT60), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n940), .A2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(new_n247), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n940), .A2(new_n689), .A3(new_n979), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n982), .A2(new_n926), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT122), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT61), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n984), .A2(new_n985), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n925), .B1(new_n980), .B2(new_n981), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n990), .A2(new_n986), .A3(new_n987), .A4(new_n983), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n989), .A2(new_n991), .ZN(G66));
  NOR2_X1   g806(.A1(new_n865), .A2(new_n869), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n993), .A2(new_n466), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT123), .Z(new_n995));
  OAI21_X1  g809(.A(G953), .B1(new_n468), .B2(new_n555), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n932), .B1(G898), .B2(new_n189), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n997), .B(new_n998), .ZN(G69));
  NOR2_X1   g813(.A1(new_n393), .A2(new_n394), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n1000), .B(new_n444), .ZN(new_n1001));
  XNOR2_X1  g815(.A(KEYINPUT124), .B(KEYINPUT125), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n1001), .B(new_n1002), .Z(new_n1003));
  INV_X1    g817(.A(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(G227), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n466), .A2(G900), .ZN(new_n1006));
  AND2_X1   g820(.A1(new_n726), .A2(new_n892), .ZN(new_n1007));
  INV_X1    g821(.A(KEYINPUT62), .ZN(new_n1008));
  OR2_X1    g822(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1009), .A2(new_n189), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n412), .A2(new_n773), .A3(new_n867), .ZN(new_n1012));
  OR2_X1    g826(.A1(new_n710), .A2(new_n1012), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n1011), .A2(new_n805), .A3(new_n812), .A4(new_n1013), .ZN(new_n1014));
  OAI221_X1 g828(.A(new_n1004), .B1(new_n1005), .B2(new_n1006), .C1(new_n1010), .C2(new_n1014), .ZN(new_n1015));
  AND4_X1   g829(.A1(new_n412), .A2(new_n795), .A3(new_n708), .A4(new_n763), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n779), .A2(new_n782), .A3(new_n785), .ZN(new_n1017));
  NOR3_X1   g831(.A1(new_n1016), .A2(new_n854), .A3(new_n1017), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1018), .A2(new_n805), .A3(new_n812), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT126), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND4_X1  g835(.A1(new_n1018), .A2(KEYINPUT126), .A3(new_n805), .A4(new_n812), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n466), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n1003), .B1(G227), .B2(new_n1006), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n1015), .B1(new_n1023), .B2(new_n1024), .ZN(G72));
  NAND2_X1  g839(.A1(G472), .A2(G902), .ZN(new_n1026));
  XOR2_X1   g840(.A(new_n1026), .B(KEYINPUT63), .Z(new_n1027));
  NAND2_X1  g841(.A1(new_n1009), .A2(new_n993), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n1027), .B1(new_n1028), .B2(new_n1014), .ZN(new_n1029));
  NOR2_X1   g843(.A1(new_n372), .A2(new_n341), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n1030), .A2(new_n364), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n925), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g846(.A1(new_n1021), .A2(new_n1022), .A3(new_n993), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1033), .A2(new_n1027), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n1034), .A2(new_n364), .A3(new_n1030), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n397), .A2(new_n406), .ZN(new_n1036));
  OAI211_X1 g850(.A(new_n1027), .B(new_n1036), .C1(new_n891), .C2(new_n902), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n1032), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g852(.A(KEYINPUT127), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g854(.A1(new_n1032), .A2(new_n1035), .A3(KEYINPUT127), .A4(new_n1037), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1040), .A2(new_n1041), .ZN(G57));
endmodule


