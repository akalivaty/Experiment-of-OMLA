//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 0 0 1 1 1 1 0 0 1 0 0 0 1 1 1 1 1 1 0 1 1 0 0 0 1 1 1 0 1 1 1 1 0 0 0 1 0 1 0 1 1 0 0 1 0 0 0 1 0 0 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:47 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n567,
    new_n568, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n582, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n616,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT64), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n452), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT66), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  OAI21_X1  g036(.A(new_n460), .B1(new_n461), .B2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n463), .A2(KEYINPUT67), .A3(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n461), .A2(G2104), .ZN(new_n465));
  NAND4_X1  g040(.A1(new_n462), .A2(new_n464), .A3(G137), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G101), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n465), .A2(new_n471), .A3(G125), .ZN(new_n472));
  INV_X1    g047(.A(G113), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n472), .B1(new_n473), .B2(new_n463), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  AND3_X1   g052(.A1(new_n462), .A2(new_n465), .A3(new_n464), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(KEYINPUT68), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n462), .A2(new_n465), .A3(new_n464), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g057(.A(G2105), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n469), .B1(new_n479), .B2(new_n482), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n469), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n484), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  INV_X1    g065(.A(G138), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n462), .A2(new_n464), .A3(new_n492), .A4(new_n465), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  OAI211_X1 g069(.A(G138), .B(new_n469), .C1(new_n494), .C2(KEYINPUT70), .ZN(new_n495));
  AND2_X1   g070(.A1(new_n494), .A2(KEYINPUT70), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AND2_X1   g072(.A1(new_n465), .A2(new_n471), .ZN(new_n498));
  AOI22_X1  g073(.A1(KEYINPUT4), .A2(new_n493), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  AND2_X1   g074(.A1(G126), .A2(G2105), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n462), .A2(new_n464), .A3(new_n465), .A4(new_n500), .ZN(new_n501));
  OAI21_X1  g076(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(G114), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G2105), .ZN(new_n505));
  AOI21_X1  g080(.A(KEYINPUT69), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n469), .A2(G114), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT69), .ZN(new_n508));
  NOR3_X1   g083(.A1(new_n507), .A2(new_n502), .A3(new_n508), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n501), .B1(new_n506), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n499), .A2(new_n510), .ZN(G164));
  NAND2_X1  g086(.A1(G75), .A2(G543), .ZN(new_n512));
  AND2_X1   g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G62), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n512), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G543), .ZN(new_n518));
  OR2_X1    g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n517), .A2(G651), .B1(G50), .B2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G88), .ZN(new_n523));
  NOR2_X1   g098(.A1(KEYINPUT6), .A2(G651), .ZN(new_n524));
  AND2_X1   g099(.A1(KEYINPUT6), .A2(G651), .ZN(new_n525));
  OAI22_X1  g100(.A1(new_n524), .A2(new_n525), .B1(new_n513), .B2(new_n514), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT71), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n519), .A2(new_n520), .ZN(new_n529));
  XNOR2_X1  g104(.A(KEYINPUT5), .B(G543), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n529), .A2(new_n530), .A3(KEYINPUT71), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n522), .B1(new_n523), .B2(new_n532), .ZN(G303));
  INV_X1    g108(.A(G303), .ZN(G166));
  NAND3_X1  g109(.A1(new_n528), .A2(G89), .A3(new_n531), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT72), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT7), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n535), .A2(new_n536), .A3(new_n538), .ZN(new_n539));
  AND2_X1   g114(.A1(G63), .A2(G651), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n521), .A2(G51), .B1(new_n530), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n536), .B1(new_n535), .B2(new_n538), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n542), .A2(new_n543), .ZN(G286));
  INV_X1    g119(.A(G286), .ZN(G168));
  INV_X1    g120(.A(G651), .ZN(new_n546));
  INV_X1    g121(.A(G64), .ZN(new_n547));
  INV_X1    g122(.A(G77), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n515), .A2(new_n547), .B1(new_n548), .B2(new_n518), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT73), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n546), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n551), .B1(new_n550), .B2(new_n549), .ZN(new_n552));
  AND2_X1   g127(.A1(new_n528), .A2(new_n531), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G90), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n521), .A2(G52), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n552), .A2(new_n554), .A3(new_n555), .ZN(G301));
  INV_X1    g131(.A(G301), .ZN(G171));
  NAND2_X1  g132(.A1(new_n553), .A2(G81), .ZN(new_n558));
  NAND2_X1  g133(.A1(G68), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(G56), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n515), .B2(new_n560), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n561), .A2(G651), .B1(G43), .B2(new_n521), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n558), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  NAND4_X1  g140(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND4_X1  g143(.A1(G319), .A2(G483), .A3(G661), .A4(new_n568), .ZN(G188));
  NAND3_X1  g144(.A1(new_n528), .A2(G91), .A3(new_n531), .ZN(new_n570));
  OAI211_X1 g145(.A(G53), .B(G543), .C1(new_n525), .C2(new_n524), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n571), .A2(KEYINPUT74), .A3(KEYINPUT9), .ZN(new_n572));
  NAND2_X1  g147(.A1(KEYINPUT74), .A2(KEYINPUT9), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n521), .A2(G53), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(G78), .A2(G543), .ZN(new_n576));
  INV_X1    g151(.A(G65), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n515), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(G651), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n570), .A2(new_n575), .A3(new_n579), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT75), .ZN(G299));
  INV_X1    g156(.A(G74), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n515), .A2(new_n582), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n583), .A2(G651), .B1(new_n521), .B2(G49), .ZN(new_n584));
  INV_X1    g159(.A(G87), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n532), .B2(new_n585), .ZN(G288));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G61), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n515), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n589), .A2(G651), .B1(G48), .B2(new_n521), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n528), .A2(G86), .A3(new_n531), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(G305));
  NAND2_X1  g167(.A1(new_n521), .A2(G47), .ZN(new_n593));
  INV_X1    g168(.A(G85), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n532), .B2(new_n594), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT76), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n530), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n597), .A2(new_n546), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT77), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n596), .A2(KEYINPUT77), .A3(new_n598), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(G301), .A2(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n521), .A2(G54), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n530), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(new_n546), .ZN(new_n607));
  AND3_X1   g182(.A1(new_n528), .A2(G92), .A3(new_n531), .ZN(new_n608));
  OR2_X1    g183(.A1(new_n608), .A2(KEYINPUT10), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(KEYINPUT10), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n607), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n604), .B1(new_n611), .B2(G868), .ZN(G284));
  OAI21_X1  g187(.A(new_n604), .B1(new_n611), .B2(G868), .ZN(G321));
  INV_X1    g188(.A(G868), .ZN(new_n614));
  NOR2_X1   g189(.A1(G286), .A2(new_n614), .ZN(new_n615));
  XOR2_X1   g190(.A(G299), .B(KEYINPUT78), .Z(new_n616));
  AOI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(new_n614), .ZN(G280));
  XOR2_X1   g192(.A(G280), .B(KEYINPUT79), .Z(G297));
  INV_X1    g193(.A(new_n611), .ZN(new_n619));
  INV_X1    g194(.A(G860), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n619), .B1(G559), .B2(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT80), .ZN(G148));
  NAND2_X1  g197(.A1(new_n563), .A2(new_n614), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n619), .A2(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(new_n614), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g201(.A1(new_n485), .A2(G123), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n469), .A2(G111), .ZN(new_n628));
  OAI21_X1  g203(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n629));
  AND3_X1   g204(.A1(new_n483), .A2(KEYINPUT81), .A3(G135), .ZN(new_n630));
  AOI21_X1  g205(.A(KEYINPUT81), .B1(new_n483), .B2(G135), .ZN(new_n631));
  OAI221_X1 g206(.A(new_n627), .B1(new_n628), .B2(new_n629), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n632), .A2(G2096), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(G2096), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n463), .A2(G2105), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n498), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT12), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT13), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2100), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n633), .A2(new_n634), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT82), .ZN(G156));
  INV_X1    g216(.A(KEYINPUT14), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2427), .B(G2430), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT84), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n647), .B1(new_n644), .B2(new_n645), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n648), .B(new_n649), .Z(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n648), .B(new_n649), .ZN(new_n655));
  INV_X1    g230(.A(new_n653), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2451), .B(G2454), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT85), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n654), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n660), .A2(G14), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n659), .B1(new_n654), .B2(new_n657), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n661), .A2(new_n662), .ZN(G401));
  XNOR2_X1  g238(.A(G2084), .B(G2090), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2072), .B(G2078), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT86), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n666), .B(KEYINPUT17), .Z(new_n669));
  INV_X1    g244(.A(new_n667), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n664), .B(new_n668), .C1(new_n669), .C2(new_n670), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n670), .A2(new_n664), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n666), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT18), .Z(new_n674));
  NOR2_X1   g249(.A1(new_n667), .A2(new_n664), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n669), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n671), .A2(new_n674), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT87), .ZN(new_n678));
  XNOR2_X1  g253(.A(G2096), .B(G2100), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(G227));
  XOR2_X1   g256(.A(G1971), .B(G1976), .Z(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1956), .B(G2474), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1961), .B(G1966), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT20), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n685), .A2(new_n686), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n684), .A2(new_n687), .A3(new_n690), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(new_n684), .B2(new_n690), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(G1991), .B(G1996), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(G1981), .B(G1986), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT89), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n695), .B(new_n699), .ZN(G229));
  NOR2_X1   g275(.A1(G6), .A2(G16), .ZN(new_n701));
  INV_X1    g276(.A(G305), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n701), .B1(new_n702), .B2(G16), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT32), .ZN(new_n704));
  INV_X1    g279(.A(G1981), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  MUX2_X1   g281(.A(G23), .B(G288), .S(G16), .Z(new_n707));
  XOR2_X1   g282(.A(KEYINPUT33), .B(G1976), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(G16), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G22), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G166), .B2(new_n710), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(G1971), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT91), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n709), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  OAI211_X1 g290(.A(new_n706), .B(new_n715), .C1(new_n714), .C2(new_n713), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT34), .Z(new_n717));
  OR2_X1    g292(.A1(G16), .A2(G24), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G290), .B2(new_n710), .ZN(new_n719));
  INV_X1    g294(.A(G1986), .ZN(new_n720));
  AND2_X1   g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(G29), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G25), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n485), .A2(G119), .ZN(new_n724));
  OAI21_X1  g299(.A(KEYINPUT90), .B1(G95), .B2(G2105), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  NOR3_X1   g301(.A1(KEYINPUT90), .A2(G95), .A3(G2105), .ZN(new_n727));
  OAI221_X1 g302(.A(G2104), .B1(G107), .B2(new_n469), .C1(new_n726), .C2(new_n727), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n724), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n483), .A2(G131), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n723), .B1(new_n732), .B2(new_n722), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT35), .B(G1991), .Z(new_n734));
  XOR2_X1   g309(.A(new_n733), .B(new_n734), .Z(new_n735));
  NOR2_X1   g310(.A1(new_n719), .A2(new_n720), .ZN(new_n736));
  NOR3_X1   g311(.A1(new_n721), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n717), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT36), .ZN(new_n739));
  NOR2_X1   g314(.A1(G171), .A2(new_n710), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G5), .B2(new_n710), .ZN(new_n741));
  INV_X1    g316(.A(G1961), .ZN(new_n742));
  INV_X1    g317(.A(G2084), .ZN(new_n743));
  AND2_X1   g318(.A1(KEYINPUT24), .A2(G34), .ZN(new_n744));
  NOR2_X1   g319(.A1(KEYINPUT24), .A2(G34), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n722), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT96), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(new_n476), .B2(new_n722), .ZN(new_n748));
  AOI22_X1  g323(.A1(new_n741), .A2(new_n742), .B1(new_n743), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(G27), .A2(G29), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G164), .B2(G29), .ZN(new_n751));
  INV_X1    g326(.A(G2078), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n749), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n722), .A2(G33), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT25), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n498), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n758), .A2(new_n469), .ZN(new_n759));
  AOI211_X1 g334(.A(new_n757), .B(new_n759), .C1(G139), .C2(new_n483), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n755), .B1(new_n760), .B2(new_n722), .ZN(new_n761));
  XOR2_X1   g336(.A(KEYINPUT95), .B(G2072), .Z(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n722), .A2(G32), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n483), .A2(G141), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n485), .A2(G129), .ZN(new_n766));
  NAND3_X1  g341(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT26), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n767), .A2(new_n768), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n769), .A2(new_n770), .B1(G105), .B2(new_n635), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n765), .A2(new_n766), .A3(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n764), .B1(new_n773), .B2(new_n722), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT27), .B(G1996), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n763), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n564), .A2(G16), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G16), .B2(G19), .ZN(new_n779));
  INV_X1    g354(.A(G1341), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n779), .A2(new_n780), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT31), .B(G11), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT97), .ZN(new_n784));
  INV_X1    g359(.A(G28), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n785), .A2(KEYINPUT30), .ZN(new_n786));
  AOI21_X1  g361(.A(G29), .B1(new_n785), .B2(KEYINPUT30), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n784), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n781), .A2(new_n782), .A3(new_n788), .ZN(new_n789));
  OAI22_X1  g364(.A1(new_n741), .A2(new_n742), .B1(new_n743), .B2(new_n748), .ZN(new_n790));
  NOR4_X1   g365(.A1(new_n754), .A2(new_n777), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n774), .A2(new_n776), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n710), .A2(G21), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G168), .B2(new_n710), .ZN(new_n794));
  INV_X1    g369(.A(G1966), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n791), .A2(new_n792), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n710), .A2(G20), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT23), .ZN(new_n799));
  INV_X1    g374(.A(G299), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(new_n710), .ZN(new_n801));
  INV_X1    g376(.A(G1956), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n710), .A2(G4), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(new_n611), .B2(new_n710), .ZN(new_n805));
  OAI22_X1  g380(.A1(new_n805), .A2(G1348), .B1(new_n632), .B2(new_n722), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(G1348), .B2(new_n805), .ZN(new_n807));
  NOR2_X1   g382(.A1(G29), .A2(G35), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(G162), .B2(G29), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT29), .B(G2090), .Z(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n803), .A2(new_n807), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n722), .A2(G26), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT28), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n483), .A2(G140), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT92), .ZN(new_n816));
  OAI21_X1  g391(.A(KEYINPUT94), .B1(G104), .B2(G2105), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  NOR3_X1   g393(.A1(KEYINPUT94), .A2(G104), .A3(G2105), .ZN(new_n819));
  OAI221_X1 g394(.A(G2104), .B1(G116), .B2(new_n469), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n485), .A2(KEYINPUT93), .A3(G128), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  AOI21_X1  g397(.A(KEYINPUT93), .B1(new_n485), .B2(G128), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n820), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n816), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n814), .B1(new_n825), .B2(new_n722), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(G2067), .ZN(new_n827));
  NOR3_X1   g402(.A1(new_n797), .A2(new_n812), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n739), .A2(new_n828), .ZN(G150));
  INV_X1    g404(.A(G150), .ZN(G311));
  NAND2_X1  g405(.A1(new_n521), .A2(G55), .ZN(new_n831));
  AOI22_X1  g406(.A1(new_n530), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n831), .B1(new_n832), .B2(new_n546), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n833), .B1(new_n553), .B2(G93), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n834), .A2(new_n620), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT37), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n611), .A2(G559), .ZN(new_n837));
  XNOR2_X1  g412(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(G93), .ZN(new_n840));
  OAI221_X1 g415(.A(new_n831), .B1(new_n546), .B2(new_n832), .C1(new_n532), .C2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n563), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n834), .A2(new_n558), .A3(new_n562), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n839), .B(new_n844), .Z(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(KEYINPUT39), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT99), .Z(new_n847));
  OAI21_X1  g422(.A(new_n620), .B1(new_n845), .B2(KEYINPUT39), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n836), .B1(new_n847), .B2(new_n848), .ZN(G145));
  XNOR2_X1  g424(.A(new_n632), .B(new_n476), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n489), .ZN(new_n851));
  INV_X1    g426(.A(G164), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(new_n816), .B2(new_n824), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT92), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n815), .B(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n820), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT93), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n479), .A2(new_n482), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(G2105), .ZN(new_n859));
  INV_X1    g434(.A(G128), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n857), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n856), .B1(new_n861), .B2(new_n821), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n855), .A2(new_n862), .A3(G164), .ZN(new_n863));
  AND3_X1   g438(.A1(new_n853), .A2(new_n772), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n772), .B1(new_n853), .B2(new_n863), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT100), .ZN(new_n866));
  OAI22_X1  g441(.A1(new_n864), .A2(new_n865), .B1(new_n866), .B2(new_n760), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n483), .A2(G142), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n485), .A2(G130), .ZN(new_n869));
  OAI21_X1  g444(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n870));
  INV_X1    g445(.A(G118), .ZN(new_n871));
  AOI22_X1  g446(.A1(new_n870), .A2(KEYINPUT101), .B1(new_n871), .B2(G2105), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n872), .B1(KEYINPUT101), .B2(new_n870), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n868), .A2(new_n869), .A3(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(new_n637), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(new_n731), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NOR3_X1   g452(.A1(new_n816), .A2(new_n824), .A3(new_n852), .ZN(new_n878));
  AOI21_X1  g453(.A(G164), .B1(new_n855), .B2(new_n862), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n773), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n853), .A2(new_n772), .A3(new_n863), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n760), .B(new_n866), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n867), .A2(new_n877), .A3(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT102), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g461(.A1(new_n867), .A2(KEYINPUT102), .A3(new_n877), .A4(new_n883), .ZN(new_n887));
  AND2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n760), .A2(new_n866), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n890), .B1(new_n880), .B2(new_n881), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n876), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(KEYINPUT103), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n877), .B1(new_n867), .B2(new_n883), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT103), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n851), .B1(new_n888), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n886), .A2(new_n887), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n894), .A2(new_n851), .ZN(new_n900));
  AOI21_X1  g475(.A(G37), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g478(.A(G303), .B(G288), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n601), .A2(G305), .A3(new_n602), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(G305), .B1(new_n601), .B2(new_n602), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n905), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(G290), .A2(new_n702), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n910), .A2(new_n904), .A3(new_n906), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(KEYINPUT106), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n912), .A2(KEYINPUT42), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT104), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n916), .B(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n624), .B(new_n844), .ZN(new_n919));
  NOR2_X1   g494(.A1(G299), .A2(new_n611), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(G299), .A2(new_n611), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n921), .A2(new_n922), .A3(KEYINPUT41), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT41), .ZN(new_n924));
  INV_X1    g499(.A(new_n922), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n924), .B1(new_n925), .B2(new_n920), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n919), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n925), .A2(new_n920), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n928), .B1(new_n919), .B2(new_n929), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n915), .A2(new_n918), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n930), .B1(new_n915), .B2(new_n918), .ZN(new_n932));
  OAI21_X1  g507(.A(G868), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n933), .B1(G868), .B2(new_n834), .ZN(G295));
  OAI21_X1  g509(.A(new_n933), .B1(G868), .B2(new_n834), .ZN(G331));
  INV_X1    g510(.A(KEYINPUT107), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n842), .A2(new_n843), .A3(G301), .ZN(new_n937));
  AOI21_X1  g512(.A(G301), .B1(new_n842), .B2(new_n843), .ZN(new_n938));
  OAI21_X1  g513(.A(G286), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n844), .A2(G171), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n842), .A2(new_n843), .A3(G301), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n940), .A2(G168), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n939), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n936), .B1(new_n943), .B2(new_n929), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n923), .A2(new_n926), .A3(new_n942), .A4(new_n939), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n912), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(G37), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n909), .A2(new_n944), .A3(new_n911), .A4(new_n945), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(KEYINPUT43), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT43), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n947), .A2(new_n952), .A3(new_n948), .A4(new_n949), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT108), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT44), .B1(new_n955), .B2(new_n952), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n954), .B(new_n956), .ZN(G397));
  INV_X1    g532(.A(KEYINPUT126), .ZN(new_n958));
  INV_X1    g533(.A(G1384), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n959), .B1(new_n499), .B2(new_n510), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT45), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(KEYINPUT109), .B(G40), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n470), .A2(new_n475), .A3(new_n963), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g540(.A(G290), .B(new_n720), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(G2067), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n825), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(G2067), .B1(new_n816), .B2(new_n824), .ZN(new_n970));
  INV_X1    g545(.A(G1996), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n772), .B(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n969), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n731), .B(new_n734), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n965), .B1(new_n967), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(G8), .ZN(new_n979));
  AND3_X1   g554(.A1(new_n470), .A2(new_n475), .A3(new_n963), .ZN(new_n980));
  OAI211_X1 g555(.A(KEYINPUT45), .B(new_n959), .C1(new_n499), .C2(new_n510), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n962), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n795), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n964), .B1(new_n960), .B2(KEYINPUT50), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT50), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n985), .B(new_n959), .C1(new_n499), .C2(new_n510), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n984), .A2(new_n743), .A3(new_n986), .ZN(new_n987));
  AOI211_X1 g562(.A(new_n979), .B(G286), .C1(new_n983), .C2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G1971), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n982), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G2090), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n984), .A2(new_n991), .A3(new_n986), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(G303), .A2(G8), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT55), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n997));
  OR2_X1    g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n993), .A2(new_n998), .A3(G8), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n988), .A2(new_n999), .A3(KEYINPUT63), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n998), .B1(new_n993), .B2(G8), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n497), .A2(new_n498), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n503), .A2(KEYINPUT69), .A3(new_n505), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n508), .B1(new_n507), .B2(new_n502), .ZN(new_n1006));
  AOI22_X1  g581(.A1(new_n478), .A2(new_n500), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(G1384), .B1(new_n1004), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n980), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G1976), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1009), .B(G8), .C1(new_n1010), .C2(G288), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(KEYINPUT52), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT111), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT49), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n590), .A2(new_n591), .A3(new_n705), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n705), .B1(new_n590), .B2(new_n591), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n1013), .B(new_n1014), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1017), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1019), .A2(new_n1015), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n979), .B1(new_n980), .B2(new_n1008), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1018), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  XOR2_X1   g598(.A(KEYINPUT110), .B(G1976), .Z(new_n1024));
  AOI21_X1  g599(.A(KEYINPUT52), .B1(G288), .B2(new_n1024), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n1022), .B(new_n1025), .C1(new_n1010), .C2(G288), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1012), .A2(new_n1023), .A3(new_n1026), .ZN(new_n1027));
  OAI21_X1  g602(.A(KEYINPUT113), .B1(new_n1001), .B2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n996), .A2(new_n997), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n960), .A2(KEYINPUT50), .ZN(new_n1030));
  AND3_X1   g605(.A1(new_n1030), .A2(new_n980), .A3(new_n986), .ZN(new_n1031));
  AOI22_X1  g606(.A1(new_n1031), .A2(new_n991), .B1(new_n982), .B2(new_n989), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1029), .B1(new_n1032), .B2(new_n979), .ZN(new_n1033));
  AND3_X1   g608(.A1(new_n1012), .A2(new_n1023), .A3(new_n1026), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT113), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1000), .A2(new_n1028), .A3(new_n1036), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1033), .A2(new_n1034), .A3(new_n988), .A4(new_n999), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT63), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g615(.A1(G288), .A2(G1976), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1016), .B1(new_n1023), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1022), .ZN(new_n1043));
  OAI22_X1  g618(.A1(new_n999), .A2(new_n1027), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT112), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT112), .ZN(new_n1046));
  OAI221_X1 g621(.A(new_n1046), .B1(new_n1042), .B2(new_n1043), .C1(new_n999), .C2(new_n1027), .ZN(new_n1047));
  AOI22_X1  g622(.A1(new_n1037), .A2(new_n1040), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n979), .B1(new_n983), .B2(new_n987), .ZN(new_n1049));
  OAI21_X1  g624(.A(G8), .B1(new_n542), .B2(new_n543), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(KEYINPUT118), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT118), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1052), .B(G8), .C1(new_n542), .C2(new_n543), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  NOR4_X1   g629(.A1(new_n1049), .A2(new_n1054), .A3(KEYINPUT119), .A4(KEYINPUT51), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1049), .A2(new_n1054), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT51), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1051), .A2(KEYINPUT119), .A3(new_n1053), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n983), .A2(new_n987), .ZN(new_n1060));
  AOI22_X1  g635(.A1(new_n1058), .A2(new_n1059), .B1(new_n1054), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1055), .B1(new_n1057), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n752), .A2(KEYINPUT53), .ZN(new_n1064));
  OR2_X1    g639(.A1(new_n982), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1066), .B1(new_n982), .B2(G2078), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n980), .B1(new_n1008), .B2(new_n985), .ZN(new_n1068));
  INV_X1    g643(.A(new_n986), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n742), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n1065), .A2(new_n1067), .A3(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1063), .B1(new_n1071), .B2(G301), .ZN(new_n1072));
  INV_X1    g647(.A(G40), .ZN(new_n1073));
  NOR3_X1   g648(.A1(new_n476), .A2(new_n1073), .A3(new_n1064), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1074), .A2(new_n962), .A3(new_n981), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1067), .A2(new_n1070), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(KEYINPUT120), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT120), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1067), .A2(new_n1078), .A3(new_n1070), .A4(new_n1075), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1077), .A2(G171), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1072), .A2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1076), .A2(G171), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n982), .A2(new_n1064), .ZN(new_n1083));
  AOI21_X1  g658(.A(G1961), .B1(new_n984), .B2(new_n986), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(G301), .B1(new_n1085), .B2(new_n1067), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1063), .B1(new_n1082), .B2(new_n1086), .ZN(new_n1087));
  AND3_X1   g662(.A1(new_n1033), .A2(new_n999), .A3(new_n1034), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1062), .A2(new_n1081), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n802), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT114), .ZN(new_n1091));
  OR2_X1    g666(.A1(new_n1091), .A2(KEYINPUT57), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n570), .A2(new_n575), .A3(new_n579), .A4(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1091), .A2(KEYINPUT57), .ZN(new_n1094));
  XOR2_X1   g669(.A(new_n1094), .B(KEYINPUT115), .Z(new_n1095));
  XNOR2_X1  g670(.A(new_n1093), .B(new_n1095), .ZN(new_n1096));
  XNOR2_X1  g671(.A(KEYINPUT56), .B(G2072), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n962), .A2(new_n980), .A3(new_n981), .A4(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1090), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  XOR2_X1   g675(.A(new_n1093), .B(new_n1095), .Z(new_n1101));
  INV_X1    g676(.A(new_n1098), .ZN(new_n1102));
  AOI21_X1  g677(.A(G1956), .B1(new_n984), .B2(new_n986), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1101), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(G1348), .B1(new_n984), .B2(new_n986), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n980), .A2(new_n1008), .A3(new_n968), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n611), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1100), .B1(new_n1104), .B2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1104), .A2(KEYINPUT117), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT117), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1090), .A2(new_n1098), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1111), .B1(new_n1112), .B2(new_n1101), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1099), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT61), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1104), .A2(new_n1099), .A3(KEYINPUT61), .ZN(new_n1117));
  OAI211_X1 g692(.A(KEYINPUT60), .B(new_n1106), .C1(new_n1031), .C2(G1348), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT60), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1119), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1118), .A2(new_n1120), .A3(new_n611), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1117), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT59), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n962), .A2(new_n971), .A3(new_n980), .A4(new_n981), .ZN(new_n1124));
  XNOR2_X1  g699(.A(KEYINPUT116), .B(KEYINPUT58), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n1125), .B(G1341), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1009), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1124), .A2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1123), .B1(new_n1128), .B2(new_n564), .ZN(new_n1129));
  AOI211_X1 g704(.A(KEYINPUT59), .B(new_n563), .C1(new_n1124), .C2(new_n1127), .ZN(new_n1130));
  OAI22_X1  g705(.A1(new_n1129), .A2(new_n1130), .B1(new_n1118), .B2(new_n611), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1122), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1109), .B1(new_n1116), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1048), .B1(new_n1089), .B2(new_n1133), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1086), .A2(new_n1033), .A3(new_n999), .A4(new_n1034), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1060), .A2(G8), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1136), .A2(new_n1058), .A3(new_n1137), .A4(new_n1059), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1059), .A2(new_n1058), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1054), .A2(new_n1060), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1138), .B1(new_n1141), .B2(new_n1056), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT62), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1135), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  OR2_X1    g719(.A1(new_n1144), .A2(KEYINPUT122), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1146), .B1(new_n1144), .B2(KEYINPUT122), .ZN(new_n1147));
  AOI22_X1  g722(.A1(new_n1134), .A2(KEYINPUT121), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT121), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n1048), .B(new_n1149), .C1(new_n1089), .C2(new_n1133), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n978), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n969), .A2(new_n773), .A3(new_n970), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(new_n965), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n965), .A2(new_n971), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1154), .B(KEYINPUT46), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(KEYINPUT47), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT47), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1153), .A2(new_n1158), .A3(new_n1155), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n732), .A2(new_n734), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1160), .B(KEYINPUT123), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n969), .B1(new_n1161), .B2(new_n973), .ZN(new_n1162));
  AOI22_X1  g737(.A1(new_n1157), .A2(new_n1159), .B1(new_n965), .B2(new_n1162), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n601), .A2(new_n720), .A3(new_n602), .A4(new_n965), .ZN(new_n1164));
  AND2_X1   g739(.A1(new_n1164), .A2(KEYINPUT124), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1164), .A2(KEYINPUT124), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT48), .ZN(new_n1167));
  OR3_X1    g742(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n976), .A2(new_n965), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1167), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1163), .A2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1172), .A2(KEYINPUT125), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT125), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1174), .B1(new_n1163), .B2(new_n1171), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n958), .B1(new_n1151), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1134), .A2(KEYINPUT121), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1178), .A2(new_n1150), .A3(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1180), .A2(new_n977), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n1172), .B(KEYINPUT125), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1181), .A2(KEYINPUT126), .A3(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1177), .A2(new_n1183), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g759(.A(G319), .ZN(new_n1186));
  NOR2_X1   g760(.A1(G229), .A2(new_n1186), .ZN(new_n1187));
  OAI211_X1 g761(.A(new_n1187), .B(new_n680), .C1(new_n661), .C2(new_n662), .ZN(new_n1188));
  AOI21_X1  g762(.A(new_n1188), .B1(new_n951), .B2(new_n953), .ZN(new_n1189));
  INV_X1    g763(.A(new_n851), .ZN(new_n1190));
  XNOR2_X1  g764(.A(new_n894), .B(KEYINPUT103), .ZN(new_n1191));
  AOI21_X1  g765(.A(new_n1190), .B1(new_n1191), .B2(new_n899), .ZN(new_n1192));
  NAND2_X1  g766(.A1(new_n899), .A2(new_n900), .ZN(new_n1193));
  NAND2_X1  g767(.A1(new_n1193), .A2(new_n948), .ZN(new_n1194));
  OAI211_X1 g768(.A(new_n1189), .B(KEYINPUT127), .C1(new_n1192), .C2(new_n1194), .ZN(new_n1195));
  INV_X1    g769(.A(new_n1195), .ZN(new_n1196));
  AOI21_X1  g770(.A(KEYINPUT127), .B1(new_n902), .B2(new_n1189), .ZN(new_n1197));
  NOR2_X1   g771(.A1(new_n1196), .A2(new_n1197), .ZN(G308));
  NAND2_X1  g772(.A1(new_n902), .A2(new_n1189), .ZN(G225));
endmodule


