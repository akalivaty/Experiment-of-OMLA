//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 1 0 0 1 1 1 0 1 1 1 1 1 0 1 1 0 0 0 0 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 1 1 0 0 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:14 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n539, new_n540, new_n541, new_n542,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n551, new_n553,
    new_n554, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n605, new_n606, new_n608, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1178;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT65), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT66), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT67), .ZN(new_n455));
  OR2_X1    g030(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT68), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  AOI22_X1  g033(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  AOI22_X1  g035(.A1(new_n460), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT69), .B(G2105), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  AND2_X1   g044(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n470));
  NOR2_X1   g045(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n471));
  OAI211_X1 g046(.A(new_n467), .B(new_n469), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G137), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n466), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n463), .A2(new_n474), .ZN(G160));
  INV_X1    g050(.A(new_n462), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(new_n460), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(G2105), .ZN(new_n479));
  AND2_X1   g054(.A1(new_n460), .A2(new_n479), .ZN(new_n480));
  AOI22_X1  g055(.A1(new_n478), .A2(G124), .B1(new_n480), .B2(G136), .ZN(new_n481));
  OAI221_X1 g056(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n462), .C2(G112), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT70), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  INV_X1    g060(.A(G138), .ZN(new_n486));
  OAI21_X1  g061(.A(KEYINPUT4), .B1(new_n472), .B2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n462), .A2(new_n460), .A3(new_n488), .A4(G138), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  OR2_X1    g065(.A1(G102), .A2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n491), .A2(new_n493), .A3(G2104), .ZN(new_n494));
  AND2_X1   g069(.A1(G126), .A2(G2105), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n467), .A2(new_n469), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT71), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n494), .A2(new_n496), .A3(KEYINPUT71), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n490), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT5), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n508), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT6), .B(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT72), .B(G88), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G50), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n513), .A2(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OR2_X1    g092(.A1(new_n511), .A2(new_n517), .ZN(G303));
  INV_X1    g093(.A(G303), .ZN(G166));
  XNOR2_X1  g094(.A(KEYINPUT74), .B(KEYINPUT7), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT75), .ZN(new_n521));
  NAND4_X1  g096(.A1(new_n521), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT75), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n520), .B(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(new_n513), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G89), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n522), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT76), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n515), .A2(KEYINPUT73), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n515), .A2(KEYINPUT73), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G51), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n508), .A2(G63), .A3(G651), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n530), .A2(new_n535), .A3(new_n536), .ZN(G286));
  INV_X1    g112(.A(G286), .ZN(G168));
  AOI22_X1  g113(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n510), .ZN(new_n540));
  XOR2_X1   g115(.A(new_n540), .B(KEYINPUT77), .Z(new_n541));
  AOI22_X1  g116(.A1(new_n534), .A2(G52), .B1(G90), .B2(new_n527), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  AND3_X1   g119(.A1(new_n531), .A2(G43), .A3(new_n532), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n508), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  INV_X1    g121(.A(G81), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n546), .A2(new_n510), .B1(new_n513), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n551), .A2(new_n554), .ZN(G188));
  INV_X1    g130(.A(new_n515), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G53), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT78), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  OAI21_X1  g134(.A(KEYINPUT79), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n560), .B1(KEYINPUT79), .B2(new_n559), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n508), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n562));
  OAI22_X1  g137(.A1(new_n557), .A2(new_n561), .B1(new_n562), .B2(new_n510), .ZN(new_n563));
  INV_X1    g138(.A(G53), .ZN(new_n564));
  OAI22_X1  g139(.A1(new_n515), .A2(new_n564), .B1(new_n558), .B2(new_n559), .ZN(new_n565));
  INV_X1    g140(.A(G91), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n566), .B2(new_n513), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(G299));
  NAND2_X1  g144(.A1(new_n527), .A2(G87), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n556), .A2(G49), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(G288));
  NAND2_X1  g148(.A1(new_n527), .A2(G86), .ZN(new_n574));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G61), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n507), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(G651), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n556), .A2(G48), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n574), .A2(new_n578), .A3(new_n579), .ZN(G305));
  NAND2_X1  g155(.A1(G72), .A2(G543), .ZN(new_n581));
  INV_X1    g156(.A(G60), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n507), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(G651), .ZN(new_n584));
  INV_X1    g159(.A(G85), .ZN(new_n585));
  INV_X1    g160(.A(G47), .ZN(new_n586));
  OAI221_X1 g161(.A(new_n584), .B1(new_n585), .B2(new_n513), .C1(new_n533), .C2(new_n586), .ZN(G290));
  NAND2_X1  g162(.A1(new_n534), .A2(G54), .ZN(new_n588));
  AND3_X1   g163(.A1(new_n508), .A2(G92), .A3(new_n512), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n589), .B(KEYINPUT10), .ZN(new_n590));
  NAND2_X1  g165(.A1(G79), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G66), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n507), .B2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT80), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n510), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n595), .B1(new_n594), .B2(new_n593), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n588), .A2(new_n590), .A3(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(G868), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(G171), .B2(new_n598), .ZN(G284));
  OAI21_X1  g175(.A(new_n599), .B1(G171), .B2(new_n598), .ZN(G321));
  NAND2_X1  g176(.A1(G299), .A2(new_n598), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(G168), .B2(new_n598), .ZN(G297));
  OAI21_X1  g178(.A(new_n602), .B1(G168), .B2(new_n598), .ZN(G280));
  INV_X1    g179(.A(G860), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n597), .B1(G559), .B2(new_n605), .ZN(new_n606));
  XOR2_X1   g181(.A(new_n606), .B(KEYINPUT81), .Z(G148));
  INV_X1    g182(.A(new_n549), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(new_n598), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n597), .A2(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(new_n598), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g187(.A1(new_n460), .A2(new_n465), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT12), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(KEYINPUT13), .Z(new_n615));
  OR2_X1    g190(.A1(new_n615), .A2(G2100), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n478), .A2(G123), .B1(new_n480), .B2(G135), .ZN(new_n617));
  OAI221_X1 g192(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n462), .C2(G111), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(G2096), .Z(new_n620));
  NAND2_X1  g195(.A1(new_n615), .A2(G2100), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n616), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT82), .Z(G156));
  XNOR2_X1  g198(.A(G2427), .B(G2430), .ZN(new_n624));
  XNOR2_X1  g199(.A(KEYINPUT83), .B(G2438), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT15), .B(G2435), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n626), .A2(new_n627), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n628), .A2(KEYINPUT14), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2443), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2451), .B(G2454), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2446), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n631), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G1341), .B(G1348), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT85), .ZN(new_n639));
  OAI21_X1  g214(.A(G14), .B1(new_n636), .B2(new_n637), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n639), .A2(new_n640), .ZN(G401));
  XOR2_X1   g216(.A(G2084), .B(G2090), .Z(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G2067), .B(G2678), .Z(new_n644));
  NOR2_X1   g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2072), .B(G2078), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT18), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n643), .A2(new_n644), .ZN(new_n649));
  AND3_X1   g224(.A1(new_n649), .A2(KEYINPUT17), .A3(new_n646), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n646), .B1(new_n649), .B2(KEYINPUT17), .ZN(new_n651));
  NOR3_X1   g226(.A1(new_n650), .A2(new_n651), .A3(new_n645), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2096), .B(G2100), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(G227));
  XNOR2_X1  g230(.A(G1971), .B(G1976), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT86), .B(KEYINPUT19), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G1956), .B(G2474), .Z(new_n659));
  XOR2_X1   g234(.A(G1961), .B(G1966), .Z(new_n660));
  AND2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT20), .Z(new_n663));
  NOR2_X1   g238(.A1(new_n659), .A2(new_n660), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n658), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT87), .ZN(new_n666));
  NOR3_X1   g241(.A1(new_n658), .A2(new_n664), .A3(new_n661), .ZN(new_n667));
  NOR3_X1   g242(.A1(new_n663), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G1991), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(G1996), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1981), .B(G1986), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(G1996), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n669), .B(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(new_n671), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n677));
  AND3_X1   g252(.A1(new_n672), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n677), .B1(new_n672), .B2(new_n676), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(G229));
  MUX2_X1   g256(.A(G6), .B(G305), .S(G16), .Z(new_n682));
  XOR2_X1   g257(.A(KEYINPUT32), .B(G1981), .Z(new_n683));
  XOR2_X1   g258(.A(new_n682), .B(new_n683), .Z(new_n684));
  XOR2_X1   g259(.A(KEYINPUT88), .B(G16), .Z(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G22), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(G166), .B2(new_n686), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G1971), .ZN(new_n689));
  NOR2_X1   g264(.A1(G16), .A2(G23), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT89), .Z(new_n691));
  INV_X1    g266(.A(G16), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n691), .B1(G288), .B2(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT33), .B(G1976), .Z(new_n694));
  XOR2_X1   g269(.A(new_n693), .B(new_n694), .Z(new_n695));
  NOR3_X1   g270(.A1(new_n684), .A2(new_n689), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT90), .B(KEYINPUT34), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n696), .A2(new_n697), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n686), .A2(G24), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n584), .B1(new_n585), .B2(new_n513), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(new_n534), .B2(G47), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n700), .B1(new_n702), .B2(new_n686), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(G1986), .Z(new_n704));
  AOI22_X1  g279(.A1(new_n478), .A2(G119), .B1(new_n480), .B2(G131), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n462), .A2(G107), .ZN(new_n706));
  OAI21_X1  g281(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  MUX2_X1   g283(.A(G25), .B(new_n708), .S(G29), .Z(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT35), .B(G1991), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n709), .B(new_n710), .Z(new_n711));
  NAND4_X1  g286(.A1(new_n698), .A2(new_n699), .A3(new_n704), .A4(new_n711), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT36), .Z(new_n713));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G35), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G162), .B2(new_n714), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT29), .B(G2090), .Z(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n686), .A2(G19), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(new_n549), .B2(new_n686), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT91), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(G1341), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n714), .A2(G33), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n724));
  AOI22_X1  g299(.A1(new_n480), .A2(G139), .B1(new_n724), .B2(KEYINPUT25), .ZN(new_n725));
  AOI22_X1  g300(.A1(new_n460), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n726));
  OAI221_X1 g301(.A(new_n725), .B1(KEYINPUT25), .B2(new_n724), .C1(new_n462), .C2(new_n726), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT93), .Z(new_n728));
  OAI21_X1  g303(.A(new_n723), .B1(new_n728), .B2(new_n714), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(G2072), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n718), .A2(new_n722), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n714), .A2(G26), .ZN(new_n732));
  NOR2_X1   g307(.A1(G104), .A2(G2105), .ZN(new_n733));
  OAI21_X1  g308(.A(G2104), .B1(new_n733), .B2(KEYINPUT92), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n462), .A2(G116), .ZN(new_n735));
  AOI211_X1 g310(.A(new_n734), .B(new_n735), .C1(KEYINPUT92), .C2(new_n733), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n480), .A2(G140), .ZN(new_n737));
  INV_X1    g312(.A(G128), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n737), .B1(new_n738), .B2(new_n477), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n732), .B1(new_n741), .B2(new_n714), .ZN(new_n742));
  MUX2_X1   g317(.A(new_n732), .B(new_n742), .S(KEYINPUT28), .Z(new_n743));
  OR2_X1    g318(.A1(new_n743), .A2(G2067), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n686), .A2(G20), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT23), .Z(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(G299), .B2(G16), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(G1956), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n743), .A2(G2067), .ZN(new_n749));
  NOR2_X1   g324(.A1(G5), .A2(G16), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G171), .B2(G16), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(G1961), .ZN(new_n752));
  NAND4_X1  g327(.A1(new_n744), .A2(new_n748), .A3(new_n749), .A4(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n692), .A2(G4), .ZN(new_n754));
  INV_X1    g329(.A(new_n597), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n754), .B1(new_n755), .B2(new_n692), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G1348), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n714), .A2(G27), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G164), .B2(new_n714), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(G2078), .Z(new_n760));
  OR2_X1    g335(.A1(G29), .A2(G32), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n480), .A2(G141), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT95), .Z(new_n763));
  NAND2_X1  g338(.A1(new_n478), .A2(G129), .ZN(new_n764));
  NAND3_X1  g339(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT26), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  AOI22_X1  g343(.A1(new_n767), .A2(new_n768), .B1(G105), .B2(new_n465), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n763), .A2(new_n764), .A3(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n761), .B1(new_n770), .B2(new_n714), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT27), .B(G1996), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT30), .B(G28), .ZN(new_n774));
  OR2_X1    g349(.A1(KEYINPUT31), .A2(G11), .ZN(new_n775));
  NAND2_X1  g350(.A1(KEYINPUT31), .A2(G11), .ZN(new_n776));
  AOI22_X1  g351(.A1(new_n774), .A2(new_n714), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n619), .B2(new_n714), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT24), .ZN(new_n779));
  INV_X1    g354(.A(G34), .ZN(new_n780));
  AOI21_X1  g355(.A(G29), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n779), .B2(new_n780), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G160), .B2(new_n714), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n778), .B1(G2084), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n760), .A2(new_n773), .A3(new_n784), .ZN(new_n785));
  NOR4_X1   g360(.A1(new_n731), .A2(new_n753), .A3(new_n757), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n692), .A2(G21), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G168), .B2(new_n692), .ZN(new_n788));
  INV_X1    g363(.A(G1966), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n729), .A2(G2072), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT94), .Z(new_n792));
  OR2_X1    g367(.A1(new_n783), .A2(G2084), .ZN(new_n793));
  OAI221_X1 g368(.A(new_n793), .B1(new_n771), .B2(new_n772), .C1(new_n751), .C2(G1961), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT96), .Z(new_n795));
  NAND4_X1  g370(.A1(new_n786), .A2(new_n790), .A3(new_n792), .A4(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n713), .A2(new_n796), .ZN(G311));
  INV_X1    g372(.A(G311), .ZN(G150));
  NAND2_X1  g373(.A1(new_n755), .A2(G559), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n800));
  XOR2_X1   g375(.A(new_n799), .B(new_n800), .Z(new_n801));
  NAND2_X1  g376(.A1(new_n527), .A2(G93), .ZN(new_n802));
  AOI22_X1  g377(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n803));
  INV_X1    g378(.A(G55), .ZN(new_n804));
  OAI221_X1 g379(.A(new_n802), .B1(new_n510), .B2(new_n803), .C1(new_n533), .C2(new_n804), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(new_n549), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n801), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n801), .A2(new_n806), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n807), .A2(new_n605), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n805), .A2(G860), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT97), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT37), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n809), .A2(new_n812), .ZN(G145));
  XNOR2_X1  g388(.A(new_n619), .B(G160), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n484), .B(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n480), .A2(G142), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n462), .A2(G118), .ZN(new_n817));
  OAI21_X1  g392(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n816), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n478), .A2(KEYINPUT99), .A3(G130), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT99), .ZN(new_n821));
  INV_X1    g396(.A(G130), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n821), .B1(new_n477), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n819), .B1(new_n820), .B2(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n815), .B(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n708), .B(new_n614), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n497), .B1(new_n487), .B2(new_n489), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT98), .Z(new_n829));
  XNOR2_X1  g404(.A(new_n770), .B(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(new_n741), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(new_n728), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n727), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n827), .A2(new_n835), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n825), .A2(new_n826), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n825), .A2(new_n826), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n837), .A2(new_n833), .A3(new_n834), .A4(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(G37), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n836), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g417(.A(G303), .B(KEYINPUT102), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(G305), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT101), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n702), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n702), .A2(new_n846), .ZN(new_n849));
  OAI21_X1  g424(.A(G288), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n849), .ZN(new_n851));
  INV_X1    g426(.A(G288), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n851), .A2(new_n852), .A3(new_n847), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(KEYINPUT103), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT103), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n850), .A2(new_n853), .A3(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n845), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  NAND4_X1  g433(.A1(new_n844), .A2(new_n856), .A3(new_n853), .A4(new_n850), .ZN(new_n859));
  AND2_X1   g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(KEYINPUT42), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n858), .A2(new_n859), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT42), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n608), .B(new_n805), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT100), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n610), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n755), .A2(G299), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n597), .A2(new_n568), .ZN(new_n870));
  AND3_X1   g445(.A1(new_n869), .A2(KEYINPUT41), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(KEYINPUT41), .B1(new_n869), .B2(new_n870), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n868), .A2(new_n874), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n867), .A2(new_n610), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n869), .A2(new_n870), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n867), .A2(new_n610), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n598), .B1(new_n865), .B2(new_n880), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n861), .A2(new_n875), .A3(new_n864), .A4(new_n879), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT104), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AOI22_X1  g460(.A1(new_n881), .A2(new_n882), .B1(new_n598), .B2(new_n805), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n885), .B1(new_n886), .B2(new_n884), .ZN(G295));
  OAI21_X1  g462(.A(new_n885), .B1(new_n886), .B2(new_n884), .ZN(G331));
  INV_X1    g463(.A(KEYINPUT44), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT43), .ZN(new_n890));
  NAND2_X1  g465(.A1(G286), .A2(new_n866), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NOR2_X1   g467(.A1(G286), .A2(new_n866), .ZN(new_n893));
  OAI21_X1  g468(.A(G301), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(G168), .A2(new_n806), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n895), .A2(new_n891), .A3(G171), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n894), .A2(new_n877), .A3(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n873), .B1(new_n894), .B2(new_n896), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n862), .A2(KEYINPUT105), .ZN(new_n901));
  AOI21_X1  g476(.A(G37), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OAI211_X1 g477(.A(KEYINPUT105), .B(new_n862), .C1(new_n898), .C2(new_n899), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n890), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n862), .B1(new_n898), .B2(new_n899), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n894), .A2(new_n896), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(new_n874), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n907), .A2(new_n860), .A3(new_n897), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n905), .A2(new_n840), .A3(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n909), .A2(KEYINPUT43), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n889), .B1(new_n904), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n901), .A2(new_n907), .A3(new_n897), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n903), .A2(new_n912), .A3(new_n890), .A4(new_n840), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(KEYINPUT106), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n889), .B1(new_n909), .B2(KEYINPUT43), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT106), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n902), .A2(new_n916), .A3(new_n890), .A4(new_n903), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n914), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n911), .A2(new_n918), .ZN(G397));
  INV_X1    g494(.A(KEYINPUT45), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n920), .B1(new_n828), .B2(G1384), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(G40), .ZN(new_n923));
  NOR3_X1   g498(.A1(new_n463), .A2(new_n474), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n770), .B(G1996), .ZN(new_n927));
  INV_X1    g502(.A(G2067), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n740), .B(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n708), .B(new_n710), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n932), .B(KEYINPUT107), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(G290), .B(G1986), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n926), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT53), .ZN(new_n937));
  INV_X1    g512(.A(G1384), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n501), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n939), .A2(KEYINPUT108), .A3(new_n920), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT108), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n494), .A2(new_n496), .A3(KEYINPUT71), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT71), .B1(new_n494), .B2(new_n496), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(G1384), .B1(new_n944), .B2(new_n490), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n941), .B1(new_n945), .B2(KEYINPUT45), .ZN(new_n946));
  INV_X1    g521(.A(new_n474), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n947), .B(G40), .C1(new_n461), .C2(new_n462), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n828), .A2(G1384), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n948), .B1(new_n949), .B2(KEYINPUT45), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n940), .A2(new_n946), .A3(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n937), .B1(new_n951), .B2(G2078), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT124), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI211_X1 g529(.A(KEYINPUT124), .B(new_n937), .C1(new_n951), .C2(G2078), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n487), .A2(new_n489), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n938), .B1(new_n956), .B2(new_n497), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n924), .B1(new_n957), .B2(KEYINPUT50), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT50), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n945), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  OR2_X1    g536(.A1(new_n961), .A2(G1961), .ZN(new_n962));
  NOR3_X1   g537(.A1(new_n937), .A2(new_n923), .A3(G2078), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT125), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n461), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n476), .B1(new_n461), .B2(new_n964), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n947), .B(new_n963), .C1(new_n965), .C2(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n967), .B1(KEYINPUT45), .B2(new_n949), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n968), .A2(KEYINPUT126), .A3(new_n921), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT126), .B1(new_n968), .B2(new_n921), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n954), .A2(new_n955), .A3(new_n962), .A4(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(G301), .B(KEYINPUT54), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n962), .A2(new_n955), .ZN(new_n976));
  AOI211_X1 g551(.A(new_n920), .B(G1384), .C1(new_n944), .C2(new_n490), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n948), .B1(new_n977), .B2(KEYINPUT112), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n921), .A2(KEYINPUT112), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n945), .A2(KEYINPUT45), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  OR3_X1    g557(.A1(new_n982), .A2(new_n937), .A3(G2078), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n976), .A2(new_n954), .A3(new_n983), .A4(new_n973), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n975), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n852), .A2(G1976), .ZN(new_n986));
  INV_X1    g561(.A(G1976), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT52), .B1(G288), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n949), .A2(new_n924), .ZN(new_n989));
  AOI21_X1  g564(.A(KEYINPUT110), .B1(new_n989), .B2(G8), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT110), .ZN(new_n991));
  INV_X1    g566(.A(G8), .ZN(new_n992));
  AOI211_X1 g567(.A(new_n991), .B(new_n992), .C1(new_n949), .C2(new_n924), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n986), .B(new_n988), .C1(new_n990), .C2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT49), .ZN(new_n995));
  INV_X1    g570(.A(G86), .ZN(new_n996));
  INV_X1    g571(.A(G48), .ZN(new_n997));
  OAI22_X1  g572(.A1(new_n513), .A2(new_n996), .B1(new_n515), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n578), .ZN(new_n999));
  OAI21_X1  g574(.A(G1981), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G1981), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n574), .A2(new_n1001), .A3(new_n578), .A4(new_n579), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n995), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1000), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1004), .A2(KEYINPUT49), .ZN(new_n1005));
  OAI22_X1  g580(.A1(new_n1003), .A2(new_n1005), .B1(new_n990), .B2(new_n993), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n989), .A2(G8), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n991), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n989), .A2(KEYINPUT110), .A3(G8), .ZN(new_n1009));
  AOI22_X1  g584(.A1(new_n1008), .A2(new_n1009), .B1(G1976), .B2(new_n852), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n1011));
  OAI211_X1 g586(.A(new_n994), .B(new_n1006), .C1(new_n1010), .C2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G1971), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n951), .A2(new_n1014), .ZN(new_n1015));
  OR3_X1    g590(.A1(new_n958), .A2(G2090), .A3(new_n960), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n992), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT109), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1018), .B(KEYINPUT55), .C1(G166), .C2(new_n992), .ZN(new_n1019));
  XNOR2_X1  g594(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n1020));
  NAND3_X1  g595(.A1(G303), .A2(G8), .A3(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1017), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n499), .A2(new_n500), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n959), .B(new_n938), .C1(new_n956), .C2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(KEYINPUT50), .B1(new_n828), .B2(G1384), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1025), .A2(new_n924), .A3(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1027), .A2(G2090), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1028), .B1(new_n1014), .B2(new_n951), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1023), .B1(new_n1029), .B2(new_n992), .ZN(new_n1030));
  AND3_X1   g605(.A1(new_n1013), .A2(new_n1022), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n985), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G2084), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n961), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT113), .ZN(new_n1035));
  AOI22_X1  g610(.A1(KEYINPUT112), .A2(new_n921), .B1(new_n945), .B2(KEYINPUT45), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n501), .A2(KEYINPUT112), .A3(KEYINPUT45), .A4(new_n938), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(new_n924), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1035), .B(new_n789), .C1(new_n1036), .C2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1034), .A2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1035), .B1(new_n982), .B2(new_n789), .ZN(new_n1041));
  OAI21_X1  g616(.A(G8), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT123), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n789), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT113), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1046), .A2(new_n1034), .A3(new_n1039), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1047), .A2(KEYINPUT123), .A3(G8), .ZN(new_n1048));
  NOR2_X1   g623(.A1(G168), .A2(new_n992), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1049), .A2(KEYINPUT51), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1044), .A2(new_n1048), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT122), .ZN(new_n1052));
  NOR3_X1   g627(.A1(new_n958), .A2(new_n960), .A3(G2084), .ZN(new_n1053));
  AOI21_X1  g628(.A(G1966), .B1(new_n978), .B2(new_n981), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1053), .B1(new_n1054), .B2(new_n1035), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n992), .B1(new_n1055), .B2(new_n1046), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1052), .B(KEYINPUT51), .C1(new_n1056), .C2(new_n1049), .ZN(new_n1057));
  OAI211_X1 g632(.A(KEYINPUT51), .B(G8), .C1(new_n1047), .C2(G286), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT122), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1051), .A2(new_n1057), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1049), .A2(new_n1047), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1032), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  XOR2_X1   g637(.A(KEYINPUT119), .B(G1996), .Z(new_n1063));
  NAND4_X1  g638(.A1(new_n940), .A2(new_n946), .A3(new_n950), .A4(new_n1063), .ZN(new_n1064));
  XOR2_X1   g639(.A(KEYINPUT58), .B(G1341), .Z(new_n1065));
  NAND2_X1  g640(.A1(new_n989), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n608), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT120), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1068), .A2(KEYINPUT59), .ZN(new_n1069));
  AND2_X1   g644(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1068), .A2(KEYINPUT59), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1071), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT117), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT57), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n568), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n1077));
  NOR2_X1   g652(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1077), .B(new_n1079), .C1(new_n563), .C2(new_n567), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1076), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  XOR2_X1   g657(.A(KEYINPUT115), .B(G1956), .Z(new_n1083));
  NAND2_X1  g658(.A1(new_n1027), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT116), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1027), .A2(KEYINPUT116), .A3(new_n1083), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  XNOR2_X1  g663(.A(KEYINPUT56), .B(G2072), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n940), .A2(new_n946), .A3(new_n950), .A4(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1082), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1091));
  AND3_X1   g666(.A1(new_n1027), .A2(KEYINPUT116), .A3(new_n1083), .ZN(new_n1092));
  AOI21_X1  g667(.A(KEYINPUT116), .B1(new_n1027), .B2(new_n1083), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1082), .B(new_n1090), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(KEYINPUT61), .B1(new_n1091), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1090), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(new_n1081), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT61), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1098), .A2(new_n1099), .A3(new_n1094), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1073), .B1(new_n1096), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT60), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n939), .A2(KEYINPUT50), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n948), .B1(new_n949), .B2(new_n959), .ZN(new_n1104));
  AOI21_X1  g679(.A(G1348), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n989), .A2(G2067), .ZN(new_n1106));
  OAI21_X1  g681(.A(KEYINPUT118), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(G1348), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1108), .B1(new_n958), .B2(new_n960), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT118), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1106), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1102), .B1(new_n1107), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1107), .A2(new_n1112), .A3(new_n1102), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT121), .ZN(new_n1116));
  AND3_X1   g691(.A1(new_n1115), .A2(new_n1116), .A3(new_n755), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1116), .B1(new_n1115), .B2(new_n755), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1114), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1115), .A2(new_n755), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(KEYINPUT121), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1115), .A2(new_n1116), .A3(new_n755), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1121), .A2(new_n1113), .A3(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1101), .A2(new_n1119), .A3(new_n1123), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n1107), .A2(new_n1112), .A3(new_n755), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1091), .B1(new_n1125), .B2(new_n1094), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1062), .A2(new_n1127), .ZN(new_n1128));
  AND3_X1   g703(.A1(new_n1006), .A2(new_n987), .A3(new_n852), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n1002), .B(KEYINPUT111), .ZN(new_n1130));
  OAI22_X1  g705(.A1(new_n1129), .A2(new_n1130), .B1(new_n993), .B2(new_n990), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1131), .B1(new_n1022), .B2(new_n1012), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1056), .A2(G168), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1031), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT63), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  OR2_X1    g712(.A1(new_n1017), .A2(KEYINPUT114), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1017), .A2(KEYINPUT114), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1138), .A2(new_n1023), .A3(new_n1139), .ZN(new_n1140));
  AND2_X1   g715(.A1(new_n1013), .A2(new_n1022), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1140), .A2(new_n1134), .A3(new_n1141), .A4(KEYINPUT63), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1132), .B1(new_n1137), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1128), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n976), .A2(new_n954), .A3(new_n983), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1031), .A2(G171), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT62), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1060), .A2(KEYINPUT62), .A3(new_n1061), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1146), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n936), .B1(new_n1144), .B2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n708), .A2(new_n710), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n931), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n741), .A2(new_n928), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n925), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n926), .B1(new_n930), .B2(new_n770), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n926), .A2(KEYINPUT46), .A3(new_n673), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT46), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1159), .B1(new_n925), .B2(G1996), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1157), .A2(new_n1158), .A3(new_n1160), .ZN(new_n1161));
  XOR2_X1   g736(.A(new_n1161), .B(KEYINPUT47), .Z(new_n1162));
  NOR2_X1   g737(.A1(G290), .A2(G1986), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n926), .A2(KEYINPUT48), .A3(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(KEYINPUT48), .B1(new_n926), .B2(new_n1163), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1165), .B1(new_n934), .B2(new_n926), .ZN(new_n1166));
  AOI211_X1 g741(.A(new_n1156), .B(new_n1162), .C1(new_n1164), .C2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1152), .A2(new_n1167), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g743(.A1(new_n904), .A2(new_n910), .ZN(new_n1170));
  INV_X1    g744(.A(G319), .ZN(new_n1171));
  NOR2_X1   g745(.A1(G227), .A2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g746(.A(new_n1172), .B1(new_n639), .B2(new_n640), .ZN(new_n1173));
  INV_X1    g747(.A(KEYINPUT127), .ZN(new_n1174));
  XNOR2_X1  g748(.A(new_n1173), .B(new_n1174), .ZN(new_n1175));
  NAND3_X1  g749(.A1(new_n1175), .A2(new_n680), .A3(new_n841), .ZN(new_n1176));
  NOR2_X1   g750(.A1(new_n1170), .A2(new_n1176), .ZN(G308));
  AND2_X1   g751(.A1(new_n680), .A2(new_n841), .ZN(new_n1178));
  OAI211_X1 g752(.A(new_n1178), .B(new_n1175), .C1(new_n904), .C2(new_n910), .ZN(G225));
endmodule


