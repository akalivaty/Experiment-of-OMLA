//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 0 0 1 1 1 0 0 0 1 0 0 0 1 0 0 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 0 0 0 1 1 0 1 1 1 0 0 1 1 0 0 1 0 1 1 0 0 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:25 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023;
  XNOR2_X1  g000(.A(KEYINPUT67), .B(G953), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G227), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT77), .ZN(new_n189));
  XNOR2_X1  g003(.A(G110), .B(G140), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G143), .ZN(new_n194));
  INV_X1    g008(.A(G128), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(KEYINPUT1), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n197));
  INV_X1    g011(.A(G143), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n197), .B1(new_n198), .B2(G146), .ZN(new_n199));
  NOR3_X1   g013(.A1(new_n193), .A2(KEYINPUT64), .A3(G143), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n194), .B(new_n196), .C1(new_n199), .C2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT81), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n198), .A2(G146), .ZN(new_n203));
  OAI21_X1  g017(.A(KEYINPUT64), .B1(new_n193), .B2(G143), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n197), .A2(new_n198), .A3(G146), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n195), .B1(new_n194), .B2(KEYINPUT1), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n201), .B(new_n202), .C1(new_n206), .C2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n209));
  INV_X1    g023(.A(G107), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n209), .B1(new_n210), .B2(G104), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(G104), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G101), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n210), .A2(KEYINPUT79), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT79), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G107), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n215), .A2(new_n217), .A3(G104), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT78), .B(KEYINPUT3), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n213), .B(new_n214), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT79), .B(G107), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n212), .B1(new_n221), .B2(G104), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G101), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n206), .A2(KEYINPUT81), .A3(new_n196), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n208), .A2(new_n220), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT10), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n223), .A2(new_n220), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT1), .ZN(new_n229));
  OAI21_X1  g043(.A(G128), .B1(new_n203), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n198), .A2(G146), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n194), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n226), .B1(new_n233), .B2(new_n201), .ZN(new_n234));
  AOI22_X1  g048(.A1(new_n225), .A2(new_n226), .B1(new_n228), .B2(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n213), .B1(new_n218), .B2(new_n219), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(KEYINPUT80), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT80), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n213), .B(new_n238), .C1(new_n218), .C2(new_n219), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n237), .A2(G101), .A3(new_n239), .ZN(new_n240));
  AND2_X1   g054(.A1(new_n220), .A2(KEYINPUT4), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n214), .A2(KEYINPUT4), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n237), .A2(new_n239), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(KEYINPUT0), .A2(G128), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  OR2_X1    g060(.A1(KEYINPUT0), .A2(G128), .ZN(new_n247));
  AND2_X1   g061(.A1(new_n247), .A2(new_n245), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n206), .A2(new_n246), .B1(new_n248), .B2(new_n232), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n242), .A2(new_n244), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G134), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(G137), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n252), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(G137), .ZN(new_n258));
  INV_X1    g072(.A(G137), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G134), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n258), .B1(new_n260), .B2(new_n251), .ZN(new_n261));
  INV_X1    g075(.A(G131), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n262), .A2(KEYINPUT66), .ZN(new_n263));
  NOR3_X1   g077(.A1(new_n257), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n263), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n259), .A2(G134), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n266), .B1(new_n252), .B2(new_n256), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n251), .B1(new_n260), .B2(new_n253), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n265), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n264), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n235), .A2(new_n250), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT82), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT82), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n235), .A2(new_n250), .A3(new_n273), .A4(new_n270), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g089(.A(KEYINPUT83), .B(KEYINPUT12), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n227), .A2(new_n201), .A3(new_n233), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n225), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n276), .B1(new_n278), .B2(new_n270), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n270), .B1(new_n225), .B2(new_n277), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n280), .B1(KEYINPUT83), .B2(KEYINPUT12), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n192), .B1(new_n275), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n275), .A2(KEYINPUT84), .A3(new_n192), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n270), .B1(new_n235), .B2(new_n250), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n191), .B1(new_n272), .B2(new_n274), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n289), .A2(KEYINPUT84), .ZN(new_n290));
  OAI211_X1 g104(.A(G469), .B(new_n284), .C1(new_n288), .C2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G469), .ZN(new_n292));
  INV_X1    g106(.A(G902), .ZN(new_n293));
  AOI221_X4 g107(.A(new_n191), .B1(new_n279), .B2(new_n281), .C1(new_n272), .C2(new_n274), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n192), .B1(new_n275), .B2(new_n287), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n292), .B(new_n293), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n292), .A2(new_n293), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n291), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT85), .ZN(new_n300));
  XNOR2_X1  g114(.A(KEYINPUT9), .B(G234), .ZN(new_n301));
  OAI21_X1  g115(.A(G221), .B1(new_n301), .B2(G902), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n299), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n300), .B1(new_n299), .B2(new_n302), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(G214), .B1(G237), .B2(G902), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n233), .A2(new_n201), .ZN(new_n308));
  INV_X1    g122(.A(G125), .ZN(new_n309));
  MUX2_X1   g123(.A(new_n249), .B(new_n308), .S(new_n309), .Z(new_n310));
  INV_X1    g124(.A(G224), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n311), .A2(G953), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n310), .B(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(G110), .B(G122), .ZN(new_n315));
  INV_X1    g129(.A(G119), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G116), .ZN(new_n317));
  INV_X1    g131(.A(G116), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G119), .ZN(new_n319));
  AND2_X1   g133(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n320), .A2(KEYINPUT5), .ZN(new_n321));
  OAI21_X1  g135(.A(G113), .B1(new_n317), .B2(KEYINPUT5), .ZN(new_n322));
  INV_X1    g136(.A(new_n320), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT2), .B(G113), .ZN(new_n324));
  OAI22_X1  g138(.A1(new_n321), .A2(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n325), .A2(new_n227), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  AND2_X1   g141(.A1(new_n240), .A2(new_n241), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n320), .B(new_n324), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n244), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n327), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT86), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n315), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  AND2_X1   g148(.A1(new_n244), .A2(new_n330), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n326), .B1(new_n335), .B2(new_n242), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT86), .ZN(new_n337));
  AND3_X1   g151(.A1(new_n334), .A2(KEYINPUT6), .A3(new_n337), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n327), .B(new_n315), .C1(new_n328), .C2(new_n331), .ZN(new_n339));
  AOI22_X1  g153(.A1(new_n334), .A2(new_n337), .B1(KEYINPUT6), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n314), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(G210), .B1(G237), .B2(G902), .ZN(new_n342));
  OAI21_X1  g156(.A(KEYINPUT7), .B1(new_n311), .B2(G953), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n310), .B(new_n344), .ZN(new_n345));
  XOR2_X1   g159(.A(new_n315), .B(KEYINPUT8), .Z(new_n346));
  NAND2_X1  g160(.A1(new_n325), .A2(new_n227), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n346), .B1(new_n327), .B2(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(G902), .B1(new_n349), .B2(new_n339), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n341), .A2(new_n342), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT89), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n339), .A2(KEYINPUT6), .ZN(new_n354));
  INV_X1    g168(.A(new_n315), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n355), .B1(new_n336), .B2(KEYINPUT86), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n332), .A2(new_n333), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n354), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n334), .A2(KEYINPUT6), .A3(new_n337), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n313), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n350), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(KEYINPUT89), .A3(new_n342), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n353), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n341), .A2(KEYINPUT87), .A3(new_n350), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT87), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n366), .B1(new_n360), .B2(new_n361), .ZN(new_n367));
  XOR2_X1   g181(.A(new_n342), .B(KEYINPUT88), .Z(new_n368));
  NAND3_X1  g182(.A1(new_n365), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n307), .B1(new_n364), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G475), .ZN(new_n371));
  INV_X1    g185(.A(G953), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(KEYINPUT67), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT67), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G953), .ZN(new_n375));
  INV_X1    g189(.A(G237), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n373), .A2(new_n375), .A3(G214), .A4(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n198), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n187), .A2(G143), .A3(G214), .A4(new_n376), .ZN(new_n379));
  NAND2_X1  g193(.A1(KEYINPUT18), .A2(G131), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n380), .B(KEYINPUT90), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n378), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT91), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n378), .A2(new_n379), .A3(KEYINPUT91), .A4(new_n381), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n380), .B1(new_n378), .B2(new_n379), .ZN(new_n387));
  INV_X1    g201(.A(G140), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(G125), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n309), .A2(G140), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n391), .A2(G146), .ZN(new_n392));
  NOR3_X1   g206(.A1(new_n388), .A2(KEYINPUT72), .A3(G125), .ZN(new_n393));
  XNOR2_X1  g207(.A(G125), .B(G140), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n393), .B1(new_n394), .B2(KEYINPUT72), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n392), .B1(new_n395), .B2(G146), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n387), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n386), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n262), .B1(new_n378), .B2(new_n379), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(KEYINPUT17), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n378), .A2(new_n379), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G131), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n378), .A2(new_n379), .A3(new_n262), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n400), .B1(new_n404), .B2(KEYINPUT17), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT73), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n389), .A2(new_n390), .A3(KEYINPUT72), .ZN(new_n407));
  OR3_X1    g221(.A1(new_n388), .A2(KEYINPUT72), .A3(G125), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n407), .A2(new_n408), .A3(KEYINPUT16), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT16), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n389), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n406), .B1(new_n412), .B2(G146), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(G146), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n409), .A2(KEYINPUT73), .A3(new_n193), .A4(new_n411), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n398), .B1(new_n405), .B2(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(G113), .B(G122), .ZN(new_n418));
  XNOR2_X1  g232(.A(KEYINPUT92), .B(G104), .ZN(new_n419));
  XOR2_X1   g233(.A(new_n418), .B(new_n419), .Z(new_n420));
  NAND2_X1  g234(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n420), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n422), .B(new_n398), .C1(new_n405), .C2(new_n416), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n371), .B1(new_n424), .B2(new_n293), .ZN(new_n425));
  NOR2_X1   g239(.A1(G475), .A2(G902), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT93), .ZN(new_n427));
  AOI211_X1 g241(.A(new_n387), .B(new_n396), .C1(new_n384), .C2(new_n385), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT19), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n429), .B1(new_n407), .B2(new_n408), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n394), .A2(KEYINPUT19), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n193), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n378), .A2(new_n379), .A3(new_n262), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n414), .B(new_n432), .C1(new_n433), .C2(new_n399), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n427), .B(new_n420), .C1(new_n428), .C2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n423), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n398), .A2(new_n434), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n427), .B1(new_n438), .B2(new_n420), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n426), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(KEYINPUT20), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n193), .B1(new_n409), .B2(new_n411), .ZN(new_n442));
  INV_X1    g256(.A(new_n431), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n443), .B1(new_n395), .B2(new_n429), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n442), .B1(new_n444), .B2(new_n193), .ZN(new_n445));
  AOI22_X1  g259(.A1(new_n386), .A2(new_n397), .B1(new_n445), .B2(new_n404), .ZN(new_n446));
  OAI21_X1  g260(.A(KEYINPUT93), .B1(new_n446), .B2(new_n422), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n447), .A2(new_n423), .A3(new_n436), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT20), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n448), .A2(new_n449), .A3(new_n426), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n425), .B1(new_n441), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n318), .A2(G122), .ZN(new_n452));
  OAI21_X1  g266(.A(KEYINPUT94), .B1(new_n452), .B2(KEYINPUT14), .ZN(new_n453));
  INV_X1    g267(.A(G122), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(G116), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n452), .A2(KEYINPUT14), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n453), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NOR3_X1   g271(.A1(new_n452), .A2(KEYINPUT94), .A3(KEYINPUT14), .ZN(new_n458));
  OAI21_X1  g272(.A(G107), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n198), .A2(G128), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n195), .A2(G143), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(G134), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n460), .A2(new_n461), .A3(new_n255), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n455), .A2(new_n452), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  AOI22_X1  g280(.A1(new_n463), .A2(new_n464), .B1(new_n466), .B2(new_n221), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n459), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT13), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n460), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(new_n461), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n460), .A2(new_n469), .ZN(new_n472));
  OAI21_X1  g286(.A(G134), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n466), .A2(new_n221), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n221), .A2(new_n455), .A3(new_n452), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n473), .B(new_n464), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(G217), .ZN(new_n477));
  NOR3_X1   g291(.A1(new_n301), .A2(new_n477), .A3(G953), .ZN(new_n478));
  AND3_X1   g292(.A1(new_n468), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n478), .B1(new_n468), .B2(new_n476), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n293), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT95), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(G478), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n484), .A2(KEYINPUT15), .ZN(new_n485));
  OAI211_X1 g299(.A(KEYINPUT95), .B(new_n293), .C1(new_n479), .C2(new_n480), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n483), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  OR2_X1    g301(.A1(new_n481), .A2(new_n485), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(G952), .ZN(new_n490));
  AOI211_X1 g304(.A(G953), .B(new_n490), .C1(G234), .C2(G237), .ZN(new_n491));
  AOI211_X1 g305(.A(new_n293), .B(new_n187), .C1(G234), .C2(G237), .ZN(new_n492));
  XNOR2_X1  g306(.A(KEYINPUT21), .B(G898), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n451), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  XOR2_X1   g311(.A(G119), .B(G128), .Z(new_n498));
  XNOR2_X1  g312(.A(KEYINPUT24), .B(G110), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT23), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n501), .B1(new_n316), .B2(G128), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n195), .A2(KEYINPUT23), .A3(G119), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n502), .B(new_n503), .C1(G119), .C2(new_n195), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n500), .B1(new_n504), .B2(G110), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n505), .B(KEYINPUT75), .ZN(new_n506));
  OR3_X1    g320(.A1(new_n506), .A2(new_n392), .A3(new_n442), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT74), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n498), .A2(new_n499), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n509), .B1(G110), .B2(new_n504), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n416), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n508), .B1(new_n416), .B2(new_n510), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n507), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n187), .A2(G221), .A3(G234), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT22), .B(G137), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n514), .B(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n507), .B(new_n516), .C1(new_n511), .C2(new_n512), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n518), .A2(new_n293), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(KEYINPUT25), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT25), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n518), .A2(new_n522), .A3(new_n293), .A4(new_n519), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n477), .B1(G234), .B2(new_n293), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n521), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n524), .A2(G902), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n518), .A2(new_n519), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(KEYINPUT76), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT76), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n518), .A2(new_n529), .A3(new_n519), .A4(new_n526), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n525), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n194), .B(new_n246), .C1(new_n199), .C2(new_n200), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n232), .A2(new_n245), .A3(new_n247), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n267), .A2(new_n265), .A3(new_n268), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n263), .B1(new_n257), .B2(new_n261), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n262), .B1(new_n257), .B2(new_n261), .ZN(new_n538));
  NOR3_X1   g352(.A1(new_n256), .A2(new_n266), .A3(new_n262), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  AOI22_X1  g354(.A1(new_n538), .A2(new_n540), .B1(new_n201), .B2(new_n233), .ZN(new_n541));
  NOR3_X1   g355(.A1(new_n537), .A2(new_n541), .A3(KEYINPUT30), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT30), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n249), .B1(new_n264), .B2(new_n269), .ZN(new_n544));
  AOI21_X1  g358(.A(G131), .B1(new_n267), .B2(new_n268), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n308), .B1(new_n545), .B2(new_n539), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n543), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n330), .B1(new_n542), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT69), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n187), .A2(G210), .A3(new_n376), .ZN(new_n550));
  XOR2_X1   g364(.A(KEYINPUT68), .B(KEYINPUT27), .Z(new_n551));
  XNOR2_X1  g365(.A(new_n550), .B(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(KEYINPUT26), .B(G101), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n552), .B(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n544), .A2(new_n546), .A3(new_n329), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n548), .A2(new_n549), .A3(new_n554), .A4(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT31), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n555), .ZN(new_n559));
  OAI21_X1  g373(.A(KEYINPUT30), .B1(new_n537), .B2(new_n541), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n544), .A2(new_n546), .A3(new_n543), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n559), .B1(new_n562), .B2(new_n330), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n563), .A2(new_n549), .A3(KEYINPUT31), .A4(new_n554), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n558), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n329), .B1(new_n544), .B2(new_n546), .ZN(new_n566));
  OAI21_X1  g380(.A(KEYINPUT28), .B1(new_n559), .B2(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(KEYINPUT70), .B1(new_n559), .B2(KEYINPUT28), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT70), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT28), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n555), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n567), .A2(new_n568), .A3(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n554), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n565), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(G472), .A2(G902), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n575), .A2(KEYINPUT32), .A3(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT32), .ZN(new_n578));
  AOI22_X1  g392(.A1(new_n558), .A2(new_n564), .B1(new_n573), .B2(new_n572), .ZN(new_n579));
  INV_X1    g393(.A(new_n576), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT71), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n577), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n575), .A2(KEYINPUT71), .A3(KEYINPUT32), .A4(new_n576), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n548), .A2(new_n555), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n573), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n567), .A2(new_n568), .A3(new_n554), .A4(new_n571), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT29), .ZN(new_n589));
  AND3_X1   g403(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n293), .B1(new_n588), .B2(new_n589), .ZN(new_n591));
  OAI21_X1  g405(.A(G472), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n531), .B1(new_n585), .B2(new_n592), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n305), .A2(new_n370), .A3(new_n497), .A4(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(G101), .ZN(G3));
  INV_X1    g409(.A(new_n342), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n596), .B1(new_n360), .B2(new_n361), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n351), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n306), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n441), .A2(new_n450), .ZN(new_n600));
  INV_X1    g414(.A(new_n425), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT33), .ZN(new_n603));
  INV_X1    g417(.A(new_n480), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT96), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n606), .B1(new_n479), .B2(new_n480), .ZN(new_n607));
  INV_X1    g421(.A(new_n479), .ZN(new_n608));
  OAI211_X1 g422(.A(new_n608), .B(new_n604), .C1(new_n605), .C2(new_n603), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n484), .A2(G902), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n483), .A2(new_n486), .ZN(new_n612));
  AOI22_X1  g426(.A1(new_n610), .A2(new_n611), .B1(new_n612), .B2(new_n484), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n602), .A2(new_n614), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n599), .A2(new_n494), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(G902), .B1(new_n565), .B2(new_n574), .ZN(new_n617));
  INV_X1    g431(.A(G472), .ZN(new_n618));
  OAI22_X1  g432(.A1(new_n617), .A2(new_n618), .B1(new_n580), .B2(new_n579), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n531), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n305), .A2(new_n616), .A3(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT34), .B(G104), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G6));
  INV_X1    g437(.A(KEYINPUT97), .ZN(new_n624));
  INV_X1    g438(.A(new_n450), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n449), .B1(new_n448), .B2(new_n426), .ZN(new_n626));
  OAI211_X1 g440(.A(new_n601), .B(new_n489), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n624), .B1(new_n627), .B2(new_n494), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n307), .B1(new_n351), .B2(new_n597), .ZN(new_n629));
  INV_X1    g443(.A(new_n494), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n451), .A2(KEYINPUT97), .A3(new_n630), .A4(new_n489), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n628), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT98), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n628), .A2(new_n629), .A3(KEYINPUT98), .A4(new_n631), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n636), .A2(new_n305), .A3(new_n620), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT35), .B(G107), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G9));
  NOR2_X1   g453(.A1(new_n517), .A2(KEYINPUT36), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n513), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n526), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n525), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n497), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n644), .A2(new_n619), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n305), .A2(new_n370), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT37), .B(G110), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(KEYINPUT99), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n646), .B(new_n648), .ZN(G12));
  OR2_X1    g463(.A1(new_n289), .A2(KEYINPUT84), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n286), .B1(new_n289), .B2(KEYINPUT84), .ZN(new_n651));
  AOI211_X1 g465(.A(new_n292), .B(new_n283), .C1(new_n650), .C2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n296), .A2(new_n298), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n302), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(KEYINPUT85), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n299), .A2(new_n300), .A3(new_n302), .ZN(new_n656));
  INV_X1    g470(.A(G900), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n491), .B1(new_n492), .B2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n627), .A2(new_n658), .ZN(new_n659));
  AND3_X1   g473(.A1(new_n629), .A2(new_n659), .A3(new_n643), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n585), .A2(new_n592), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n655), .A2(new_n656), .A3(new_n660), .A4(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G128), .ZN(G30));
  OAI21_X1  g477(.A(new_n573), .B1(new_n559), .B2(new_n566), .ZN(new_n664));
  OR2_X1    g478(.A1(new_n664), .A2(KEYINPUT100), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n563), .A2(new_n554), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n664), .A2(KEYINPUT100), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  AOI21_X1  g482(.A(G902), .B1(new_n668), .B2(KEYINPUT101), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n669), .B1(KEYINPUT101), .B2(new_n668), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(G472), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n585), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(KEYINPUT102), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n451), .B1(new_n488), .B2(new_n487), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n306), .ZN(new_n676));
  AOI21_X1  g490(.A(KEYINPUT89), .B1(new_n362), .B2(new_n342), .ZN(new_n677));
  NOR4_X1   g491(.A1(new_n360), .A2(new_n361), .A3(new_n352), .A4(new_n596), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n369), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(KEYINPUT38), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT38), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n364), .A2(new_n681), .A3(new_n369), .ZN(new_n682));
  AOI211_X1 g496(.A(new_n643), .B(new_n676), .C1(new_n680), .C2(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(new_n658), .B(KEYINPUT39), .Z(new_n684));
  NAND2_X1  g498(.A1(new_n305), .A2(new_n684), .ZN(new_n685));
  OAI211_X1 g499(.A(new_n674), .B(new_n683), .C1(KEYINPUT40), .C2(new_n685), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n685), .A2(KEYINPUT40), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(new_n198), .ZN(G45));
  NOR3_X1   g503(.A1(new_n451), .A2(new_n613), .A3(new_n658), .ZN(new_n690));
  AND3_X1   g504(.A1(new_n629), .A2(new_n690), .A3(new_n643), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n655), .A2(new_n656), .A3(new_n661), .A4(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G146), .ZN(G48));
  INV_X1    g507(.A(new_n592), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n694), .B1(new_n583), .B2(new_n584), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n275), .A2(new_n287), .ZN(new_n696));
  AOI22_X1  g510(.A1(new_n696), .A2(new_n191), .B1(new_n289), .B2(new_n282), .ZN(new_n697));
  OAI211_X1 g511(.A(KEYINPUT103), .B(G469), .C1(new_n697), .C2(G902), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n696), .A2(new_n191), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n289), .A2(new_n282), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(KEYINPUT103), .A2(G469), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n701), .A2(new_n293), .A3(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n698), .A2(new_n703), .A3(new_n302), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n695), .A2(new_n531), .A3(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT104), .ZN(new_n706));
  AND3_X1   g520(.A1(new_n705), .A2(new_n706), .A3(new_n616), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n706), .B1(new_n705), .B2(new_n616), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XOR2_X1   g523(.A(KEYINPUT41), .B(G113), .Z(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G15));
  NAND2_X1  g525(.A1(new_n636), .A2(new_n705), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G116), .ZN(G18));
  NOR2_X1   g527(.A1(new_n695), .A2(new_n644), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n704), .A2(new_n599), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G119), .ZN(G21));
  NOR2_X1   g531(.A1(new_n704), .A2(new_n494), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n629), .A2(new_n675), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n528), .A2(new_n530), .ZN(new_n720));
  INV_X1    g534(.A(new_n524), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n721), .B1(new_n520), .B2(KEYINPUT25), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n720), .B1(new_n523), .B2(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n554), .B1(new_n572), .B2(KEYINPUT105), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n724), .B1(KEYINPUT105), .B2(new_n572), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n580), .B1(new_n725), .B2(new_n565), .ZN(new_n726));
  OAI21_X1  g540(.A(KEYINPUT106), .B1(new_n617), .B2(new_n618), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT106), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n728), .B(G472), .C1(new_n579), .C2(G902), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n726), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n718), .A2(new_n719), .A3(new_n723), .A4(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G122), .ZN(G24));
  NAND2_X1  g546(.A1(new_n727), .A2(new_n729), .ZN(new_n733));
  INV_X1    g547(.A(new_n726), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n733), .A2(new_n643), .A3(new_n690), .A4(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n629), .A2(new_n302), .A3(new_n698), .A4(new_n703), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(new_n309), .ZN(G27));
  OAI211_X1 g552(.A(new_n369), .B(new_n306), .C1(new_n677), .C2(new_n678), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n299), .A2(new_n302), .ZN(new_n741));
  INV_X1    g555(.A(new_n690), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n742), .A2(KEYINPUT42), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n593), .A2(new_n740), .A3(new_n741), .A4(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT42), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n577), .A2(new_n581), .A3(new_n592), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n723), .A2(new_n690), .A3(new_n746), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n739), .A2(new_n747), .A3(new_n654), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n744), .B1(new_n745), .B2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(new_n262), .ZN(G33));
  NOR2_X1   g564(.A1(new_n739), .A2(new_n654), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n751), .A2(new_n593), .A3(new_n659), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G134), .ZN(G36));
  OAI21_X1  g567(.A(new_n284), .B1(new_n288), .B2(new_n290), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT45), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n292), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n283), .B1(new_n650), .B2(new_n651), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(KEYINPUT45), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n297), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n296), .B1(new_n759), .B2(KEYINPUT46), .ZN(new_n760));
  OAI21_X1  g574(.A(G469), .B1(new_n757), .B2(KEYINPUT45), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n754), .A2(new_n755), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT46), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n763), .A2(new_n764), .A3(new_n297), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n302), .B1(new_n760), .B2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(KEYINPUT107), .B(KEYINPUT108), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n767), .A2(new_n684), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n768), .B1(new_n767), .B2(new_n684), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n451), .A2(new_n614), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(KEYINPUT43), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT43), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n451), .A2(new_n614), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(KEYINPUT109), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n777), .A2(new_n619), .A3(new_n643), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT110), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT44), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n778), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n740), .B1(new_n778), .B2(new_n780), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n779), .B1(new_n778), .B2(new_n780), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n781), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n771), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G137), .ZN(G39));
  INV_X1    g600(.A(KEYINPUT47), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n766), .A2(new_n787), .ZN(new_n788));
  OAI211_X1 g602(.A(KEYINPUT47), .B(new_n302), .C1(new_n760), .C2(new_n765), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NOR4_X1   g604(.A1(new_n661), .A2(new_n739), .A3(new_n742), .A4(new_n723), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G140), .ZN(G42));
  INV_X1    g607(.A(new_n491), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n776), .A2(new_n794), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n730), .A2(new_n723), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AOI211_X1 g611(.A(new_n490), .B(G953), .C1(new_n797), .C2(new_n715), .ZN(new_n798));
  NOR4_X1   g612(.A1(new_n739), .A2(new_n704), .A3(new_n794), .A4(new_n531), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n673), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n798), .B1(new_n800), .B2(new_n615), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n739), .A2(new_n704), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT114), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n802), .A2(new_n803), .A3(new_n795), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n803), .B1(new_n802), .B2(new_n795), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n723), .B(new_n746), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n806), .A2(KEYINPUT48), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(KEYINPUT48), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n801), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT115), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n698), .A2(new_n703), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n788), .B(new_n789), .C1(new_n302), .C2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n795), .A2(new_n796), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n813), .A2(new_n739), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n680), .A2(new_n682), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n704), .A2(new_n306), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n797), .A2(new_n816), .A3(KEYINPUT50), .A4(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT50), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n680), .A2(new_n682), .A3(new_n817), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n819), .B1(new_n813), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n730), .A2(new_n643), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n823), .B1(new_n804), .B2(new_n805), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n673), .A2(new_n451), .A3(new_n613), .A4(new_n799), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n822), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n815), .A2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT51), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n810), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AOI211_X1 g643(.A(KEYINPUT115), .B(KEYINPUT51), .C1(new_n815), .C2(new_n826), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n809), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n822), .A2(new_n824), .A3(new_n825), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n832), .B1(new_n812), .B2(new_n814), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n833), .A2(KEYINPUT116), .A3(KEYINPUT51), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n815), .A2(new_n826), .A3(KEYINPUT51), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT116), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(KEYINPUT117), .B1(new_n831), .B2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n840));
  OR2_X1    g654(.A1(new_n735), .A2(new_n736), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n643), .A2(new_n658), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n741), .A2(new_n672), .A3(new_n719), .A4(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n662), .A2(new_n692), .A3(new_n841), .A4(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT52), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n629), .A2(new_n659), .A3(new_n643), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n695), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n737), .B1(new_n305), .B2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n849), .A2(KEYINPUT52), .A3(new_n692), .A4(new_n843), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n846), .A2(new_n850), .A3(KEYINPUT112), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT112), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n844), .A2(new_n852), .A3(new_n845), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n655), .A2(new_n370), .A3(new_n656), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n661), .A2(new_n497), .A3(new_n723), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n716), .B(new_n731), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n705), .A2(new_n706), .A3(new_n616), .ZN(new_n858));
  INV_X1    g672(.A(new_n708), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n494), .B1(new_n615), .B2(new_n627), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n861), .A2(new_n679), .A3(new_n306), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n305), .A2(new_n620), .A3(new_n862), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n646), .A2(new_n863), .A3(new_n712), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n489), .A2(new_n658), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n865), .B(new_n601), .C1(new_n625), .C2(new_n626), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT111), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT111), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n451), .A2(new_n868), .A3(new_n865), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n867), .A2(new_n643), .A3(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n695), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n871), .A2(new_n655), .A3(new_n656), .A4(new_n740), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n751), .A2(new_n690), .A3(new_n823), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n872), .A2(new_n752), .A3(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n874), .A2(new_n749), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n860), .A2(new_n864), .A3(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n840), .B1(new_n854), .B2(new_n876), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n872), .A2(new_n752), .A3(new_n873), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n751), .A2(new_n593), .A3(new_n743), .ZN(new_n879));
  INV_X1    g693(.A(new_n747), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n745), .B1(new_n751), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n878), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n629), .A2(new_n675), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n884), .A2(new_n704), .A3(new_n494), .ZN(new_n885));
  AOI22_X1  g699(.A1(new_n885), .A2(new_n796), .B1(new_n714), .B2(new_n715), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n594), .B(new_n886), .C1(new_n707), .C2(new_n708), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n646), .A2(new_n863), .A3(new_n712), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n883), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n846), .A2(new_n850), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n889), .A2(KEYINPUT53), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n877), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(KEYINPUT54), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n889), .A2(KEYINPUT53), .A3(new_n853), .A4(new_n851), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n846), .A2(new_n850), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n840), .B1(new_n876), .B2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT113), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT54), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n894), .A2(new_n896), .A3(new_n897), .A4(new_n898), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n893), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g714(.A(KEYINPUT115), .B1(new_n833), .B2(KEYINPUT51), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n827), .A2(new_n810), .A3(new_n828), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n834), .A2(new_n837), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT117), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n903), .A2(new_n904), .A3(new_n905), .A4(new_n809), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n894), .A2(new_n898), .A3(new_n896), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(KEYINPUT113), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n839), .A2(new_n900), .A3(new_n906), .A4(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n490), .A2(new_n372), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n811), .A2(KEYINPUT49), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n811), .A2(KEYINPUT49), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n451), .A2(new_n614), .A3(new_n306), .A4(new_n302), .ZN(new_n914));
  NOR4_X1   g728(.A1(new_n912), .A2(new_n913), .A3(new_n531), .A4(new_n914), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n673), .A2(new_n915), .A3(new_n816), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n911), .A2(new_n916), .ZN(G75));
  NOR3_X1   g731(.A1(new_n338), .A2(new_n340), .A3(new_n314), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n918), .A2(new_n360), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT55), .ZN(new_n920));
  AOI21_X1  g734(.A(KEYINPUT53), .B1(new_n889), .B2(new_n890), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n860), .A2(KEYINPUT53), .A3(new_n875), .A4(new_n864), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n854), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n924), .A2(new_n293), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(G210), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT56), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n920), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n187), .A2(G952), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n920), .A2(new_n927), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n930), .B1(new_n925), .B2(new_n368), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n928), .A2(new_n929), .A3(new_n931), .ZN(G51));
  OAI21_X1  g746(.A(KEYINPUT54), .B1(new_n921), .B2(new_n923), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n933), .A2(KEYINPUT118), .A3(new_n907), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT118), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n935), .B(KEYINPUT54), .C1(new_n921), .C2(new_n923), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n297), .B(KEYINPUT57), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n934), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n701), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n925), .A2(new_n763), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n929), .B1(new_n939), .B2(new_n940), .ZN(G54));
  NAND3_X1  g755(.A1(new_n925), .A2(KEYINPUT58), .A3(G475), .ZN(new_n942));
  INV_X1    g756(.A(new_n448), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n942), .A2(new_n943), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n944), .A2(new_n945), .A3(new_n929), .ZN(G60));
  INV_X1    g760(.A(new_n610), .ZN(new_n947));
  XNOR2_X1  g761(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n484), .A2(new_n293), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n948), .B(new_n949), .Z(new_n950));
  NOR2_X1   g764(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n934), .A2(new_n936), .A3(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT120), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n934), .A2(KEYINPUT120), .A3(new_n936), .A4(new_n951), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n908), .A2(new_n893), .A3(new_n899), .ZN(new_n957));
  INV_X1    g771(.A(new_n950), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n929), .B1(new_n959), .B2(new_n947), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n956), .A2(new_n960), .ZN(G63));
  NAND2_X1  g775(.A1(G217), .A2(G902), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(KEYINPUT60), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n924), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n641), .ZN(new_n965));
  INV_X1    g779(.A(new_n929), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n518), .A2(new_n519), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n967), .B1(new_n924), .B2(new_n963), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n965), .A2(new_n966), .A3(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT61), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(G66));
  NAND2_X1  g785(.A1(new_n860), .A2(new_n864), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT121), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n187), .ZN(new_n974));
  OAI21_X1  g788(.A(G953), .B1(new_n493), .B2(new_n311), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT122), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  OAI211_X1 g791(.A(new_n358), .B(new_n359), .C1(G898), .C2(new_n187), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n977), .B(new_n978), .ZN(G69));
  NAND2_X1  g793(.A1(new_n785), .A2(new_n792), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT62), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n849), .A2(new_n692), .ZN(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  OAI211_X1 g797(.A(new_n981), .B(new_n983), .C1(new_n686), .C2(new_n687), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n615), .A2(new_n627), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n593), .A2(new_n740), .A3(new_n985), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n685), .A2(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  AND2_X1   g802(.A1(new_n984), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(KEYINPUT62), .B1(new_n688), .B2(new_n982), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n187), .B1(new_n980), .B2(new_n991), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n562), .B(new_n444), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n993), .B(KEYINPUT123), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT125), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n187), .B1(G227), .B2(G900), .ZN(new_n996));
  AOI22_X1  g810(.A1(new_n992), .A2(new_n994), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OR2_X1    g811(.A1(new_n996), .A2(new_n995), .ZN(new_n998));
  INV_X1    g812(.A(new_n187), .ZN(new_n999));
  AOI22_X1  g813(.A1(new_n771), .A2(new_n784), .B1(new_n790), .B2(new_n791), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n983), .A2(new_n882), .A3(new_n752), .ZN(new_n1001));
  AND3_X1   g815(.A1(new_n719), .A2(new_n723), .A3(new_n746), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1001), .B1(new_n771), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n999), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n999), .A2(new_n657), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1005), .B(KEYINPUT124), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n993), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  AND3_X1   g821(.A1(new_n997), .A2(new_n998), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n998), .B1(new_n997), .B2(new_n1007), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n1008), .A2(new_n1009), .ZN(G72));
  NAND2_X1  g824(.A1(G472), .A2(G902), .ZN(new_n1011));
  XOR2_X1   g825(.A(new_n1011), .B(KEYINPUT63), .Z(new_n1012));
  XOR2_X1   g826(.A(new_n1012), .B(KEYINPUT126), .Z(new_n1013));
  NAND3_X1  g827(.A1(new_n1000), .A2(new_n990), .A3(new_n989), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1013), .B1(new_n1014), .B2(new_n973), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n1015), .A2(new_n554), .A3(new_n586), .ZN(new_n1016));
  INV_X1    g830(.A(new_n1012), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1017), .B1(new_n587), .B2(new_n666), .ZN(new_n1018));
  XNOR2_X1  g832(.A(new_n1018), .B(KEYINPUT127), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n929), .B1(new_n892), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1013), .B1(new_n1021), .B2(new_n973), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n1022), .A2(new_n573), .A3(new_n563), .ZN(new_n1023));
  AND3_X1   g837(.A1(new_n1016), .A2(new_n1020), .A3(new_n1023), .ZN(G57));
endmodule


