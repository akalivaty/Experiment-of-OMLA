//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 0 1 0 0 1 0 1 1 0 0 1 0 1 0 1 0 0 1 0 1 1 0 0 0 0 1 1 0 0 0 1 0 0 1 1 0 1 0 1 0 0 1 1 0 1 0 0 1 1 1 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:44 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n649, new_n650, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n665, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958;
  INV_X1    g000(.A(G104), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT3), .B1(new_n187), .B2(G107), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT3), .ZN(new_n189));
  INV_X1    g003(.A(G107), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G104), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n187), .A2(G107), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n188), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G101), .ZN(new_n194));
  INV_X1    g008(.A(G101), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n188), .A2(new_n191), .A3(new_n195), .A4(new_n192), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n194), .A2(KEYINPUT4), .A3(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT4), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n193), .A2(new_n198), .A3(G101), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  XOR2_X1   g014(.A(KEYINPUT2), .B(G113), .Z(new_n201));
  XNOR2_X1  g015(.A(G116), .B(G119), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n202), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT68), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT68), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n201), .A2(new_n206), .A3(new_n202), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n203), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  OR2_X1    g022(.A1(new_n200), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G116), .ZN(new_n210));
  NOR3_X1   g024(.A1(new_n210), .A2(KEYINPUT5), .A3(G119), .ZN(new_n211));
  XOR2_X1   g025(.A(new_n211), .B(KEYINPUT80), .Z(new_n212));
  NAND2_X1  g026(.A1(new_n202), .A2(KEYINPUT5), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(G113), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n205), .A2(new_n207), .ZN(new_n215));
  INV_X1    g029(.A(new_n192), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n187), .A2(G107), .ZN(new_n217));
  OAI21_X1  g031(.A(G101), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AND2_X1   g032(.A1(new_n218), .A2(new_n196), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n214), .A2(new_n215), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n209), .A2(new_n220), .ZN(new_n221));
  XOR2_X1   g035(.A(G110), .B(G122), .Z(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT82), .B(KEYINPUT6), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n222), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n209), .A2(new_n220), .A3(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n223), .A2(KEYINPUT6), .A3(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT81), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n223), .A2(KEYINPUT81), .A3(KEYINPUT6), .A4(new_n227), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n225), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G146), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n233), .A2(G143), .ZN(new_n234));
  AND2_X1   g048(.A1(KEYINPUT64), .A2(G143), .ZN(new_n235));
  NOR2_X1   g049(.A1(KEYINPUT64), .A2(G143), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n234), .B1(new_n237), .B2(new_n233), .ZN(new_n238));
  XOR2_X1   g052(.A(KEYINPUT0), .B(G128), .Z(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT65), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT65), .ZN(new_n242));
  NOR3_X1   g056(.A1(new_n235), .A2(new_n236), .A3(G146), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n242), .B(new_n239), .C1(new_n243), .C2(new_n234), .ZN(new_n244));
  INV_X1    g058(.A(G143), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n245), .A2(G146), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT64), .B(G143), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n246), .B1(new_n247), .B2(G146), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n248), .A2(KEYINPUT0), .A3(G128), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n241), .A2(new_n244), .A3(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G125), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G224), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n253), .A2(G953), .ZN(new_n254));
  OAI21_X1  g068(.A(G146), .B1(new_n235), .B2(new_n236), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT1), .ZN(new_n256));
  INV_X1    g070(.A(new_n246), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n255), .A2(new_n256), .A3(G128), .A4(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G128), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n259), .B1(new_n257), .B2(KEYINPUT1), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n258), .B1(new_n238), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(new_n251), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  OR3_X1    g077(.A1(new_n252), .A2(new_n254), .A3(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n254), .B1(new_n252), .B2(new_n263), .ZN(new_n265));
  AND2_X1   g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(G902), .B1(new_n232), .B2(new_n266), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n264), .B(new_n265), .C1(KEYINPUT7), .C2(new_n254), .ZN(new_n268));
  OR4_X1    g082(.A1(KEYINPUT7), .A2(new_n252), .A3(new_n263), .A4(new_n254), .ZN(new_n269));
  XOR2_X1   g083(.A(new_n222), .B(KEYINPUT8), .Z(new_n270));
  INV_X1    g084(.A(new_n220), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n219), .B1(new_n214), .B2(new_n215), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n268), .A2(new_n269), .A3(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT83), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n268), .A2(new_n273), .A3(new_n269), .A4(KEYINPUT83), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n276), .A2(new_n277), .A3(new_n227), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n267), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(G210), .B1(G237), .B2(G902), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n267), .A2(new_n278), .A3(new_n280), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(G214), .B1(G237), .B2(G902), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n285), .B(KEYINPUT78), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n286), .B(KEYINPUT79), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n237), .A2(new_n233), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n259), .B1(new_n290), .B2(KEYINPUT1), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n258), .B1(new_n291), .B2(new_n248), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n219), .ZN(new_n293));
  OR2_X1    g107(.A1(new_n261), .A2(new_n219), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n293), .A2(new_n294), .A3(KEYINPUT77), .ZN(new_n295));
  INV_X1    g109(.A(G134), .ZN(new_n296));
  OAI21_X1  g110(.A(KEYINPUT11), .B1(new_n296), .B2(G137), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT11), .ZN(new_n298));
  INV_X1    g112(.A(G137), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n298), .A2(new_n299), .A3(G134), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n296), .A2(G137), .ZN(new_n302));
  INV_X1    g116(.A(G131), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(KEYINPUT66), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT66), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G131), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n301), .A2(new_n302), .A3(new_n307), .ZN(new_n308));
  AOI22_X1  g122(.A1(new_n297), .A2(new_n300), .B1(new_n296), .B2(G137), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n308), .B1(new_n303), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n261), .A2(new_n219), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT77), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n295), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT12), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n315), .B(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n261), .A2(KEYINPUT10), .A3(new_n219), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n318), .B1(new_n250), .B2(new_n200), .ZN(new_n319));
  AOI21_X1  g133(.A(KEYINPUT10), .B1(new_n292), .B2(new_n219), .ZN(new_n320));
  NOR3_X1   g134(.A1(new_n319), .A2(new_n320), .A3(new_n310), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(G110), .B(G140), .ZN(new_n323));
  INV_X1    g137(.A(G953), .ZN(new_n324));
  AND2_X1   g138(.A1(new_n324), .A2(G227), .ZN(new_n325));
  XOR2_X1   g139(.A(new_n323), .B(new_n325), .Z(new_n326));
  AND2_X1   g140(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n317), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n310), .B1(new_n319), .B2(new_n320), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n326), .B1(new_n322), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G469), .ZN(new_n333));
  INV_X1    g147(.A(G902), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n327), .A2(new_n329), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n315), .B(KEYINPUT12), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n337), .A2(new_n321), .ZN(new_n338));
  OAI211_X1 g152(.A(G469), .B(new_n336), .C1(new_n338), .C2(new_n326), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n333), .A2(new_n334), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n335), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  XOR2_X1   g156(.A(KEYINPUT9), .B(G234), .Z(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(G221), .B1(new_n344), .B2(G902), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT93), .ZN(new_n348));
  XNOR2_X1  g162(.A(G116), .B(G122), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT88), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n349), .B(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n190), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT91), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n245), .A2(G128), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n354), .B1(new_n247), .B2(G128), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n355), .B(new_n296), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT14), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n349), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n210), .A2(KEYINPUT14), .A3(G122), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(G107), .A3(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT91), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n351), .A2(new_n361), .A3(new_n190), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n353), .A2(new_n356), .A3(new_n360), .A4(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n355), .A2(KEYINPUT13), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n247), .A2(G128), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n365), .B(G134), .C1(KEYINPUT13), .C2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n354), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n368), .B1(new_n237), .B2(new_n259), .ZN(new_n369));
  OAI21_X1  g183(.A(KEYINPUT89), .B1(new_n369), .B2(G134), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT89), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n355), .A2(new_n371), .A3(new_n296), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n367), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT90), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n349), .B(KEYINPUT88), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G107), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n352), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n374), .A2(new_n375), .A3(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(new_n373), .A3(new_n367), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT90), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n364), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G217), .ZN(new_n383));
  NOR3_X1   g197(.A1(new_n344), .A2(new_n383), .A3(G953), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n384), .ZN(new_n386));
  AOI211_X1 g200(.A(new_n386), .B(new_n364), .C1(new_n379), .C2(new_n381), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n334), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G478), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n389), .A2(KEYINPUT15), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n348), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n375), .B1(new_n374), .B2(new_n378), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n380), .A2(KEYINPUT90), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n363), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n386), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n382), .A2(new_n384), .ZN(new_n396));
  AOI21_X1  g210(.A(G902), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n390), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n397), .A2(KEYINPUT93), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n391), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT92), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n401), .B1(new_n397), .B2(new_n398), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n388), .A2(KEYINPUT92), .A3(new_n390), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n324), .A2(G952), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n406), .B1(G234), .B2(G237), .ZN(new_n407));
  XOR2_X1   g221(.A(KEYINPUT21), .B(G898), .Z(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(G234), .A2(G237), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n410), .A2(G902), .A3(G953), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n407), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  NOR3_X1   g227(.A1(new_n251), .A2(KEYINPUT16), .A3(G140), .ZN(new_n414));
  INV_X1    g228(.A(G140), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n415), .B1(new_n251), .B2(KEYINPUT75), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT75), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n417), .A2(G125), .A3(G140), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n414), .B1(new_n419), .B2(KEYINPUT16), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n420), .A2(G146), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n420), .A2(G146), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(G237), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT71), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT71), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(G237), .ZN(new_n427));
  AOI21_X1  g241(.A(G953), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(G214), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n237), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n428), .A2(new_n245), .A3(G214), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n433), .A2(KEYINPUT17), .A3(new_n304), .A4(new_n306), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n432), .B(new_n307), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n423), .B(new_n434), .C1(new_n435), .C2(KEYINPUT17), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT18), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n437), .A2(new_n303), .ZN(new_n438));
  OAI21_X1  g252(.A(KEYINPUT85), .B1(new_n433), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n433), .A2(new_n438), .ZN(new_n440));
  XNOR2_X1  g254(.A(G125), .B(G140), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n233), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n442), .B1(new_n233), .B2(new_n419), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT85), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n432), .B(new_n444), .C1(new_n437), .C2(new_n303), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n439), .A2(new_n440), .A3(new_n443), .A4(new_n445), .ZN(new_n446));
  XNOR2_X1  g260(.A(G113), .B(G122), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n447), .B(new_n187), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n436), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n448), .B1(new_n436), .B2(new_n446), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n334), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(G475), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n420), .A2(G146), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT19), .ZN(new_n455));
  AOI21_X1  g269(.A(KEYINPUT86), .B1(new_n441), .B2(new_n455), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n419), .A2(new_n455), .ZN(new_n457));
  MUX2_X1   g271(.A(new_n456), .B(KEYINPUT86), .S(new_n457), .Z(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n233), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n435), .A2(new_n454), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n446), .ZN(new_n461));
  INV_X1    g275(.A(new_n448), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n449), .ZN(new_n464));
  NOR2_X1   g278(.A1(G475), .A2(G902), .ZN(new_n465));
  XOR2_X1   g279(.A(new_n465), .B(KEYINPUT87), .Z(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n468), .A2(KEYINPUT20), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT84), .B(KEYINPUT20), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n471), .B1(new_n464), .B2(new_n467), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n453), .B1(new_n469), .B2(new_n472), .ZN(new_n473));
  NOR3_X1   g287(.A1(new_n405), .A2(new_n413), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n289), .A2(new_n347), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n296), .A2(KEYINPUT67), .A3(G137), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n299), .A2(G134), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(KEYINPUT67), .B1(new_n296), .B2(G137), .ZN(new_n480));
  OAI21_X1  g294(.A(G131), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n308), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT69), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n308), .A2(new_n481), .A3(KEYINPUT69), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(new_n261), .A3(new_n485), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n310), .A2(new_n241), .A3(new_n244), .A4(new_n249), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n486), .A2(new_n208), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n261), .A2(new_n308), .A3(new_n481), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT30), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT70), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n486), .A2(KEYINPUT30), .A3(new_n487), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n486), .A2(KEYINPUT70), .A3(KEYINPUT30), .A4(new_n487), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n208), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n489), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  XNOR2_X1  g314(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n501), .B(G101), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n428), .A2(G210), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n502), .B(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(KEYINPUT73), .B1(new_n500), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT73), .ZN(new_n506));
  INV_X1    g320(.A(new_n504), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n208), .B1(new_n496), .B2(new_n497), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n506), .B(new_n507), .C1(new_n508), .C2(new_n489), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n488), .A2(KEYINPUT28), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT28), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n486), .A2(new_n511), .A3(new_n208), .A4(new_n487), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n491), .A2(new_n499), .ZN(new_n514));
  AND2_X1   g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(KEYINPUT29), .B1(new_n515), .B2(new_n504), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n505), .A2(new_n509), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n486), .A2(new_n487), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n499), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n513), .A2(KEYINPUT29), .A3(new_n504), .A4(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n517), .A2(new_n334), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(G472), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n488), .A2(new_n504), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n523), .B1(new_n498), .B2(new_n499), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT31), .ZN(new_n525));
  OAI21_X1  g339(.A(KEYINPUT72), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n504), .B1(new_n513), .B2(new_n514), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n527), .B1(new_n524), .B2(new_n525), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT72), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n529), .B(KEYINPUT31), .C1(new_n508), .C2(new_n523), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n526), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  NOR2_X1   g345(.A1(G472), .A2(G902), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT32), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n531), .A2(KEYINPUT32), .A3(new_n532), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n522), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(KEYINPUT74), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT74), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n522), .A2(new_n535), .A3(new_n539), .A4(new_n536), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n259), .A2(G119), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(KEYINPUT23), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n259), .A2(G119), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n545), .A2(new_n542), .ZN(new_n547));
  XOR2_X1   g361(.A(KEYINPUT24), .B(G110), .Z(new_n548));
  OAI22_X1  g362(.A1(new_n546), .A2(G110), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n549), .A2(new_n454), .A3(new_n442), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n546), .A2(G110), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n547), .A2(new_n548), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n551), .B(new_n552), .C1(new_n421), .C2(new_n422), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n324), .A2(G221), .A3(G234), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n555), .B(KEYINPUT22), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n556), .B(G137), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n554), .B(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  OR3_X1    g373(.A1(new_n559), .A2(KEYINPUT25), .A3(G902), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n383), .B1(G234), .B2(new_n334), .ZN(new_n561));
  OAI21_X1  g375(.A(KEYINPUT25), .B1(new_n559), .B2(G902), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n561), .A2(G902), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n558), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(KEYINPUT76), .B1(new_n541), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT76), .ZN(new_n569));
  AOI211_X1 g383(.A(new_n569), .B(new_n566), .C1(new_n538), .C2(new_n540), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n476), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(G101), .ZN(G3));
  NAND2_X1  g386(.A1(new_n531), .A2(new_n334), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT94), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(G472), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n573), .B(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n576), .A2(new_n567), .A3(new_n347), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(KEYINPUT95), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n389), .A2(new_n334), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT96), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n394), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n395), .A2(new_n581), .A3(KEYINPUT33), .A4(new_n396), .ZN(new_n582));
  OAI21_X1  g396(.A(KEYINPUT33), .B1(new_n382), .B2(KEYINPUT96), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n583), .B1(new_n385), .B2(new_n387), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n579), .B1(new_n585), .B2(G478), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n397), .A2(new_n389), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n473), .ZN(new_n589));
  INV_X1    g403(.A(new_n286), .ZN(new_n590));
  INV_X1    g404(.A(new_n413), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n284), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n578), .A2(new_n589), .A3(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(KEYINPUT34), .B(G104), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n593), .B(new_n594), .ZN(G6));
  AOI22_X1  g409(.A1(new_n391), .A2(new_n399), .B1(new_n402), .B2(new_n403), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n468), .A2(new_n470), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT97), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n464), .A2(new_n471), .A3(new_n467), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  AOI211_X1 g414(.A(new_n470), .B(new_n466), .C1(new_n463), .C2(new_n449), .ZN(new_n601));
  OAI21_X1  g415(.A(KEYINPUT97), .B1(new_n472), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n600), .A2(new_n602), .A3(new_n453), .ZN(new_n603));
  NOR3_X1   g417(.A1(new_n592), .A2(new_n596), .A3(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n578), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(KEYINPUT35), .B(G107), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(G9));
  INV_X1    g422(.A(new_n576), .ZN(new_n609));
  INV_X1    g423(.A(new_n557), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n610), .A2(KEYINPUT36), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n554), .B(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n564), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n563), .A2(new_n613), .ZN(new_n614));
  NOR3_X1   g428(.A1(new_n475), .A2(new_n609), .A3(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(KEYINPUT37), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(G110), .ZN(G12));
  INV_X1    g431(.A(new_n614), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n286), .B1(new_n282), .B2(new_n283), .ZN(new_n619));
  INV_X1    g433(.A(new_n407), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n620), .B1(G900), .B2(new_n411), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n600), .A2(new_n602), .A3(new_n453), .A4(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n622), .A2(new_n596), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n619), .A2(new_n623), .A3(new_n347), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n541), .A2(new_n618), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(G128), .ZN(G30));
  AND3_X1   g440(.A1(new_n531), .A2(KEYINPUT32), .A3(new_n532), .ZN(new_n627));
  AOI21_X1  g441(.A(KEYINPUT32), .B1(new_n531), .B2(new_n532), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n504), .B1(new_n519), .B2(new_n488), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n334), .B1(new_n524), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(G472), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n405), .A2(new_n473), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n634), .A2(new_n286), .A3(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(new_n621), .B(KEYINPUT98), .Z(new_n637));
  XOR2_X1   g451(.A(new_n637), .B(KEYINPUT39), .Z(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n347), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n640), .A2(KEYINPUT40), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n641), .A2(new_n618), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n284), .B(KEYINPUT38), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n640), .A2(KEYINPUT40), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n636), .A2(new_n642), .A3(new_n643), .A4(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(new_n237), .ZN(G45));
  NAND2_X1  g460(.A1(new_n284), .A2(new_n590), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n647), .A2(new_n346), .ZN(new_n648));
  AND4_X1   g462(.A1(new_n473), .A2(new_n586), .A3(new_n587), .A4(new_n621), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n541), .A2(new_n618), .A3(new_n648), .A4(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(G146), .ZN(G48));
  AOI21_X1  g465(.A(new_n566), .B1(new_n538), .B2(new_n540), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n592), .A2(new_n589), .ZN(new_n653));
  INV_X1    g467(.A(new_n345), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n330), .B1(new_n317), .B2(new_n327), .ZN(new_n655));
  OAI21_X1  g469(.A(G469), .B1(new_n655), .B2(G902), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT99), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n335), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  OAI211_X1 g472(.A(KEYINPUT99), .B(G469), .C1(new_n655), .C2(G902), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n654), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(KEYINPUT100), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n652), .A2(new_n653), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(KEYINPUT41), .B(G113), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G15));
  NAND3_X1  g478(.A1(new_n652), .A2(new_n604), .A3(new_n661), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G116), .ZN(G18));
  AOI21_X1  g480(.A(new_n614), .B1(new_n538), .B2(new_n540), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n619), .A2(new_n660), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n667), .A2(new_n474), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G119), .ZN(G21));
  INV_X1    g485(.A(new_n473), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n592), .A2(new_n596), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n573), .A2(G472), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n524), .A2(new_n525), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n513), .A2(new_n519), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n507), .B1(new_n676), .B2(KEYINPUT101), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n676), .A2(KEYINPUT101), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n675), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n524), .A2(new_n525), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n532), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  AND3_X1   g495(.A1(new_n674), .A2(new_n567), .A3(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n673), .A2(new_n661), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G122), .ZN(G24));
  NAND4_X1  g498(.A1(new_n649), .A2(new_n681), .A3(new_n618), .A4(new_n674), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n668), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(new_n251), .ZN(G27));
  NAND3_X1  g501(.A1(new_n282), .A2(new_n283), .A3(new_n590), .ZN(new_n688));
  AND3_X1   g502(.A1(new_n342), .A2(KEYINPUT102), .A3(new_n345), .ZN(new_n689));
  AOI21_X1  g503(.A(KEYINPUT102), .B1(new_n342), .B2(new_n345), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n652), .A2(new_n649), .A3(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT42), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n536), .B(KEYINPUT103), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n695), .A2(new_n535), .A3(new_n522), .ZN(new_n696));
  AND2_X1   g510(.A1(new_n696), .A2(new_n567), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n697), .A2(KEYINPUT42), .A3(new_n649), .A4(new_n691), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G131), .ZN(G33));
  NAND3_X1  g514(.A1(new_n652), .A2(new_n623), .A3(new_n691), .ZN(new_n701));
  XNOR2_X1  g515(.A(KEYINPUT104), .B(G134), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G36));
  NAND2_X1  g517(.A1(new_n588), .A2(new_n672), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT43), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n588), .A2(KEYINPUT43), .A3(new_n672), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n708), .A2(new_n609), .A3(new_n618), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n688), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n708), .A2(KEYINPUT44), .A3(new_n609), .A4(new_n618), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT105), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT46), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n336), .B1(new_n338), .B2(new_n326), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT45), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  OAI211_X1 g534(.A(KEYINPUT45), .B(new_n336), .C1(new_n338), .C2(new_n326), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n720), .A2(new_n721), .A3(G469), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n717), .B1(new_n723), .B2(new_n340), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n722), .A2(KEYINPUT46), .A3(new_n341), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n724), .A2(new_n335), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n345), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n727), .A2(new_n638), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n711), .A2(KEYINPUT105), .A3(new_n712), .A4(new_n713), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n716), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G137), .ZN(G39));
  INV_X1    g545(.A(KEYINPUT47), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n727), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n726), .A2(KEYINPUT47), .A3(new_n345), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n541), .A2(new_n567), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n735), .A2(new_n649), .A3(new_n712), .A4(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G140), .ZN(G42));
  NAND2_X1  g552(.A1(new_n658), .A2(new_n659), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT49), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n287), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OR4_X1    g555(.A1(new_n566), .A2(new_n741), .A3(new_n704), .A4(new_n654), .ZN(new_n742));
  INV_X1    g556(.A(new_n739), .ZN(new_n743));
  OAI22_X1  g557(.A1(new_n742), .A2(KEYINPUT106), .B1(KEYINPUT49), .B2(new_n743), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n742), .A2(KEYINPUT106), .ZN(new_n745));
  OR4_X1    g559(.A1(new_n643), .A2(new_n744), .A3(new_n745), .A4(new_n633), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n620), .B1(new_n706), .B2(new_n707), .ZN(new_n747));
  AND2_X1   g561(.A1(new_n747), .A2(new_n682), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT109), .ZN(new_n749));
  INV_X1    g563(.A(new_n660), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n749), .B1(new_n750), .B2(new_n590), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n750), .A2(new_n749), .A3(new_n590), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n643), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n748), .A2(new_n751), .A3(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT50), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n748), .A2(new_n753), .A3(KEYINPUT50), .A4(new_n751), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n743), .A2(new_n345), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n712), .B(new_n748), .C1(new_n735), .C2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n758), .A2(new_n760), .A3(KEYINPUT110), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(KEYINPUT51), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n750), .A2(new_n688), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n747), .A2(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n764), .A2(new_n618), .A3(new_n674), .A4(new_n681), .ZN(new_n765));
  AND4_X1   g579(.A1(new_n567), .A2(new_n634), .A3(new_n407), .A4(new_n763), .ZN(new_n766));
  INV_X1    g580(.A(new_n588), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n766), .A2(new_n672), .A3(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n758), .A2(new_n760), .A3(new_n765), .A4(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n406), .B1(new_n762), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n748), .A2(new_n669), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n766), .A2(new_n473), .A3(new_n588), .ZN(new_n772));
  AND3_X1   g586(.A1(new_n758), .A2(new_n760), .A3(new_n765), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n773), .A2(KEYINPUT51), .A3(new_n761), .A4(new_n768), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n770), .A2(new_n771), .A3(new_n772), .A4(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n764), .A2(new_n697), .ZN(new_n776));
  XOR2_X1   g590(.A(new_n776), .B(KEYINPUT48), .Z(new_n777));
  NOR2_X1   g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT111), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n596), .A2(new_n473), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n781), .B1(new_n473), .B2(new_n588), .ZN(new_n782));
  NOR4_X1   g596(.A1(new_n577), .A2(new_n782), .A3(new_n288), .A4(new_n413), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n539), .B1(new_n629), .B2(new_n522), .ZN(new_n784));
  INV_X1    g598(.A(new_n540), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n567), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n569), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n652), .A2(KEYINPUT76), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n783), .B1(new_n789), .B2(new_n476), .ZN(new_n790));
  AND4_X1   g604(.A1(new_n662), .A2(new_n665), .A3(new_n670), .A4(new_n683), .ZN(new_n791));
  INV_X1    g605(.A(new_n615), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n667), .A2(new_n596), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n622), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n794), .A2(new_n347), .A3(new_n795), .A4(new_n712), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n790), .A2(new_n791), .A3(new_n792), .A4(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n618), .A2(new_n674), .A3(new_n681), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n691), .A2(new_n649), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n699), .B(new_n701), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n797), .A2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n686), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n647), .A2(new_n635), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n614), .A2(new_n342), .A3(new_n345), .A4(new_n621), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT107), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n804), .A2(new_n805), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n803), .A2(new_n633), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n650), .A2(new_n625), .A3(new_n802), .A4(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT108), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n686), .B1(new_n667), .B2(new_n624), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n812), .A2(KEYINPUT108), .A3(new_n650), .A4(new_n808), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(KEYINPUT52), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT52), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n811), .A2(new_n816), .A3(new_n813), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n801), .A2(new_n818), .A3(KEYINPUT53), .ZN(new_n819));
  INV_X1    g633(.A(new_n783), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n571), .A2(new_n792), .A3(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n701), .B1(new_n798), .B2(new_n799), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n823), .B1(new_n694), .B2(new_n698), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n822), .A2(new_n824), .A3(new_n791), .A4(new_n796), .ZN(new_n825));
  OR2_X1    g639(.A1(new_n809), .A2(new_n816), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n825), .B1(new_n817), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n819), .B1(new_n827), .B2(KEYINPUT53), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(KEYINPUT54), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n811), .A2(new_n816), .A3(new_n813), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n816), .B1(new_n811), .B2(new_n813), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n830), .B1(new_n833), .B2(new_n825), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT54), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n817), .A2(new_n826), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n801), .A2(KEYINPUT53), .A3(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n834), .A2(new_n835), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n829), .A2(new_n838), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n775), .A2(KEYINPUT111), .A3(new_n777), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n780), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(G952), .A2(G953), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n746), .B1(new_n841), .B2(new_n842), .ZN(G75));
  NOR2_X1   g657(.A1(new_n324), .A2(G952), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n334), .B1(new_n834), .B2(new_n837), .ZN(new_n846));
  AOI21_X1  g660(.A(KEYINPUT56), .B1(new_n846), .B2(G210), .ZN(new_n847));
  XOR2_X1   g661(.A(new_n232), .B(new_n266), .Z(new_n848));
  XNOR2_X1  g662(.A(new_n848), .B(KEYINPUT112), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(KEYINPUT55), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n845), .B1(new_n847), .B2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT113), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n846), .B(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(new_n281), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT56), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n850), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n851), .B1(new_n854), .B2(new_n856), .ZN(G51));
  AOI21_X1  g671(.A(KEYINPUT53), .B1(new_n801), .B2(new_n818), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n665), .A2(new_n662), .A3(new_n670), .A4(new_n683), .ZN(new_n859));
  NOR4_X1   g673(.A1(new_n793), .A2(new_n346), .A3(new_n622), .A4(new_n688), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n821), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  AND4_X1   g675(.A1(KEYINPUT53), .A2(new_n836), .A3(new_n861), .A4(new_n824), .ZN(new_n862));
  OAI21_X1  g676(.A(KEYINPUT54), .B1(new_n858), .B2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT115), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n863), .A2(new_n864), .A3(new_n838), .ZN(new_n865));
  XOR2_X1   g679(.A(KEYINPUT114), .B(KEYINPUT57), .Z(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(new_n340), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n834), .A2(new_n837), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n868), .A2(KEYINPUT115), .A3(KEYINPUT54), .ZN(new_n869));
  OR2_X1    g683(.A1(new_n866), .A2(new_n340), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n865), .A2(new_n867), .A3(new_n869), .A4(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(new_n332), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n853), .A2(new_n723), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n844), .B1(new_n872), .B2(new_n873), .ZN(G54));
  OR2_X1    g688(.A1(new_n846), .A2(KEYINPUT113), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n846), .A2(KEYINPUT113), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n875), .A2(KEYINPUT58), .A3(G475), .A4(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(new_n464), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n853), .A2(KEYINPUT58), .A3(G475), .A4(new_n464), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n879), .A2(new_n880), .A3(new_n845), .ZN(G60));
  INV_X1    g695(.A(new_n585), .ZN(new_n882));
  XNOR2_X1  g696(.A(KEYINPUT116), .B(KEYINPUT59), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(new_n579), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n865), .A2(new_n869), .A3(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT117), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n886), .A2(new_n887), .A3(new_n845), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n887), .B1(new_n886), .B2(new_n845), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n882), .B1(new_n839), .B2(new_n884), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(G63));
  XNOR2_X1  g705(.A(KEYINPUT118), .B(KEYINPUT60), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n383), .A2(new_n334), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n892), .B(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n868), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n844), .B1(new_n895), .B2(new_n559), .ZN(new_n896));
  OR2_X1    g710(.A1(KEYINPUT119), .A2(KEYINPUT61), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n868), .A2(new_n612), .A3(new_n894), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(KEYINPUT119), .A2(KEYINPUT61), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n899), .B(new_n900), .ZN(G66));
  OAI21_X1  g715(.A(G953), .B1(new_n409), .B2(new_n253), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n822), .A2(new_n791), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT120), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n902), .B1(new_n904), .B2(G953), .ZN(new_n905));
  INV_X1    g719(.A(new_n232), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n906), .B1(G898), .B2(new_n324), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n905), .B(new_n907), .ZN(G69));
  AOI21_X1  g722(.A(new_n324), .B1(G227), .B2(G900), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT122), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n728), .A2(new_n697), .A3(new_n803), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(KEYINPUT121), .Z(new_n913));
  NAND4_X1  g727(.A1(new_n913), .A2(new_n730), .A3(new_n699), .A4(new_n737), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n812), .A2(new_n650), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n701), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n911), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n730), .A2(new_n699), .A3(new_n737), .ZN(new_n918));
  INV_X1    g732(.A(new_n916), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n918), .A2(KEYINPUT122), .A3(new_n913), .A4(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n917), .A2(new_n920), .A3(new_n324), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n498), .B(new_n458), .ZN(new_n922));
  NAND2_X1  g736(.A1(G900), .A2(G953), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT123), .ZN(new_n925));
  INV_X1    g739(.A(new_n922), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n915), .A2(new_n645), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT62), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n730), .A2(new_n737), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n789), .A2(new_n347), .A3(new_n639), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n930), .A2(new_n688), .A3(new_n782), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n928), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n926), .B1(new_n932), .B2(G953), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n924), .A2(new_n925), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n925), .B1(new_n924), .B2(new_n933), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n910), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n924), .A2(new_n933), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(KEYINPUT123), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n924), .A2(new_n925), .A3(new_n933), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n938), .A2(new_n909), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n936), .A2(new_n940), .ZN(G72));
  NAND2_X1  g755(.A1(G472), .A2(G902), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT63), .Z(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n917), .A2(new_n920), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n944), .B1(new_n945), .B2(new_n904), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n500), .B(KEYINPUT125), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n946), .A2(new_n504), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n505), .A2(new_n509), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n943), .B1(new_n949), .B2(new_n524), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT126), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n828), .A2(new_n951), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT127), .Z(new_n953));
  AOI21_X1  g767(.A(new_n944), .B1(new_n932), .B2(new_n904), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(KEYINPUT124), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n504), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n947), .B1(new_n954), .B2(KEYINPUT124), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n845), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n948), .A2(new_n953), .A3(new_n958), .ZN(G57));
endmodule


