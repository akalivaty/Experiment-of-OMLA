//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 1 0 1 1 1 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 1 0 0 0 0 1 0 0 0 0 1 1 0 0 0 0 0 0 0 1 1 0 0 1 0 0 0 1 0 0 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:53 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n444, new_n445, new_n446, new_n450, new_n452,
    new_n456, new_n457, new_n458, new_n459, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n567, new_n569, new_n570, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n643, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1206, new_n1207, new_n1208,
    new_n1209;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  INV_X1    g018(.A(G2072), .ZN(new_n444));
  INV_X1    g019(.A(G2078), .ZN(new_n445));
  NOR2_X1   g020(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g021(.A1(new_n446), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g022(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g023(.A(G452), .Z(G391));
  NAND2_X1  g024(.A1(G94), .A2(G452), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT65), .ZN(G173));
  NAND2_X1  g026(.A1(G7), .A2(G661), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g028(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g029(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g030(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT2), .Z(new_n457));
  NOR4_X1   g032(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n457), .A2(new_n459), .ZN(G325));
  INV_X1    g035(.A(G325), .ZN(G261));
  AOI22_X1  g036(.A1(new_n457), .A2(G2106), .B1(G567), .B2(new_n459), .ZN(new_n462));
  XOR2_X1   g037(.A(new_n462), .B(KEYINPUT66), .Z(G319));
  AND2_X1   g038(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n466), .A2(new_n467), .A3(G137), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(KEYINPUT3), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT3), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G2104), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n475), .A2(new_n477), .A3(G125), .ZN(new_n478));
  NAND2_X1  g053(.A1(G113), .A2(G2104), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n466), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n473), .A2(new_n480), .ZN(G160));
  NOR2_X1   g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT69), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n466), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT68), .ZN(new_n485));
  AND2_X1   g060(.A1(new_n467), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n467), .A2(new_n485), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n469), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(G136), .ZN(new_n489));
  INV_X1    g064(.A(G124), .ZN(new_n490));
  OAI22_X1  g065(.A1(new_n486), .A2(new_n487), .B1(new_n465), .B2(new_n464), .ZN(new_n491));
  OAI221_X1 g066(.A(new_n484), .B1(new_n488), .B2(new_n489), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  AND2_X1   g068(.A1(G126), .A2(G2105), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n467), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT70), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G2105), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n496), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n469), .A2(G114), .ZN(new_n502));
  NOR3_X1   g077(.A1(new_n502), .A2(new_n497), .A3(KEYINPUT70), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n495), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n466), .A2(new_n467), .A3(G138), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n506), .A2(KEYINPUT71), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n507), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n466), .A2(new_n467), .A3(new_n509), .A4(G138), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n504), .B1(new_n508), .B2(new_n510), .ZN(G164));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  OAI21_X1  g087(.A(KEYINPUT73), .B1(new_n512), .B2(KEYINPUT5), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT73), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n514), .A2(new_n515), .A3(G543), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n513), .A2(new_n516), .B1(KEYINPUT5), .B2(new_n512), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT74), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT72), .A2(G651), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT6), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n519), .B(new_n520), .ZN(new_n521));
  AND3_X1   g096(.A1(new_n517), .A2(new_n518), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n518), .B1(new_n517), .B2(new_n521), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G88), .ZN(new_n525));
  NAND2_X1  g100(.A1(G75), .A2(G543), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT75), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n513), .A2(new_n516), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n512), .A2(KEYINPUT5), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(G62), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n527), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  AND2_X1   g107(.A1(new_n521), .A2(G543), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n532), .A2(G651), .B1(new_n533), .B2(G50), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n525), .A2(new_n534), .ZN(G303));
  INV_X1    g110(.A(G303), .ZN(G166));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(KEYINPUT7), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n537), .A2(KEYINPUT7), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n533), .A2(G51), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n530), .A2(KEYINPUT76), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT76), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n517), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n541), .A2(G63), .A3(new_n543), .A4(G651), .ZN(new_n544));
  AND2_X1   g119(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n524), .A2(G89), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(G286));
  INV_X1    g122(.A(G286), .ZN(G168));
  INV_X1    g123(.A(G651), .ZN(new_n549));
  NAND2_X1  g124(.A1(G77), .A2(G543), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n541), .A2(new_n543), .ZN(new_n551));
  INV_X1    g126(.A(G64), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n549), .B1(new_n553), .B2(KEYINPUT77), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n554), .B1(KEYINPUT77), .B2(new_n553), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n524), .A2(G90), .B1(G52), .B2(new_n533), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(new_n556), .ZN(G301));
  INV_X1    g132(.A(G301), .ZN(G171));
  XNOR2_X1  g133(.A(KEYINPUT78), .B(G81), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n524), .A2(new_n559), .B1(G43), .B2(new_n533), .ZN(new_n560));
  AND3_X1   g135(.A1(new_n541), .A2(G56), .A3(new_n543), .ZN(new_n561));
  AND2_X1   g136(.A1(G68), .A2(G543), .ZN(new_n562));
  OAI21_X1  g137(.A(G651), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(G153));
  AND3_X1   g141(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G36), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n567), .A2(new_n570), .ZN(G188));
  AND3_X1   g146(.A1(new_n521), .A2(G53), .A3(G543), .ZN(new_n572));
  XOR2_X1   g147(.A(new_n572), .B(KEYINPUT9), .Z(new_n573));
  INV_X1    g148(.A(G91), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n517), .A2(new_n521), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(KEYINPUT74), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n517), .A2(new_n518), .A3(new_n521), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n573), .B1(new_n574), .B2(new_n578), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n517), .B(KEYINPUT79), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(G65), .ZN(new_n581));
  NAND2_X1  g156(.A1(G78), .A2(G543), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n549), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  OR2_X1    g158(.A1(new_n579), .A2(new_n583), .ZN(G299));
  AND3_X1   g159(.A1(new_n521), .A2(G49), .A3(G543), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n585), .B1(new_n524), .B2(G87), .ZN(new_n586));
  AOI21_X1  g161(.A(G74), .B1(new_n541), .B2(new_n543), .ZN(new_n587));
  NOR3_X1   g162(.A1(new_n587), .A2(KEYINPUT80), .A3(new_n549), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT80), .ZN(new_n589));
  INV_X1    g164(.A(G74), .ZN(new_n590));
  AND3_X1   g165(.A1(new_n528), .A2(new_n542), .A3(new_n529), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n542), .B1(new_n528), .B2(new_n529), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n589), .B1(new_n593), .B2(G651), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n586), .B1(new_n588), .B2(new_n594), .ZN(G288));
  INV_X1    g170(.A(KEYINPUT81), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n517), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n597), .B2(new_n549), .ZN(new_n598));
  NAND2_X1  g173(.A1(G73), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G61), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n530), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n601), .A2(KEYINPUT81), .A3(G651), .ZN(new_n602));
  AND3_X1   g177(.A1(new_n598), .A2(new_n602), .A3(KEYINPUT82), .ZN(new_n603));
  AOI21_X1  g178(.A(KEYINPUT82), .B1(new_n598), .B2(new_n602), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n533), .A2(G48), .ZN(new_n606));
  INV_X1    g181(.A(G86), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n578), .B2(new_n607), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(G305));
  AOI22_X1  g185(.A1(new_n524), .A2(G85), .B1(G47), .B2(new_n533), .ZN(new_n611));
  AND3_X1   g186(.A1(new_n541), .A2(G60), .A3(new_n543), .ZN(new_n612));
  AND2_X1   g187(.A1(G72), .A2(G543), .ZN(new_n613));
  OAI21_X1  g188(.A(G651), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n611), .A2(new_n614), .ZN(G290));
  NAND2_X1  g190(.A1(G301), .A2(G868), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n517), .A2(KEYINPUT79), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n517), .A2(KEYINPUT79), .ZN(new_n619));
  OAI21_X1  g194(.A(G66), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(G79), .A2(G543), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n549), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n533), .A2(G54), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(KEYINPUT83), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(KEYINPUT83), .ZN(new_n626));
  AOI22_X1  g201(.A1(new_n580), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n626), .B(new_n623), .C1(new_n627), .C2(new_n549), .ZN(new_n628));
  INV_X1    g203(.A(G92), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n578), .A2(new_n629), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n630), .A2(KEYINPUT10), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(KEYINPUT10), .ZN(new_n632));
  AOI22_X1  g207(.A1(new_n625), .A2(new_n628), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n616), .B1(G868), .B2(new_n633), .ZN(G284));
  OAI21_X1  g209(.A(new_n616), .B1(G868), .B2(new_n633), .ZN(G321));
  NAND2_X1  g210(.A1(G286), .A2(G868), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n636), .A2(KEYINPUT84), .ZN(new_n637));
  INV_X1    g212(.A(G868), .ZN(new_n638));
  NAND2_X1  g213(.A1(G299), .A2(new_n638), .ZN(new_n639));
  AND2_X1   g214(.A1(new_n636), .A2(KEYINPUT84), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n637), .B1(new_n639), .B2(new_n640), .ZN(G297));
  AOI21_X1  g216(.A(new_n637), .B1(new_n639), .B2(new_n640), .ZN(G280));
  INV_X1    g217(.A(G559), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n633), .B1(new_n643), .B2(G860), .ZN(G148));
  NAND2_X1  g219(.A1(new_n564), .A2(new_n638), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n625), .A2(new_n628), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n631), .A2(new_n632), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n648), .A2(G559), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n645), .B1(new_n649), .B2(new_n638), .ZN(G323));
  XNOR2_X1  g225(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI221_X1 g226(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n466), .C2(G111), .ZN(new_n652));
  INV_X1    g227(.A(G123), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n652), .B1(new_n491), .B2(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n488), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n654), .B1(G135), .B2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT85), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n657), .A2(G2096), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(G2096), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n467), .A2(new_n471), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT12), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT13), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G2100), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n658), .A2(new_n659), .A3(new_n663), .ZN(G156));
  XNOR2_X1  g239(.A(G2427), .B(G2438), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2430), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT15), .B(G2435), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n666), .A2(new_n667), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n668), .A2(KEYINPUT14), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2451), .B(G2454), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT16), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n670), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2443), .B(G2446), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1341), .B(G1348), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT86), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n678), .B(G14), .C1(new_n676), .C2(new_n675), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(G401));
  XNOR2_X1  g255(.A(G2072), .B(G2078), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT17), .Z(new_n682));
  XNOR2_X1  g257(.A(G2067), .B(G2678), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT87), .Z(new_n684));
  OR2_X1    g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G2084), .B(G2090), .Z(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n684), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n685), .B(new_n687), .C1(new_n688), .C2(new_n681), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(KEYINPUT88), .Z(new_n690));
  NAND3_X1  g265(.A1(new_n686), .A2(new_n683), .A3(new_n681), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT18), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n688), .A2(new_n687), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n692), .B1(new_n693), .B2(new_n682), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(G2096), .B(G2100), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(G227));
  XOR2_X1   g272(.A(G1971), .B(G1976), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT19), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1956), .B(G2474), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1961), .B(G1966), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  NOR3_X1   g278(.A1(new_n699), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n699), .A2(new_n702), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT89), .B(KEYINPUT20), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  AOI211_X1 g282(.A(new_n704), .B(new_n707), .C1(new_n699), .C2(new_n703), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT90), .ZN(new_n709));
  XOR2_X1   g284(.A(G1981), .B(G1986), .Z(new_n710));
  XNOR2_X1  g285(.A(G1991), .B(G1996), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n709), .B(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(G229));
  INV_X1    g291(.A(G16), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G6), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(new_n609), .B2(new_n717), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT32), .B(G1981), .Z(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n576), .A2(G87), .A3(new_n577), .ZN(new_n722));
  INV_X1    g297(.A(new_n585), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(KEYINPUT80), .B1(new_n587), .B2(new_n549), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n593), .A2(new_n589), .A3(G651), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n724), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n727), .A2(new_n717), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n717), .B2(G23), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT33), .B(G1976), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n729), .A2(new_n730), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n717), .A2(G22), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G166), .B2(new_n717), .ZN(new_n734));
  INV_X1    g309(.A(G1971), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  AND4_X1   g311(.A1(new_n721), .A2(new_n731), .A3(new_n732), .A4(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT34), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n737), .A2(new_n738), .ZN(new_n740));
  OAI221_X1 g315(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n466), .C2(G107), .ZN(new_n741));
  INV_X1    g316(.A(G131), .ZN(new_n742));
  INV_X1    g317(.A(G119), .ZN(new_n743));
  OAI221_X1 g318(.A(new_n741), .B1(new_n488), .B2(new_n742), .C1(new_n743), .C2(new_n491), .ZN(new_n744));
  MUX2_X1   g319(.A(G25), .B(new_n744), .S(G29), .Z(new_n745));
  XOR2_X1   g320(.A(KEYINPUT35), .B(G1991), .Z(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(G1986), .ZN(new_n748));
  INV_X1    g323(.A(G290), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(G16), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G16), .B2(G24), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n747), .B1(new_n748), .B2(new_n751), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(new_n748), .B2(new_n751), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n739), .A2(new_n740), .A3(new_n753), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT91), .B(KEYINPUT36), .Z(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n467), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n757), .A2(new_n466), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT95), .Z(new_n759));
  NAND2_X1  g334(.A1(new_n655), .A2(G139), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT25), .Z(new_n762));
  NAND3_X1  g337(.A1(new_n759), .A2(new_n760), .A3(new_n762), .ZN(new_n763));
  MUX2_X1   g338(.A(G33), .B(new_n763), .S(G29), .Z(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(new_n444), .ZN(new_n765));
  INV_X1    g340(.A(G29), .ZN(new_n766));
  INV_X1    g341(.A(new_n491), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n767), .A2(G129), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n655), .A2(G141), .ZN(new_n769));
  NAND3_X1  g344(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT26), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n770), .A2(new_n771), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n772), .A2(new_n773), .B1(G105), .B2(new_n471), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n768), .A2(new_n769), .A3(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n776), .A2(new_n766), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n766), .B2(G32), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT27), .B(G1996), .ZN(new_n779));
  OAI221_X1 g354(.A(new_n765), .B1(new_n766), .B2(new_n657), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(G168), .A2(new_n717), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n717), .B2(G21), .ZN(new_n782));
  INV_X1    g357(.A(G1966), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT24), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n766), .B1(new_n785), .B2(G34), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(new_n785), .B2(G34), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G160), .B2(G29), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n788), .A2(G2084), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(G2084), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT31), .B(G11), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT30), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n792), .A2(G28), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT97), .Z(new_n794));
  OAI211_X1 g369(.A(new_n794), .B(new_n766), .C1(new_n792), .C2(G28), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n789), .A2(new_n790), .A3(new_n791), .A4(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n766), .A2(G27), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G164), .B2(new_n766), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G2078), .ZN(new_n799));
  NOR4_X1   g374(.A1(new_n780), .A2(new_n784), .A3(new_n796), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n717), .A2(G20), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT23), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n579), .A2(new_n583), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n802), .B1(new_n803), .B2(new_n717), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G1956), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n778), .A2(new_n779), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT96), .ZN(new_n807));
  AOI211_X1 g382(.A(new_n805), .B(new_n807), .C1(new_n783), .C2(new_n782), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n766), .A2(G35), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G162), .B2(new_n766), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT29), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(G2090), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n766), .A2(G26), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT28), .Z(new_n814));
  OAI221_X1 g389(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n466), .C2(G116), .ZN(new_n815));
  INV_X1    g390(.A(G140), .ZN(new_n816));
  INV_X1    g391(.A(G128), .ZN(new_n817));
  OAI221_X1 g392(.A(new_n815), .B1(new_n488), .B2(new_n816), .C1(new_n817), .C2(new_n491), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT93), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n818), .A2(new_n819), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n814), .B1(new_n822), .B2(G29), .ZN(new_n823));
  XNOR2_X1  g398(.A(KEYINPUT94), .B(G2067), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n812), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n717), .A2(G19), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(new_n565), .B2(new_n717), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(G1341), .Z(new_n829));
  NAND4_X1  g404(.A1(new_n800), .A2(new_n808), .A3(new_n826), .A4(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(G4), .A2(G16), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT92), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(new_n648), .B2(new_n717), .ZN(new_n833));
  INV_X1    g408(.A(G1348), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n717), .A2(G5), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(G171), .B2(new_n717), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(G1961), .ZN(new_n838));
  NOR3_X1   g413(.A1(new_n830), .A2(new_n835), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n756), .A2(new_n839), .ZN(G150));
  INV_X1    g415(.A(G150), .ZN(G311));
  NOR2_X1   g416(.A1(new_n648), .A2(new_n643), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT38), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n533), .A2(G55), .ZN(new_n844));
  INV_X1    g419(.A(G93), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n844), .B1(new_n578), .B2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(G67), .ZN(new_n847));
  NOR3_X1   g422(.A1(new_n591), .A2(new_n592), .A3(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(G80), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n849), .A2(new_n512), .ZN(new_n850));
  OAI21_X1  g425(.A(KEYINPUT98), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT98), .ZN(new_n852));
  INV_X1    g427(.A(new_n850), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n852), .B(new_n853), .C1(new_n551), .C2(new_n847), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n851), .A2(G651), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n846), .B1(new_n855), .B2(KEYINPUT99), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT99), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n851), .A2(new_n854), .A3(new_n857), .A4(G651), .ZN(new_n858));
  AND3_X1   g433(.A1(new_n856), .A2(new_n565), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n565), .B1(new_n856), .B2(new_n858), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n843), .B(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT39), .ZN(new_n863));
  AOI21_X1  g438(.A(G860), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n864), .B1(new_n863), .B2(new_n862), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n856), .A2(new_n858), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(G860), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n867), .B(KEYINPUT37), .Z(new_n868));
  NAND2_X1  g443(.A1(new_n865), .A2(new_n868), .ZN(G145));
  AND2_X1   g444(.A1(new_n820), .A2(new_n821), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(G164), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n508), .A2(new_n510), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n498), .A2(new_n496), .A3(new_n500), .ZN(new_n873));
  OAI21_X1  g448(.A(KEYINPUT70), .B1(new_n502), .B2(new_n497), .ZN(new_n874));
  AOI22_X1  g449(.A1(new_n873), .A2(new_n874), .B1(new_n467), .B2(new_n494), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n822), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n871), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(new_n776), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n871), .A2(new_n775), .A3(new_n877), .ZN(new_n880));
  OR2_X1    g455(.A1(new_n763), .A2(KEYINPUT100), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n763), .A2(KEYINPUT100), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n744), .B(KEYINPUT101), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(new_n661), .ZN(new_n887));
  OAI221_X1 g462(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n466), .C2(G118), .ZN(new_n888));
  INV_X1    g463(.A(G130), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n888), .B1(new_n491), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n890), .B1(G142), .B2(new_n655), .ZN(new_n891));
  XOR2_X1   g466(.A(new_n887), .B(new_n891), .Z(new_n892));
  NAND4_X1  g467(.A1(new_n879), .A2(new_n883), .A3(new_n880), .A4(new_n881), .ZN(new_n893));
  AND3_X1   g468(.A1(new_n885), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n892), .B1(new_n885), .B2(new_n893), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n657), .B(G160), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(G162), .ZN(new_n897));
  OR3_X1    g472(.A1(new_n894), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(G37), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n897), .B1(new_n894), .B2(new_n895), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g477(.A1(new_n866), .A2(new_n638), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n609), .B(G303), .ZN(new_n904));
  XNOR2_X1  g479(.A(G288), .B(G290), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(KEYINPUT102), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n905), .A2(KEYINPUT102), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n908), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n910), .A2(new_n906), .A3(new_n904), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  XOR2_X1   g487(.A(KEYINPUT103), .B(KEYINPUT42), .Z(new_n913));
  XNOR2_X1  g488(.A(new_n912), .B(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n861), .B(new_n649), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n648), .A2(G299), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n633), .A2(new_n803), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  AND3_X1   g494(.A1(new_n916), .A2(new_n917), .A3(KEYINPUT41), .ZN(new_n920));
  AOI21_X1  g495(.A(KEYINPUT41), .B1(new_n916), .B2(new_n917), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n919), .B1(new_n915), .B2(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n914), .B(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n903), .B1(new_n924), .B2(new_n638), .ZN(G295));
  OAI21_X1  g500(.A(new_n903), .B1(new_n924), .B2(new_n638), .ZN(G331));
  INV_X1    g501(.A(new_n918), .ZN(new_n927));
  OAI21_X1  g502(.A(G171), .B1(new_n859), .B2(new_n860), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n866), .A2(new_n564), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n856), .A2(new_n565), .A3(new_n858), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n929), .A2(G301), .A3(new_n930), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n928), .A2(new_n931), .A3(G168), .ZN(new_n932));
  AOI21_X1  g507(.A(G168), .B1(new_n928), .B2(new_n931), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n927), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n928), .A2(new_n931), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(G286), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n928), .A2(new_n931), .A3(G168), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n936), .A2(new_n922), .A3(new_n937), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n909), .A2(new_n911), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n934), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(new_n899), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n939), .B1(new_n934), .B2(new_n938), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT43), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n934), .A2(new_n938), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n912), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT43), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n945), .A2(new_n946), .A3(new_n899), .A4(new_n940), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT104), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n943), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n950));
  OAI211_X1 g525(.A(KEYINPUT104), .B(KEYINPUT43), .C1(new_n941), .C2(new_n942), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n943), .A2(new_n947), .A3(KEYINPUT44), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(G397));
  INV_X1    g529(.A(KEYINPUT105), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n478), .A2(new_n479), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n472), .B(new_n468), .C1(new_n956), .C2(new_n466), .ZN(new_n957));
  INV_X1    g532(.A(G40), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n955), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(G160), .A2(KEYINPUT105), .A3(G40), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT45), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n962), .B1(G164), .B2(G1384), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  XOR2_X1   g539(.A(new_n964), .B(KEYINPUT107), .Z(new_n965));
  INV_X1    g540(.A(G2067), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n870), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n822), .A2(G2067), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n965), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n965), .A2(G1996), .A3(new_n775), .ZN(new_n970));
  INV_X1    g545(.A(G1996), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n964), .A2(new_n971), .A3(new_n776), .ZN(new_n972));
  AND3_X1   g547(.A1(new_n969), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n746), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n744), .A2(new_n974), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n744), .A2(new_n974), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n965), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n973), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n749), .A2(new_n748), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n979), .B(KEYINPUT106), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n981), .B1(new_n748), .B2(new_n749), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n978), .B1(new_n964), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT54), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT105), .B1(G160), .B2(G40), .ZN(new_n985));
  NOR4_X1   g560(.A1(new_n473), .A2(new_n480), .A3(new_n955), .A4(new_n958), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G1384), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n876), .A2(KEYINPUT45), .A3(new_n988), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n987), .A2(new_n445), .A3(new_n963), .A4(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT53), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n445), .A2(KEYINPUT53), .ZN(new_n993));
  NOR3_X1   g568(.A1(new_n957), .A2(new_n958), .A3(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n963), .A2(new_n994), .A3(new_n989), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n992), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT50), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n997), .B1(new_n876), .B2(new_n988), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n961), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT108), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n1000), .B1(G164), .B2(G1384), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n876), .A2(KEYINPUT108), .A3(new_n988), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1001), .A2(new_n997), .A3(new_n1002), .ZN(new_n1003));
  AND3_X1   g578(.A1(new_n999), .A2(new_n1003), .A3(KEYINPUT117), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT117), .B1(new_n999), .B2(new_n1003), .ZN(new_n1005));
  NOR3_X1   g580(.A1(new_n1004), .A2(new_n1005), .A3(G1961), .ZN(new_n1006));
  OR2_X1    g581(.A1(new_n1006), .A2(KEYINPUT124), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(KEYINPUT124), .ZN(new_n1008));
  AOI211_X1 g583(.A(G171), .B(new_n996), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT123), .ZN(new_n1010));
  AND2_X1   g585(.A1(new_n987), .A2(new_n989), .ZN(new_n1011));
  AOI21_X1  g586(.A(KEYINPUT108), .B1(new_n876), .B2(new_n988), .ZN(new_n1012));
  AOI211_X1 g587(.A(new_n1000), .B(G1384), .C1(new_n872), .C2(new_n875), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1011), .B1(new_n1014), .B2(KEYINPUT45), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n992), .B1(new_n1015), .B2(new_n993), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1006), .A2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1010), .B1(new_n1017), .B2(G301), .ZN(new_n1018));
  OAI211_X1 g593(.A(KEYINPUT123), .B(G171), .C1(new_n1006), .C2(new_n1016), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n984), .B1(new_n1009), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n1022));
  INV_X1    g597(.A(G8), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1023), .B1(new_n1014), .B2(new_n987), .ZN(new_n1024));
  OAI211_X1 g599(.A(G1976), .B(new_n586), .C1(new_n588), .C2(new_n594), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1022), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n987), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1027), .A2(new_n1025), .A3(G8), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1022), .B1(new_n727), .B2(G1976), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1026), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G1981), .ZN(new_n1032));
  AOI22_X1  g607(.A1(new_n524), .A2(G86), .B1(G48), .B2(new_n533), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n1032), .B(new_n1033), .C1(new_n603), .C2(new_n604), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n598), .A2(new_n602), .ZN(new_n1035));
  OAI21_X1  g610(.A(G1981), .B1(new_n608), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT49), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1034), .A2(KEYINPUT49), .A3(new_n1036), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1039), .A2(new_n1040), .A3(new_n1024), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1031), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n987), .A2(new_n989), .ZN(new_n1043));
  INV_X1    g618(.A(new_n963), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n735), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(G2090), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n999), .A2(new_n1003), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(G8), .ZN(new_n1049));
  NAND2_X1  g624(.A1(G303), .A2(G8), .ZN(new_n1050));
  XNOR2_X1  g625(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n1051));
  XNOR2_X1  g626(.A(new_n1050), .B(new_n1051), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1049), .A2(new_n1052), .ZN(new_n1053));
  OR2_X1    g628(.A1(new_n1042), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT112), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n997), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1055), .B1(new_n1056), .B2(new_n961), .ZN(new_n1057));
  OAI21_X1  g632(.A(KEYINPUT50), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1058), .A2(KEYINPUT112), .A3(new_n987), .ZN(new_n1059));
  NOR2_X1   g634(.A1(G164), .A2(G1384), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(new_n997), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1057), .A2(new_n1059), .A3(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT113), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT113), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1057), .A2(new_n1059), .A3(new_n1064), .A4(new_n1061), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1063), .A2(new_n1046), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(new_n1045), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(G8), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1054), .B1(new_n1068), .B2(new_n1052), .ZN(new_n1069));
  AND2_X1   g644(.A1(new_n1006), .A2(KEYINPUT124), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1006), .A2(KEYINPUT124), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(G171), .B1(new_n1072), .B2(new_n996), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n984), .B1(new_n1017), .B2(G301), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT45), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n783), .B1(new_n1076), .B2(new_n1043), .ZN(new_n1077));
  INV_X1    g652(.A(G2084), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n999), .A2(new_n1003), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(G8), .ZN(new_n1081));
  NAND2_X1  g656(.A1(G286), .A2(G8), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1081), .A2(KEYINPUT51), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT51), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1084), .B(G8), .C1(new_n1080), .C2(G286), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1082), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT122), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  AOI211_X1 g663(.A(KEYINPUT122), .B(new_n1082), .C1(new_n1077), .C2(new_n1079), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1083), .B(new_n1085), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1021), .A2(new_n1069), .A3(new_n1075), .A4(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT61), .ZN(new_n1092));
  INV_X1    g667(.A(G1956), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1062), .A2(new_n1093), .ZN(new_n1094));
  XNOR2_X1  g669(.A(new_n803), .B(KEYINPUT57), .ZN(new_n1095));
  XNOR2_X1  g670(.A(KEYINPUT56), .B(G2072), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n1011), .A2(new_n963), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  AND4_X1   g673(.A1(KEYINPUT116), .A2(new_n1094), .A3(new_n1095), .A4(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1097), .B1(new_n1062), .B2(new_n1093), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT116), .B1(new_n1100), .B2(new_n1095), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT119), .ZN(new_n1103));
  XNOR2_X1  g678(.A(G299), .B(KEYINPUT57), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1058), .A2(new_n987), .ZN(new_n1105));
  AOI22_X1  g680(.A1(new_n1105), .A2(new_n1055), .B1(new_n997), .B2(new_n1060), .ZN(new_n1106));
  AOI21_X1  g681(.A(G1956), .B1(new_n1106), .B2(new_n1059), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1103), .B(new_n1104), .C1(new_n1107), .C2(new_n1097), .ZN(new_n1108));
  OAI21_X1  g683(.A(KEYINPUT119), .B1(new_n1100), .B2(new_n1095), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1092), .B1(new_n1102), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(KEYINPUT120), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT120), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1113), .B(new_n1092), .C1(new_n1102), .C2(new_n1110), .ZN(new_n1114));
  OR3_X1    g689(.A1(new_n1004), .A2(new_n1005), .A3(G1348), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1027), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(new_n966), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT60), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT121), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1118), .B1(new_n633), .B2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1115), .A2(new_n1117), .A3(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n633), .A2(new_n1119), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NOR3_X1   g698(.A1(new_n1004), .A2(new_n1005), .A3(G1348), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1117), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1118), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1122), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1127), .A2(new_n1120), .A3(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1123), .A2(new_n1126), .A3(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1104), .B1(new_n1107), .B2(new_n1097), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1100), .A2(new_n1095), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1131), .A2(KEYINPUT61), .A3(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1134));
  XNOR2_X1  g709(.A(KEYINPUT118), .B(KEYINPUT58), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n1135), .B(G1341), .ZN(new_n1136));
  AOI22_X1  g711(.A1(new_n1134), .A2(new_n971), .B1(new_n1027), .B2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1137), .A2(new_n564), .ZN(new_n1138));
  XOR2_X1   g713(.A(new_n1138), .B(KEYINPUT59), .Z(new_n1139));
  AND3_X1   g714(.A1(new_n1130), .A2(new_n1133), .A3(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1112), .A2(new_n1114), .A3(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1131), .B1(new_n648), .B2(new_n1127), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1142), .B1(new_n1101), .B2(new_n1099), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1091), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT125), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1147));
  OAI21_X1  g722(.A(KEYINPUT62), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n1086), .B(new_n1087), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT62), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1149), .A2(new_n1150), .A3(new_n1085), .A4(new_n1083), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1148), .A2(new_n1020), .A3(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1042), .A2(new_n1053), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1023), .B1(new_n1066), .B2(new_n1045), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1052), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1153), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1145), .B1(new_n1152), .B2(new_n1156), .ZN(new_n1157));
  AOI22_X1  g732(.A1(new_n1090), .A2(KEYINPUT62), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1069), .A2(new_n1158), .A3(KEYINPUT125), .A4(new_n1151), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1160));
  AND3_X1   g735(.A1(new_n1034), .A2(KEYINPUT49), .A3(new_n1036), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1024), .ZN(new_n1162));
  AOI21_X1  g737(.A(KEYINPUT49), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1163));
  NOR3_X1   g738(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1028), .A2(KEYINPUT52), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1165), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT110), .ZN(new_n1167));
  NOR3_X1   g742(.A1(new_n1164), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(KEYINPUT110), .B1(new_n1031), .B2(new_n1041), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1053), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  XOR2_X1   g745(.A(new_n1024), .B(KEYINPUT111), .Z(new_n1171));
  NOR3_X1   g746(.A1(new_n1164), .A2(G1976), .A3(G288), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1034), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1171), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1170), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1049), .A2(KEYINPUT114), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT114), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1048), .A2(new_n1177), .A3(G8), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1176), .A2(new_n1052), .A3(new_n1178), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1179), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT115), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  OAI211_X1 g757(.A(new_n1179), .B(KEYINPUT115), .C1(new_n1168), .C2(new_n1169), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT63), .ZN(new_n1184));
  NOR4_X1   g759(.A1(new_n1053), .A2(new_n1184), .A3(G286), .A4(new_n1081), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1182), .A2(new_n1183), .A3(new_n1185), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1081), .A2(G286), .ZN(new_n1187));
  OAI211_X1 g762(.A(new_n1153), .B(new_n1187), .C1(new_n1154), .C2(new_n1155), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1188), .A2(new_n1184), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1175), .B1(new_n1186), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1160), .A2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n983), .B1(new_n1144), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n965), .A2(new_n775), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n964), .A2(new_n971), .ZN(new_n1194));
  XNOR2_X1  g769(.A(new_n1194), .B(KEYINPUT46), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n969), .A2(new_n1193), .A3(new_n1195), .ZN(new_n1196));
  XNOR2_X1  g771(.A(new_n1196), .B(KEYINPUT47), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n980), .A2(new_n964), .ZN(new_n1198));
  XOR2_X1   g773(.A(new_n1198), .B(KEYINPUT48), .Z(new_n1199));
  OAI21_X1  g774(.A(new_n1197), .B1(new_n1199), .B2(new_n978), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n968), .B1(new_n973), .B2(new_n975), .ZN(new_n1201));
  XNOR2_X1  g776(.A(new_n1201), .B(KEYINPUT126), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1200), .B1(new_n1202), .B2(new_n965), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1192), .A2(new_n1203), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g779(.A(new_n462), .ZN(new_n1206));
  OR2_X1    g780(.A1(G227), .A2(new_n1206), .ZN(new_n1207));
  OAI21_X1  g781(.A(new_n715), .B1(new_n1207), .B2(KEYINPUT127), .ZN(new_n1208));
  AOI211_X1 g782(.A(new_n1208), .B(G401), .C1(KEYINPUT127), .C2(new_n1207), .ZN(new_n1209));
  NAND4_X1  g783(.A1(new_n949), .A2(new_n901), .A3(new_n1209), .A4(new_n951), .ZN(G225));
  INV_X1    g784(.A(G225), .ZN(G308));
endmodule


