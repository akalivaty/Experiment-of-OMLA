

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X2 U555 ( .A(G2105), .ZN(n545) );
  NOR2_X1 U556 ( .A1(n797), .A2(n701), .ZN(n738) );
  NOR2_X1 U557 ( .A1(n709), .A2(n967), .ZN(n708) );
  BUF_X1 U558 ( .A(n738), .Z(n732) );
  XNOR2_X1 U559 ( .A(n723), .B(n722), .ZN(n727) );
  INV_X1 U560 ( .A(KEYINPUT103), .ZN(n722) );
  BUF_X1 U561 ( .A(n709), .Z(n753) );
  AND2_X1 U562 ( .A1(n760), .A2(n759), .ZN(n761) );
  AND2_X1 U563 ( .A1(n989), .A2(n842), .ZN(n524) );
  NOR2_X1 U564 ( .A1(n829), .A2(n524), .ZN(n525) );
  XNOR2_X1 U565 ( .A(KEYINPUT98), .B(n763), .ZN(n526) );
  NOR2_X1 U566 ( .A1(n768), .A2(n791), .ZN(n527) );
  INV_X1 U567 ( .A(n997), .ZN(n710) );
  AND2_X1 U568 ( .A1(n711), .A2(n710), .ZN(n712) );
  AND2_X1 U569 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U570 ( .A(KEYINPUT104), .B(KEYINPUT30), .ZN(n742) );
  XNOR2_X1 U571 ( .A(n743), .B(n742), .ZN(n744) );
  NOR2_X1 U572 ( .A1(G168), .A2(n744), .ZN(n745) );
  XNOR2_X1 U573 ( .A(n731), .B(n730), .ZN(n737) );
  AND2_X1 U574 ( .A1(n764), .A2(n526), .ZN(n767) );
  NOR2_X1 U575 ( .A1(G2104), .A2(G2105), .ZN(n550) );
  NOR2_X2 U576 ( .A1(G2104), .A2(n545), .ZN(n901) );
  NOR2_X1 U577 ( .A1(n628), .A2(G651), .ZN(n657) );
  AND2_X2 U578 ( .A1(n545), .A2(G2104), .ZN(n904) );
  INV_X1 U579 ( .A(G651), .ZN(n532) );
  NOR2_X1 U580 ( .A1(G543), .A2(n532), .ZN(n528) );
  XOR2_X1 U581 ( .A(KEYINPUT1), .B(n528), .Z(n653) );
  NAND2_X1 U582 ( .A1(G63), .A2(n653), .ZN(n530) );
  XOR2_X1 U583 ( .A(KEYINPUT0), .B(G543), .Z(n628) );
  NAND2_X1 U584 ( .A1(G51), .A2(n657), .ZN(n529) );
  NAND2_X1 U585 ( .A1(n530), .A2(n529), .ZN(n531) );
  XOR2_X1 U586 ( .A(KEYINPUT6), .B(n531), .Z(n540) );
  NOR2_X1 U587 ( .A1(n628), .A2(n532), .ZN(n651) );
  NAND2_X1 U588 ( .A1(n651), .A2(G76), .ZN(n533) );
  XNOR2_X1 U589 ( .A(KEYINPUT77), .B(n533), .ZN(n536) );
  NOR2_X1 U590 ( .A1(G543), .A2(G651), .ZN(n650) );
  NAND2_X1 U591 ( .A1(n650), .A2(G89), .ZN(n534) );
  XOR2_X1 U592 ( .A(n534), .B(KEYINPUT4), .Z(n535) );
  NOR2_X1 U593 ( .A1(n536), .A2(n535), .ZN(n537) );
  XOR2_X1 U594 ( .A(KEYINPUT78), .B(n537), .Z(n538) );
  XNOR2_X1 U595 ( .A(KEYINPUT5), .B(n538), .ZN(n539) );
  NAND2_X1 U596 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U597 ( .A(KEYINPUT7), .B(n541), .ZN(G168) );
  AND2_X1 U598 ( .A1(G2104), .A2(G2105), .ZN(n900) );
  NAND2_X1 U599 ( .A1(G113), .A2(n900), .ZN(n542) );
  XOR2_X1 U600 ( .A(KEYINPUT67), .B(n542), .Z(n549) );
  INV_X1 U601 ( .A(KEYINPUT23), .ZN(n544) );
  NAND2_X1 U602 ( .A1(G101), .A2(n904), .ZN(n543) );
  XNOR2_X1 U603 ( .A(n544), .B(n543), .ZN(n547) );
  NAND2_X1 U604 ( .A1(G125), .A2(n901), .ZN(n546) );
  AND2_X1 U605 ( .A1(n547), .A2(n546), .ZN(n548) );
  AND2_X1 U606 ( .A1(n549), .A2(n548), .ZN(n553) );
  XOR2_X1 U607 ( .A(KEYINPUT68), .B(n550), .Z(n551) );
  XNOR2_X1 U608 ( .A(KEYINPUT17), .B(n551), .ZN(n696) );
  NAND2_X1 U609 ( .A1(n696), .A2(G137), .ZN(n552) );
  NAND2_X1 U610 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X2 U611 ( .A(KEYINPUT66), .B(n554), .Z(G160) );
  BUF_X1 U612 ( .A(n696), .Z(n905) );
  NAND2_X1 U613 ( .A1(G138), .A2(n905), .ZN(n559) );
  AND2_X1 U614 ( .A1(G102), .A2(n904), .ZN(n558) );
  NAND2_X1 U615 ( .A1(G114), .A2(n900), .ZN(n556) );
  NAND2_X1 U616 ( .A1(G126), .A2(n901), .ZN(n555) );
  NAND2_X1 U617 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U618 ( .A1(n558), .A2(n557), .ZN(n697) );
  AND2_X1 U619 ( .A1(n559), .A2(n697), .ZN(G164) );
  NAND2_X1 U620 ( .A1(G64), .A2(n653), .ZN(n561) );
  NAND2_X1 U621 ( .A1(G52), .A2(n657), .ZN(n560) );
  NAND2_X1 U622 ( .A1(n561), .A2(n560), .ZN(n567) );
  NAND2_X1 U623 ( .A1(G90), .A2(n650), .ZN(n563) );
  NAND2_X1 U624 ( .A1(G77), .A2(n651), .ZN(n562) );
  NAND2_X1 U625 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U626 ( .A(KEYINPUT71), .B(n564), .ZN(n565) );
  XNOR2_X1 U627 ( .A(KEYINPUT9), .B(n565), .ZN(n566) );
  NOR2_X1 U628 ( .A1(n567), .A2(n566), .ZN(G171) );
  AND2_X1 U629 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U630 ( .A(G132), .ZN(G219) );
  INV_X1 U631 ( .A(G82), .ZN(G220) );
  INV_X1 U632 ( .A(G57), .ZN(G237) );
  XOR2_X1 U633 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U634 ( .A(KEYINPUT10), .B(KEYINPUT73), .Z(n569) );
  NAND2_X1 U635 ( .A1(G7), .A2(G661), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(G223) );
  INV_X1 U637 ( .A(G223), .ZN(n847) );
  NAND2_X1 U638 ( .A1(n847), .A2(G567), .ZN(n570) );
  XOR2_X1 U639 ( .A(KEYINPUT11), .B(n570), .Z(G234) );
  NAND2_X1 U640 ( .A1(G56), .A2(n653), .ZN(n571) );
  XOR2_X1 U641 ( .A(KEYINPUT14), .B(n571), .Z(n577) );
  NAND2_X1 U642 ( .A1(n650), .A2(G81), .ZN(n572) );
  XNOR2_X1 U643 ( .A(n572), .B(KEYINPUT12), .ZN(n574) );
  NAND2_X1 U644 ( .A1(G68), .A2(n651), .ZN(n573) );
  NAND2_X1 U645 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U646 ( .A(KEYINPUT13), .B(n575), .Z(n576) );
  NOR2_X1 U647 ( .A1(n577), .A2(n576), .ZN(n579) );
  NAND2_X1 U648 ( .A1(n657), .A2(G43), .ZN(n578) );
  NAND2_X1 U649 ( .A1(n579), .A2(n578), .ZN(n997) );
  INV_X1 U650 ( .A(G860), .ZN(n603) );
  OR2_X1 U651 ( .A1(n997), .A2(n603), .ZN(G153) );
  INV_X1 U652 ( .A(G171), .ZN(G301) );
  NAND2_X1 U653 ( .A1(G66), .A2(n653), .ZN(n581) );
  NAND2_X1 U654 ( .A1(G92), .A2(n650), .ZN(n580) );
  NAND2_X1 U655 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U656 ( .A(KEYINPUT74), .B(n582), .ZN(n586) );
  NAND2_X1 U657 ( .A1(G54), .A2(n657), .ZN(n584) );
  NAND2_X1 U658 ( .A1(G79), .A2(n651), .ZN(n583) );
  NAND2_X1 U659 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U660 ( .A1(n586), .A2(n585), .ZN(n588) );
  XNOR2_X1 U661 ( .A(KEYINPUT75), .B(KEYINPUT15), .ZN(n587) );
  XNOR2_X1 U662 ( .A(n588), .B(n587), .ZN(n917) );
  INV_X1 U663 ( .A(n917), .ZN(n987) );
  NOR2_X1 U664 ( .A1(G868), .A2(n987), .ZN(n590) );
  INV_X1 U665 ( .A(G868), .ZN(n664) );
  NOR2_X1 U666 ( .A1(n664), .A2(G301), .ZN(n589) );
  NOR2_X1 U667 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U668 ( .A(KEYINPUT76), .B(n591), .ZN(G284) );
  NAND2_X1 U669 ( .A1(G65), .A2(n653), .ZN(n593) );
  NAND2_X1 U670 ( .A1(G91), .A2(n650), .ZN(n592) );
  NAND2_X1 U671 ( .A1(n593), .A2(n592), .ZN(n597) );
  NAND2_X1 U672 ( .A1(G53), .A2(n657), .ZN(n595) );
  NAND2_X1 U673 ( .A1(G78), .A2(n651), .ZN(n594) );
  NAND2_X1 U674 ( .A1(n595), .A2(n594), .ZN(n596) );
  NOR2_X1 U675 ( .A1(n597), .A2(n596), .ZN(n598) );
  XOR2_X1 U676 ( .A(KEYINPUT72), .B(n598), .Z(G299) );
  XNOR2_X1 U677 ( .A(KEYINPUT79), .B(G868), .ZN(n599) );
  NOR2_X1 U678 ( .A1(G286), .A2(n599), .ZN(n601) );
  NOR2_X1 U679 ( .A1(G299), .A2(G868), .ZN(n600) );
  NOR2_X1 U680 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U681 ( .A(KEYINPUT80), .B(n602), .ZN(G297) );
  NAND2_X1 U682 ( .A1(n603), .A2(G559), .ZN(n604) );
  NAND2_X1 U683 ( .A1(n604), .A2(n917), .ZN(n605) );
  XNOR2_X1 U684 ( .A(n605), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U685 ( .A1(G868), .A2(n997), .ZN(n608) );
  NAND2_X1 U686 ( .A1(n917), .A2(G868), .ZN(n606) );
  NOR2_X1 U687 ( .A1(G559), .A2(n606), .ZN(n607) );
  NOR2_X1 U688 ( .A1(n608), .A2(n607), .ZN(n609) );
  XOR2_X1 U689 ( .A(KEYINPUT81), .B(n609), .Z(G282) );
  NAND2_X1 U690 ( .A1(G123), .A2(n901), .ZN(n610) );
  XNOR2_X1 U691 ( .A(n610), .B(KEYINPUT18), .ZN(n611) );
  XNOR2_X1 U692 ( .A(n611), .B(KEYINPUT82), .ZN(n613) );
  NAND2_X1 U693 ( .A1(G111), .A2(n900), .ZN(n612) );
  NAND2_X1 U694 ( .A1(n613), .A2(n612), .ZN(n617) );
  NAND2_X1 U695 ( .A1(G99), .A2(n904), .ZN(n615) );
  NAND2_X1 U696 ( .A1(G135), .A2(n905), .ZN(n614) );
  NAND2_X1 U697 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U698 ( .A1(n617), .A2(n616), .ZN(n948) );
  XNOR2_X1 U699 ( .A(G2096), .B(n948), .ZN(n619) );
  INV_X1 U700 ( .A(G2100), .ZN(n618) );
  NAND2_X1 U701 ( .A1(n619), .A2(n618), .ZN(G156) );
  NAND2_X1 U702 ( .A1(n917), .A2(G559), .ZN(n674) );
  XNOR2_X1 U703 ( .A(n997), .B(n674), .ZN(n620) );
  NOR2_X1 U704 ( .A1(n620), .A2(G860), .ZN(n627) );
  NAND2_X1 U705 ( .A1(G67), .A2(n653), .ZN(n622) );
  NAND2_X1 U706 ( .A1(G93), .A2(n650), .ZN(n621) );
  NAND2_X1 U707 ( .A1(n622), .A2(n621), .ZN(n626) );
  NAND2_X1 U708 ( .A1(G55), .A2(n657), .ZN(n624) );
  NAND2_X1 U709 ( .A1(G80), .A2(n651), .ZN(n623) );
  NAND2_X1 U710 ( .A1(n624), .A2(n623), .ZN(n625) );
  OR2_X1 U711 ( .A1(n626), .A2(n625), .ZN(n666) );
  XOR2_X1 U712 ( .A(n627), .B(n666), .Z(G145) );
  NAND2_X1 U713 ( .A1(n628), .A2(G87), .ZN(n633) );
  NAND2_X1 U714 ( .A1(G49), .A2(n657), .ZN(n630) );
  NAND2_X1 U715 ( .A1(G74), .A2(G651), .ZN(n629) );
  NAND2_X1 U716 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U717 ( .A1(n653), .A2(n631), .ZN(n632) );
  NAND2_X1 U718 ( .A1(n633), .A2(n632), .ZN(n634) );
  XOR2_X1 U719 ( .A(KEYINPUT83), .B(n634), .Z(G288) );
  NAND2_X1 U720 ( .A1(G88), .A2(n650), .ZN(n636) );
  NAND2_X1 U721 ( .A1(G75), .A2(n651), .ZN(n635) );
  NAND2_X1 U722 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U723 ( .A(KEYINPUT87), .B(n637), .ZN(n641) );
  NAND2_X1 U724 ( .A1(G62), .A2(n653), .ZN(n639) );
  NAND2_X1 U725 ( .A1(G50), .A2(n657), .ZN(n638) );
  AND2_X1 U726 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U727 ( .A1(n641), .A2(n640), .ZN(G303) );
  INV_X1 U728 ( .A(G303), .ZN(G166) );
  NAND2_X1 U729 ( .A1(G85), .A2(n650), .ZN(n643) );
  NAND2_X1 U730 ( .A1(G72), .A2(n651), .ZN(n642) );
  NAND2_X1 U731 ( .A1(n643), .A2(n642), .ZN(n648) );
  NAND2_X1 U732 ( .A1(G60), .A2(n653), .ZN(n645) );
  NAND2_X1 U733 ( .A1(G47), .A2(n657), .ZN(n644) );
  NAND2_X1 U734 ( .A1(n645), .A2(n644), .ZN(n646) );
  XOR2_X1 U735 ( .A(KEYINPUT69), .B(n646), .Z(n647) );
  NOR2_X1 U736 ( .A1(n648), .A2(n647), .ZN(n649) );
  XOR2_X1 U737 ( .A(KEYINPUT70), .B(n649), .Z(G290) );
  NAND2_X1 U738 ( .A1(G86), .A2(n650), .ZN(n662) );
  NAND2_X1 U739 ( .A1(G73), .A2(n651), .ZN(n652) );
  XNOR2_X1 U740 ( .A(n652), .B(KEYINPUT2), .ZN(n656) );
  NAND2_X1 U741 ( .A1(G61), .A2(n653), .ZN(n654) );
  XNOR2_X1 U742 ( .A(n654), .B(KEYINPUT84), .ZN(n655) );
  NAND2_X1 U743 ( .A1(n656), .A2(n655), .ZN(n660) );
  NAND2_X1 U744 ( .A1(G48), .A2(n657), .ZN(n658) );
  XNOR2_X1 U745 ( .A(KEYINPUT85), .B(n658), .ZN(n659) );
  NOR2_X1 U746 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U747 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U748 ( .A(n663), .B(KEYINPUT86), .ZN(G305) );
  NAND2_X1 U749 ( .A1(n664), .A2(n666), .ZN(n665) );
  XNOR2_X1 U750 ( .A(n665), .B(KEYINPUT90), .ZN(n678) );
  XNOR2_X1 U751 ( .A(G299), .B(G288), .ZN(n673) );
  XNOR2_X1 U752 ( .A(KEYINPUT19), .B(KEYINPUT88), .ZN(n667) );
  XOR2_X1 U753 ( .A(n667), .B(n666), .Z(n668) );
  XNOR2_X1 U754 ( .A(G166), .B(n668), .ZN(n671) );
  XNOR2_X1 U755 ( .A(G290), .B(G305), .ZN(n669) );
  XNOR2_X1 U756 ( .A(n669), .B(n997), .ZN(n670) );
  XNOR2_X1 U757 ( .A(n671), .B(n670), .ZN(n672) );
  XNOR2_X1 U758 ( .A(n673), .B(n672), .ZN(n918) );
  XNOR2_X1 U759 ( .A(KEYINPUT89), .B(n674), .ZN(n675) );
  XNOR2_X1 U760 ( .A(n918), .B(n675), .ZN(n676) );
  NAND2_X1 U761 ( .A1(G868), .A2(n676), .ZN(n677) );
  NAND2_X1 U762 ( .A1(n678), .A2(n677), .ZN(G295) );
  NAND2_X1 U763 ( .A1(G2078), .A2(G2084), .ZN(n679) );
  XOR2_X1 U764 ( .A(KEYINPUT20), .B(n679), .Z(n680) );
  NAND2_X1 U765 ( .A1(G2090), .A2(n680), .ZN(n681) );
  XNOR2_X1 U766 ( .A(KEYINPUT21), .B(n681), .ZN(n682) );
  NAND2_X1 U767 ( .A1(n682), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U768 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U769 ( .A1(G120), .A2(G69), .ZN(n683) );
  XOR2_X1 U770 ( .A(KEYINPUT91), .B(n683), .Z(n684) );
  NOR2_X1 U771 ( .A1(G237), .A2(n684), .ZN(n685) );
  XNOR2_X1 U772 ( .A(KEYINPUT92), .B(n685), .ZN(n686) );
  NAND2_X1 U773 ( .A1(n686), .A2(G108), .ZN(n851) );
  NAND2_X1 U774 ( .A1(n851), .A2(G567), .ZN(n691) );
  NOR2_X1 U775 ( .A1(G220), .A2(G219), .ZN(n687) );
  XOR2_X1 U776 ( .A(KEYINPUT22), .B(n687), .Z(n688) );
  NOR2_X1 U777 ( .A1(G218), .A2(n688), .ZN(n689) );
  NAND2_X1 U778 ( .A1(G96), .A2(n689), .ZN(n852) );
  NAND2_X1 U779 ( .A1(n852), .A2(G2106), .ZN(n690) );
  NAND2_X1 U780 ( .A1(n691), .A2(n690), .ZN(n853) );
  NAND2_X1 U781 ( .A1(G661), .A2(G483), .ZN(n692) );
  XOR2_X1 U782 ( .A(KEYINPUT93), .B(n692), .Z(n693) );
  NOR2_X1 U783 ( .A1(n853), .A2(n693), .ZN(n850) );
  NAND2_X1 U784 ( .A1(n850), .A2(G36), .ZN(G176) );
  XOR2_X1 U785 ( .A(KEYINPUT101), .B(KEYINPUT27), .Z(n703) );
  NAND2_X1 U786 ( .A1(G40), .A2(G160), .ZN(n797) );
  INV_X1 U787 ( .A(G1384), .ZN(n694) );
  AND2_X1 U788 ( .A1(G138), .A2(n694), .ZN(n695) );
  NAND2_X1 U789 ( .A1(n696), .A2(n695), .ZN(n699) );
  OR2_X1 U790 ( .A1(G1384), .A2(n697), .ZN(n698) );
  NAND2_X1 U791 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U792 ( .A(n700), .B(KEYINPUT64), .ZN(n798) );
  INV_X1 U793 ( .A(n798), .ZN(n701) );
  NAND2_X1 U794 ( .A1(G2072), .A2(n732), .ZN(n702) );
  XNOR2_X1 U795 ( .A(n703), .B(n702), .ZN(n705) );
  INV_X1 U796 ( .A(G1956), .ZN(n1019) );
  NOR2_X1 U797 ( .A1(n732), .A2(n1019), .ZN(n704) );
  NOR2_X1 U798 ( .A1(n705), .A2(n704), .ZN(n725) );
  INV_X1 U799 ( .A(G299), .ZN(n724) );
  NOR2_X1 U800 ( .A1(n725), .A2(n724), .ZN(n706) );
  XOR2_X1 U801 ( .A(n706), .B(KEYINPUT28), .Z(n729) );
  INV_X1 U802 ( .A(n738), .ZN(n709) );
  INV_X1 U803 ( .A(G1996), .ZN(n967) );
  XNOR2_X1 U804 ( .A(KEYINPUT65), .B(KEYINPUT26), .ZN(n707) );
  XNOR2_X1 U805 ( .A(n708), .B(n707), .ZN(n713) );
  NAND2_X1 U806 ( .A1(n753), .A2(G1341), .ZN(n711) );
  OR2_X1 U807 ( .A1(n917), .A2(n714), .ZN(n721) );
  NAND2_X1 U808 ( .A1(n917), .A2(n714), .ZN(n719) );
  AND2_X1 U809 ( .A1(n732), .A2(G2067), .ZN(n715) );
  XOR2_X1 U810 ( .A(n715), .B(KEYINPUT102), .Z(n717) );
  NAND2_X1 U811 ( .A1(n753), .A2(G1348), .ZN(n716) );
  NAND2_X1 U812 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U813 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U814 ( .A1(n721), .A2(n720), .ZN(n723) );
  NAND2_X1 U815 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U816 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U817 ( .A1(n729), .A2(n728), .ZN(n731) );
  INV_X1 U818 ( .A(KEYINPUT29), .ZN(n730) );
  NOR2_X1 U819 ( .A1(n732), .A2(G1961), .ZN(n735) );
  XOR2_X1 U820 ( .A(G2078), .B(KEYINPUT100), .Z(n733) );
  XNOR2_X1 U821 ( .A(KEYINPUT25), .B(n733), .ZN(n969) );
  NOR2_X1 U822 ( .A1(n753), .A2(n969), .ZN(n734) );
  NOR2_X1 U823 ( .A1(n735), .A2(n734), .ZN(n746) );
  OR2_X1 U824 ( .A1(n746), .A2(G301), .ZN(n736) );
  NAND2_X1 U825 ( .A1(n737), .A2(n736), .ZN(n751) );
  INV_X1 U826 ( .A(KEYINPUT99), .ZN(n740) );
  NAND2_X2 U827 ( .A1(G8), .A2(n709), .ZN(n791) );
  NOR2_X1 U828 ( .A1(G1966), .A2(n791), .ZN(n739) );
  XNOR2_X1 U829 ( .A(n740), .B(n739), .ZN(n765) );
  NOR2_X1 U830 ( .A1(G2084), .A2(n753), .ZN(n762) );
  NOR2_X1 U831 ( .A1(n765), .A2(n762), .ZN(n741) );
  NAND2_X1 U832 ( .A1(n741), .A2(G8), .ZN(n743) );
  XNOR2_X1 U833 ( .A(n745), .B(KEYINPUT105), .ZN(n748) );
  NAND2_X1 U834 ( .A1(n746), .A2(G301), .ZN(n747) );
  NAND2_X1 U835 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U836 ( .A(KEYINPUT31), .B(n749), .ZN(n750) );
  NAND2_X1 U837 ( .A1(n751), .A2(n750), .ZN(n764) );
  AND2_X1 U838 ( .A1(G286), .A2(G8), .ZN(n752) );
  NAND2_X1 U839 ( .A1(n764), .A2(n752), .ZN(n760) );
  INV_X1 U840 ( .A(G8), .ZN(n758) );
  NOR2_X1 U841 ( .A1(G1971), .A2(n791), .ZN(n755) );
  NOR2_X1 U842 ( .A1(G2090), .A2(n753), .ZN(n754) );
  NOR2_X1 U843 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U844 ( .A1(n756), .A2(G303), .ZN(n757) );
  OR2_X1 U845 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U846 ( .A(n761), .B(KEYINPUT32), .ZN(n784) );
  NAND2_X1 U847 ( .A1(G8), .A2(n762), .ZN(n763) );
  INV_X1 U848 ( .A(n765), .ZN(n766) );
  NAND2_X1 U849 ( .A1(n767), .A2(n766), .ZN(n783) );
  NAND2_X1 U850 ( .A1(G1976), .A2(G288), .ZN(n995) );
  INV_X1 U851 ( .A(n995), .ZN(n768) );
  OR2_X1 U852 ( .A1(KEYINPUT33), .A2(n527), .ZN(n770) );
  AND2_X1 U853 ( .A1(n783), .A2(n770), .ZN(n769) );
  AND2_X1 U854 ( .A1(n784), .A2(n769), .ZN(n777) );
  INV_X1 U855 ( .A(n770), .ZN(n775) );
  NOR2_X1 U856 ( .A1(G1976), .A2(G288), .ZN(n994) );
  NOR2_X1 U857 ( .A1(G1971), .A2(G303), .ZN(n771) );
  NOR2_X1 U858 ( .A1(n994), .A2(n771), .ZN(n773) );
  INV_X1 U859 ( .A(KEYINPUT33), .ZN(n772) );
  AND2_X1 U860 ( .A1(n773), .A2(n772), .ZN(n774) );
  NOR2_X1 U861 ( .A1(n775), .A2(n774), .ZN(n776) );
  NOR2_X1 U862 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U863 ( .A(n778), .B(KEYINPUT106), .ZN(n781) );
  NAND2_X1 U864 ( .A1(n994), .A2(KEYINPUT33), .ZN(n779) );
  NOR2_X1 U865 ( .A1(n791), .A2(n779), .ZN(n780) );
  NOR2_X1 U866 ( .A1(n781), .A2(n780), .ZN(n782) );
  XOR2_X1 U867 ( .A(G1981), .B(G305), .Z(n990) );
  NAND2_X1 U868 ( .A1(n782), .A2(n990), .ZN(n795) );
  NAND2_X1 U869 ( .A1(n784), .A2(n783), .ZN(n787) );
  NOR2_X1 U870 ( .A1(G2090), .A2(G303), .ZN(n785) );
  NAND2_X1 U871 ( .A1(G8), .A2(n785), .ZN(n786) );
  NAND2_X1 U872 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U873 ( .A1(n788), .A2(n791), .ZN(n793) );
  NOR2_X1 U874 ( .A1(G1981), .A2(G305), .ZN(n789) );
  XOR2_X1 U875 ( .A(n789), .B(KEYINPUT24), .Z(n790) );
  NOR2_X1 U876 ( .A1(n791), .A2(n790), .ZN(n792) );
  NOR2_X1 U877 ( .A1(n793), .A2(n792), .ZN(n794) );
  AND2_X1 U878 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U879 ( .A(n796), .B(KEYINPUT107), .ZN(n830) );
  NOR2_X1 U880 ( .A1(n797), .A2(n798), .ZN(n842) );
  XNOR2_X1 U881 ( .A(KEYINPUT34), .B(KEYINPUT94), .ZN(n802) );
  NAND2_X1 U882 ( .A1(G104), .A2(n904), .ZN(n800) );
  NAND2_X1 U883 ( .A1(G140), .A2(n905), .ZN(n799) );
  NAND2_X1 U884 ( .A1(n800), .A2(n799), .ZN(n801) );
  XNOR2_X1 U885 ( .A(n802), .B(n801), .ZN(n808) );
  NAND2_X1 U886 ( .A1(n900), .A2(G116), .ZN(n803) );
  XOR2_X1 U887 ( .A(KEYINPUT95), .B(n803), .Z(n805) );
  NAND2_X1 U888 ( .A1(n901), .A2(G128), .ZN(n804) );
  NAND2_X1 U889 ( .A1(n805), .A2(n804), .ZN(n806) );
  XOR2_X1 U890 ( .A(KEYINPUT35), .B(n806), .Z(n807) );
  NOR2_X1 U891 ( .A1(n808), .A2(n807), .ZN(n809) );
  XNOR2_X1 U892 ( .A(KEYINPUT36), .B(n809), .ZN(n913) );
  XNOR2_X1 U893 ( .A(KEYINPUT37), .B(G2067), .ZN(n840) );
  NOR2_X1 U894 ( .A1(n913), .A2(n840), .ZN(n943) );
  NAND2_X1 U895 ( .A1(n842), .A2(n943), .ZN(n838) );
  NAND2_X1 U896 ( .A1(G95), .A2(n904), .ZN(n811) );
  NAND2_X1 U897 ( .A1(G131), .A2(n905), .ZN(n810) );
  NAND2_X1 U898 ( .A1(n811), .A2(n810), .ZN(n815) );
  NAND2_X1 U899 ( .A1(G107), .A2(n900), .ZN(n813) );
  NAND2_X1 U900 ( .A1(G119), .A2(n901), .ZN(n812) );
  NAND2_X1 U901 ( .A1(n813), .A2(n812), .ZN(n814) );
  OR2_X1 U902 ( .A1(n815), .A2(n814), .ZN(n884) );
  AND2_X1 U903 ( .A1(n884), .A2(G1991), .ZN(n825) );
  XOR2_X1 U904 ( .A(KEYINPUT96), .B(KEYINPUT38), .Z(n817) );
  NAND2_X1 U905 ( .A1(G105), .A2(n904), .ZN(n816) );
  XNOR2_X1 U906 ( .A(n817), .B(n816), .ZN(n821) );
  NAND2_X1 U907 ( .A1(G129), .A2(n901), .ZN(n819) );
  NAND2_X1 U908 ( .A1(G141), .A2(n905), .ZN(n818) );
  NAND2_X1 U909 ( .A1(n819), .A2(n818), .ZN(n820) );
  NOR2_X1 U910 ( .A1(n821), .A2(n820), .ZN(n823) );
  NAND2_X1 U911 ( .A1(n900), .A2(G117), .ZN(n822) );
  NAND2_X1 U912 ( .A1(n823), .A2(n822), .ZN(n897) );
  AND2_X1 U913 ( .A1(n897), .A2(G1996), .ZN(n824) );
  NOR2_X1 U914 ( .A1(n825), .A2(n824), .ZN(n942) );
  INV_X1 U915 ( .A(n842), .ZN(n826) );
  NOR2_X1 U916 ( .A1(n942), .A2(n826), .ZN(n834) );
  INV_X1 U917 ( .A(n834), .ZN(n827) );
  NAND2_X1 U918 ( .A1(n838), .A2(n827), .ZN(n828) );
  XOR2_X1 U919 ( .A(KEYINPUT97), .B(n828), .Z(n829) );
  XNOR2_X1 U920 ( .A(G1986), .B(G290), .ZN(n989) );
  NAND2_X1 U921 ( .A1(n830), .A2(n525), .ZN(n845) );
  XOR2_X1 U922 ( .A(KEYINPUT109), .B(KEYINPUT39), .Z(n831) );
  XNOR2_X1 U923 ( .A(KEYINPUT108), .B(n831), .ZN(n837) );
  NOR2_X1 U924 ( .A1(G1996), .A2(n897), .ZN(n939) );
  NOR2_X1 U925 ( .A1(G1991), .A2(n884), .ZN(n949) );
  NOR2_X1 U926 ( .A1(G1986), .A2(G290), .ZN(n832) );
  NOR2_X1 U927 ( .A1(n949), .A2(n832), .ZN(n833) );
  NOR2_X1 U928 ( .A1(n834), .A2(n833), .ZN(n835) );
  NOR2_X1 U929 ( .A1(n939), .A2(n835), .ZN(n836) );
  XNOR2_X1 U930 ( .A(n837), .B(n836), .ZN(n839) );
  NAND2_X1 U931 ( .A1(n839), .A2(n838), .ZN(n841) );
  NAND2_X1 U932 ( .A1(n913), .A2(n840), .ZN(n945) );
  NAND2_X1 U933 ( .A1(n841), .A2(n945), .ZN(n843) );
  NAND2_X1 U934 ( .A1(n843), .A2(n842), .ZN(n844) );
  NAND2_X1 U935 ( .A1(n845), .A2(n844), .ZN(n846) );
  XNOR2_X1 U936 ( .A(n846), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U937 ( .A1(G2106), .A2(n847), .ZN(G217) );
  AND2_X1 U938 ( .A1(G15), .A2(G2), .ZN(n848) );
  NAND2_X1 U939 ( .A1(G661), .A2(n848), .ZN(G259) );
  NAND2_X1 U940 ( .A1(G3), .A2(G1), .ZN(n849) );
  NAND2_X1 U941 ( .A1(n850), .A2(n849), .ZN(G188) );
  XNOR2_X1 U942 ( .A(G69), .B(KEYINPUT111), .ZN(G235) );
  INV_X1 U944 ( .A(G120), .ZN(G236) );
  INV_X1 U945 ( .A(G108), .ZN(G238) );
  INV_X1 U946 ( .A(G96), .ZN(G221) );
  NOR2_X1 U947 ( .A1(n852), .A2(n851), .ZN(G325) );
  INV_X1 U948 ( .A(G325), .ZN(G261) );
  INV_X1 U949 ( .A(n853), .ZN(G319) );
  XOR2_X1 U950 ( .A(KEYINPUT41), .B(G1971), .Z(n855) );
  XNOR2_X1 U951 ( .A(G1961), .B(G1956), .ZN(n854) );
  XNOR2_X1 U952 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U953 ( .A(n856), .B(KEYINPUT114), .Z(n858) );
  XNOR2_X1 U954 ( .A(G1996), .B(G1991), .ZN(n857) );
  XNOR2_X1 U955 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U956 ( .A(G1976), .B(G1981), .Z(n860) );
  XNOR2_X1 U957 ( .A(G1986), .B(G1966), .ZN(n859) );
  XNOR2_X1 U958 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U959 ( .A(n862), .B(n861), .Z(n864) );
  XNOR2_X1 U960 ( .A(KEYINPUT113), .B(G2474), .ZN(n863) );
  XNOR2_X1 U961 ( .A(n864), .B(n863), .ZN(G229) );
  XOR2_X1 U962 ( .A(G2096), .B(KEYINPUT43), .Z(n866) );
  XNOR2_X1 U963 ( .A(G2090), .B(G2678), .ZN(n865) );
  XNOR2_X1 U964 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U965 ( .A(n867), .B(KEYINPUT112), .Z(n869) );
  XNOR2_X1 U966 ( .A(G2067), .B(G2072), .ZN(n868) );
  XNOR2_X1 U967 ( .A(n869), .B(n868), .ZN(n873) );
  XOR2_X1 U968 ( .A(KEYINPUT42), .B(G2100), .Z(n871) );
  XNOR2_X1 U969 ( .A(G2078), .B(G2084), .ZN(n870) );
  XNOR2_X1 U970 ( .A(n871), .B(n870), .ZN(n872) );
  XNOR2_X1 U971 ( .A(n873), .B(n872), .ZN(G227) );
  NAND2_X1 U972 ( .A1(G124), .A2(n901), .ZN(n874) );
  XNOR2_X1 U973 ( .A(n874), .B(KEYINPUT44), .ZN(n876) );
  NAND2_X1 U974 ( .A1(n900), .A2(G112), .ZN(n875) );
  NAND2_X1 U975 ( .A1(n876), .A2(n875), .ZN(n880) );
  NAND2_X1 U976 ( .A1(G100), .A2(n904), .ZN(n878) );
  NAND2_X1 U977 ( .A1(G136), .A2(n905), .ZN(n877) );
  NAND2_X1 U978 ( .A1(n878), .A2(n877), .ZN(n879) );
  NOR2_X1 U979 ( .A1(n880), .A2(n879), .ZN(G162) );
  XOR2_X1 U980 ( .A(KEYINPUT118), .B(KEYINPUT115), .Z(n882) );
  XNOR2_X1 U981 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n881) );
  XNOR2_X1 U982 ( .A(n882), .B(n881), .ZN(n883) );
  XOR2_X1 U983 ( .A(n883), .B(n948), .Z(n886) );
  XOR2_X1 U984 ( .A(G164), .B(n884), .Z(n885) );
  XNOR2_X1 U985 ( .A(n886), .B(n885), .ZN(n887) );
  XOR2_X1 U986 ( .A(n887), .B(G162), .Z(n899) );
  NAND2_X1 U987 ( .A1(G103), .A2(n904), .ZN(n889) );
  NAND2_X1 U988 ( .A1(G139), .A2(n905), .ZN(n888) );
  NAND2_X1 U989 ( .A1(n889), .A2(n888), .ZN(n896) );
  NAND2_X1 U990 ( .A1(n900), .A2(G115), .ZN(n890) );
  XNOR2_X1 U991 ( .A(n890), .B(KEYINPUT116), .ZN(n892) );
  NAND2_X1 U992 ( .A1(G127), .A2(n901), .ZN(n891) );
  NAND2_X1 U993 ( .A1(n892), .A2(n891), .ZN(n893) );
  XNOR2_X1 U994 ( .A(KEYINPUT117), .B(n893), .ZN(n894) );
  XNOR2_X1 U995 ( .A(KEYINPUT47), .B(n894), .ZN(n895) );
  NOR2_X1 U996 ( .A1(n896), .A2(n895), .ZN(n954) );
  XOR2_X1 U997 ( .A(n897), .B(n954), .Z(n898) );
  XNOR2_X1 U998 ( .A(n899), .B(n898), .ZN(n915) );
  NAND2_X1 U999 ( .A1(G118), .A2(n900), .ZN(n903) );
  NAND2_X1 U1000 ( .A1(G130), .A2(n901), .ZN(n902) );
  NAND2_X1 U1001 ( .A1(n903), .A2(n902), .ZN(n910) );
  NAND2_X1 U1002 ( .A1(G106), .A2(n904), .ZN(n907) );
  NAND2_X1 U1003 ( .A1(G142), .A2(n905), .ZN(n906) );
  NAND2_X1 U1004 ( .A1(n907), .A2(n906), .ZN(n908) );
  XOR2_X1 U1005 ( .A(n908), .B(KEYINPUT45), .Z(n909) );
  NOR2_X1 U1006 ( .A1(n910), .A2(n909), .ZN(n911) );
  XNOR2_X1 U1007 ( .A(n911), .B(G160), .ZN(n912) );
  XNOR2_X1 U1008 ( .A(n913), .B(n912), .ZN(n914) );
  XNOR2_X1 U1009 ( .A(n915), .B(n914), .ZN(n916) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n916), .ZN(G395) );
  XNOR2_X1 U1011 ( .A(n917), .B(G286), .ZN(n919) );
  XNOR2_X1 U1012 ( .A(n919), .B(n918), .ZN(n920) );
  XNOR2_X1 U1013 ( .A(n920), .B(G171), .ZN(n921) );
  NOR2_X1 U1014 ( .A1(G37), .A2(n921), .ZN(G397) );
  XOR2_X1 U1015 ( .A(G2438), .B(KEYINPUT110), .Z(n923) );
  XNOR2_X1 U1016 ( .A(G2443), .B(G2430), .ZN(n922) );
  XNOR2_X1 U1017 ( .A(n923), .B(n922), .ZN(n924) );
  XOR2_X1 U1018 ( .A(n924), .B(G2435), .Z(n926) );
  XNOR2_X1 U1019 ( .A(G1341), .B(G1348), .ZN(n925) );
  XNOR2_X1 U1020 ( .A(n926), .B(n925), .ZN(n930) );
  XOR2_X1 U1021 ( .A(G2451), .B(G2427), .Z(n928) );
  XNOR2_X1 U1022 ( .A(G2454), .B(G2446), .ZN(n927) );
  XNOR2_X1 U1023 ( .A(n928), .B(n927), .ZN(n929) );
  XOR2_X1 U1024 ( .A(n930), .B(n929), .Z(n931) );
  NAND2_X1 U1025 ( .A1(G14), .A2(n931), .ZN(n937) );
  NAND2_X1 U1026 ( .A1(G319), .A2(n937), .ZN(n934) );
  NOR2_X1 U1027 ( .A1(G229), .A2(G227), .ZN(n932) );
  XNOR2_X1 U1028 ( .A(KEYINPUT49), .B(n932), .ZN(n933) );
  NOR2_X1 U1029 ( .A1(n934), .A2(n933), .ZN(n936) );
  NOR2_X1 U1030 ( .A1(G395), .A2(G397), .ZN(n935) );
  NAND2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(G225) );
  INV_X1 U1032 ( .A(G225), .ZN(G308) );
  INV_X1 U1033 ( .A(n937), .ZN(G401) );
  XOR2_X1 U1034 ( .A(G2090), .B(G162), .Z(n938) );
  NOR2_X1 U1035 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1036 ( .A(KEYINPUT51), .B(n940), .Z(n941) );
  NAND2_X1 U1037 ( .A1(n942), .A2(n941), .ZN(n947) );
  INV_X1 U1038 ( .A(n943), .ZN(n944) );
  NAND2_X1 U1039 ( .A1(n945), .A2(n944), .ZN(n946) );
  NOR2_X1 U1040 ( .A1(n947), .A2(n946), .ZN(n961) );
  XOR2_X1 U1041 ( .A(G160), .B(G2084), .Z(n952) );
  NOR2_X1 U1042 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1043 ( .A(KEYINPUT119), .B(n950), .ZN(n951) );
  NOR2_X1 U1044 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1045 ( .A(KEYINPUT120), .B(n953), .Z(n959) );
  XOR2_X1 U1046 ( .A(G2072), .B(n954), .Z(n956) );
  XOR2_X1 U1047 ( .A(G164), .B(G2078), .Z(n955) );
  NOR2_X1 U1048 ( .A1(n956), .A2(n955), .ZN(n957) );
  XOR2_X1 U1049 ( .A(KEYINPUT50), .B(n957), .Z(n958) );
  NOR2_X1 U1050 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1051 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1052 ( .A(KEYINPUT52), .B(n962), .ZN(n963) );
  NAND2_X1 U1053 ( .A1(n963), .A2(G29), .ZN(n1043) );
  XNOR2_X1 U1054 ( .A(G2084), .B(G34), .ZN(n964) );
  XNOR2_X1 U1055 ( .A(n964), .B(KEYINPUT54), .ZN(n982) );
  XNOR2_X1 U1056 ( .A(G2090), .B(G35), .ZN(n979) );
  XNOR2_X1 U1057 ( .A(G2067), .B(G26), .ZN(n966) );
  XNOR2_X1 U1058 ( .A(G33), .B(G2072), .ZN(n965) );
  NOR2_X1 U1059 ( .A1(n966), .A2(n965), .ZN(n974) );
  XNOR2_X1 U1060 ( .A(G32), .B(n967), .ZN(n968) );
  NAND2_X1 U1061 ( .A1(n968), .A2(G28), .ZN(n972) );
  XOR2_X1 U1062 ( .A(G27), .B(n969), .Z(n970) );
  XNOR2_X1 U1063 ( .A(KEYINPUT121), .B(n970), .ZN(n971) );
  NOR2_X1 U1064 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1065 ( .A1(n974), .A2(n973), .ZN(n976) );
  XNOR2_X1 U1066 ( .A(G25), .B(G1991), .ZN(n975) );
  NOR2_X1 U1067 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1068 ( .A(KEYINPUT53), .B(n977), .ZN(n978) );
  NOR2_X1 U1069 ( .A1(n979), .A2(n978), .ZN(n980) );
  XOR2_X1 U1070 ( .A(KEYINPUT122), .B(n980), .Z(n981) );
  NOR2_X1 U1071 ( .A1(n982), .A2(n981), .ZN(n983) );
  XOR2_X1 U1072 ( .A(KEYINPUT123), .B(n983), .Z(n984) );
  NOR2_X1 U1073 ( .A1(G29), .A2(n984), .ZN(n985) );
  XNOR2_X1 U1074 ( .A(KEYINPUT55), .B(n985), .ZN(n986) );
  NAND2_X1 U1075 ( .A1(n986), .A2(G11), .ZN(n1041) );
  XNOR2_X1 U1076 ( .A(G16), .B(KEYINPUT56), .ZN(n1012) );
  XNOR2_X1 U1077 ( .A(G1348), .B(n987), .ZN(n988) );
  NOR2_X1 U1078 ( .A1(n989), .A2(n988), .ZN(n1010) );
  XNOR2_X1 U1079 ( .A(G1966), .B(G168), .ZN(n991) );
  NAND2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1081 ( .A(n992), .B(KEYINPUT124), .ZN(n993) );
  XNOR2_X1 U1082 ( .A(KEYINPUT57), .B(n993), .ZN(n1005) );
  INV_X1 U1083 ( .A(n994), .ZN(n996) );
  NAND2_X1 U1084 ( .A1(n996), .A2(n995), .ZN(n1003) );
  XNOR2_X1 U1085 ( .A(G171), .B(G1961), .ZN(n1001) );
  XNOR2_X1 U1086 ( .A(n997), .B(G1341), .ZN(n999) );
  XNOR2_X1 U1087 ( .A(G299), .B(G1956), .ZN(n998) );
  NOR2_X1 U1088 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1089 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NOR2_X1 U1090 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1091 ( .A1(n1005), .A2(n1004), .ZN(n1008) );
  XOR2_X1 U1092 ( .A(G1971), .B(G303), .Z(n1006) );
  XNOR2_X1 U1093 ( .A(KEYINPUT125), .B(n1006), .ZN(n1007) );
  NOR2_X1 U1094 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1095 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1096 ( .A1(n1012), .A2(n1011), .ZN(n1039) );
  INV_X1 U1097 ( .A(G16), .ZN(n1037) );
  XNOR2_X1 U1098 ( .A(G1986), .B(G24), .ZN(n1017) );
  XNOR2_X1 U1099 ( .A(G1971), .B(G22), .ZN(n1014) );
  XNOR2_X1 U1100 ( .A(G23), .B(G1976), .ZN(n1013) );
  NOR2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1102 ( .A(KEYINPUT127), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1104 ( .A(KEYINPUT58), .B(n1018), .Z(n1034) );
  XOR2_X1 U1105 ( .A(G1961), .B(G5), .Z(n1029) );
  XNOR2_X1 U1106 ( .A(G20), .B(n1019), .ZN(n1023) );
  XNOR2_X1 U1107 ( .A(G1341), .B(G19), .ZN(n1021) );
  XNOR2_X1 U1108 ( .A(G1981), .B(G6), .ZN(n1020) );
  NOR2_X1 U1109 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1110 ( .A1(n1023), .A2(n1022), .ZN(n1026) );
  XOR2_X1 U1111 ( .A(KEYINPUT59), .B(G1348), .Z(n1024) );
  XNOR2_X1 U1112 ( .A(G4), .B(n1024), .ZN(n1025) );
  NOR2_X1 U1113 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1114 ( .A(KEYINPUT60), .B(n1027), .ZN(n1028) );
  NAND2_X1 U1115 ( .A1(n1029), .A2(n1028), .ZN(n1031) );
  XNOR2_X1 U1116 ( .A(G21), .B(G1966), .ZN(n1030) );
  NOR2_X1 U1117 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XOR2_X1 U1118 ( .A(KEYINPUT126), .B(n1032), .Z(n1033) );
  NOR2_X1 U1119 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XNOR2_X1 U1120 ( .A(KEYINPUT61), .B(n1035), .ZN(n1036) );
  NAND2_X1 U1121 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  NAND2_X1 U1122 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  NOR2_X1 U1123 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  NAND2_X1 U1124 ( .A1(n1043), .A2(n1042), .ZN(n1044) );
  XOR2_X1 U1125 ( .A(KEYINPUT62), .B(n1044), .Z(G311) );
  INV_X1 U1126 ( .A(G311), .ZN(G150) );
endmodule

