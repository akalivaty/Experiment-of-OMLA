//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 1 0 1 1 1 0 0 0 1 0 1 1 1 1 1 1 0 0 0 0 1 1 1 1 1 0 1 0 1 1 1 1 1 0 1 0 1 1 1 1 0 1 0 1 0 1 0 0 1 0 0 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:01 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n449, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n567,
    new_n568, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n631, new_n632, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1213;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  XOR2_X1   g013(.A(KEYINPUT66), .B(G96), .Z(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g020(.A(KEYINPUT67), .B(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT68), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G219), .A4(G221), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  AND2_X1   g035(.A1(new_n460), .A2(G137), .ZN(new_n461));
  AND2_X1   g036(.A1(G101), .A2(G2104), .ZN(new_n462));
  OAI211_X1 g037(.A(KEYINPUT70), .B(new_n459), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT70), .ZN(new_n464));
  AOI22_X1  g039(.A1(new_n460), .A2(G137), .B1(G101), .B2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n464), .B1(new_n465), .B2(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n460), .A2(G125), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT69), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n468), .A2(new_n469), .B1(G113), .B2(G2104), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n460), .A2(KEYINPUT69), .A3(G125), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n459), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n467), .A2(new_n472), .ZN(G160));
  OR2_X1    g048(.A1(G100), .A2(G2105), .ZN(new_n474));
  OAI211_X1 g049(.A(new_n474), .B(G2104), .C1(G112), .C2(new_n459), .ZN(new_n475));
  XOR2_X1   g050(.A(new_n475), .B(KEYINPUT71), .Z(new_n476));
  INV_X1    g051(.A(KEYINPUT3), .ZN(new_n477));
  INV_X1    g052(.A(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n459), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g056(.A(G2105), .B1(new_n479), .B2(new_n480), .ZN(new_n482));
  AOI22_X1  g057(.A1(G124), .A2(new_n481), .B1(new_n482), .B2(G136), .ZN(new_n483));
  AND2_X1   g058(.A1(new_n476), .A2(new_n483), .ZN(G162));
  OAI21_X1  g059(.A(G2104), .B1(new_n459), .B2(G114), .ZN(new_n485));
  NOR2_X1   g060(.A1(G102), .A2(G2105), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT72), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n481), .A2(new_n488), .A3(G126), .ZN(new_n489));
  INV_X1    g064(.A(new_n480), .ZN(new_n490));
  NOR2_X1   g065(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n491));
  OAI211_X1 g066(.A(G126), .B(G2105), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT72), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n487), .B1(new_n489), .B2(new_n493), .ZN(new_n494));
  XOR2_X1   g069(.A(KEYINPUT73), .B(KEYINPUT4), .Z(new_n495));
  NAND3_X1  g070(.A1(new_n482), .A2(new_n495), .A3(G138), .ZN(new_n496));
  OAI211_X1 g071(.A(G138), .B(new_n459), .C1(new_n490), .C2(new_n491), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT73), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n494), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  INV_X1    g078(.A(KEYINPUT74), .ZN(new_n504));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT74), .A2(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT6), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT75), .ZN(new_n513));
  NAND4_X1  g088(.A1(new_n512), .A2(new_n513), .A3(G50), .A4(G543), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT6), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n515), .B1(new_n506), .B2(new_n507), .ZN(new_n516));
  OAI211_X1 g091(.A(G50), .B(G543), .C1(new_n516), .C2(new_n510), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(KEYINPUT75), .ZN(new_n518));
  NAND2_X1  g093(.A1(G75), .A2(G543), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT76), .ZN(new_n520));
  INV_X1    g095(.A(G62), .ZN(new_n521));
  OR2_X1    g096(.A1(KEYINPUT5), .A2(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(KEYINPUT5), .A2(G543), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n508), .B1(new_n520), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n522), .A2(new_n523), .ZN(new_n526));
  OAI211_X1 g101(.A(G88), .B(new_n526), .C1(new_n516), .C2(new_n510), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n514), .A2(new_n518), .A3(new_n525), .A4(new_n527), .ZN(G303));
  INV_X1    g103(.A(G303), .ZN(G166));
  AND2_X1   g104(.A1(new_n522), .A2(new_n523), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n530), .B1(new_n509), .B2(new_n511), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G89), .ZN(new_n532));
  INV_X1    g107(.A(G543), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n533), .B1(new_n509), .B2(new_n511), .ZN(new_n534));
  XOR2_X1   g109(.A(KEYINPUT77), .B(G51), .Z(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n537), .A2(KEYINPUT7), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(KEYINPUT7), .ZN(new_n539));
  AND2_X1   g114(.A1(G63), .A2(G651), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n538), .A2(new_n539), .B1(new_n526), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n532), .A2(new_n536), .A3(new_n541), .ZN(G286));
  INV_X1    g117(.A(G286), .ZN(G168));
  NAND2_X1  g118(.A1(new_n531), .A2(G90), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n534), .A2(G52), .ZN(new_n545));
  NAND2_X1  g120(.A1(G77), .A2(G543), .ZN(new_n546));
  INV_X1    g121(.A(G64), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n530), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(new_n508), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n544), .A2(new_n545), .A3(new_n549), .ZN(G301));
  INV_X1    g125(.A(G301), .ZN(G171));
  NAND2_X1  g126(.A1(G68), .A2(G543), .ZN(new_n552));
  INV_X1    g127(.A(G56), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n530), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(new_n508), .ZN(new_n555));
  OAI211_X1 g130(.A(G43), .B(G543), .C1(new_n516), .C2(new_n510), .ZN(new_n556));
  OAI211_X1 g131(.A(G81), .B(new_n526), .C1(new_n516), .C2(new_n510), .ZN(new_n557));
  AND3_X1   g132(.A1(new_n556), .A2(new_n557), .A3(KEYINPUT78), .ZN(new_n558));
  AOI21_X1  g133(.A(KEYINPUT78), .B1(new_n556), .B2(new_n557), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n555), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT79), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OAI211_X1 g137(.A(KEYINPUT79), .B(new_n555), .C1(new_n558), .C2(new_n559), .ZN(new_n563));
  AND2_X1   g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  NAND4_X1  g140(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND4_X1  g143(.A1(G319), .A2(G483), .A3(G661), .A4(new_n568), .ZN(G188));
  INV_X1    g144(.A(KEYINPUT9), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n534), .A2(new_n570), .A3(G53), .ZN(new_n571));
  OAI211_X1 g146(.A(G53), .B(G543), .C1(new_n516), .C2(new_n510), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(KEYINPUT9), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n571), .A2(new_n573), .B1(G91), .B2(new_n531), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT81), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT80), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n522), .A2(new_n576), .A3(new_n523), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n576), .B1(new_n522), .B2(new_n523), .ZN(new_n579));
  OAI21_X1  g154(.A(G65), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(G78), .A2(G543), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n575), .B1(new_n582), .B2(G651), .ZN(new_n583));
  INV_X1    g158(.A(G65), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n526), .A2(KEYINPUT80), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n584), .B1(new_n585), .B2(new_n577), .ZN(new_n586));
  INV_X1    g161(.A(new_n581), .ZN(new_n587));
  OAI211_X1 g162(.A(new_n575), .B(G651), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n574), .B1(new_n583), .B2(new_n589), .ZN(G299));
  NAND2_X1  g165(.A1(new_n534), .A2(G49), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n531), .A2(G87), .ZN(new_n592));
  OAI21_X1  g167(.A(G651), .B1(new_n526), .B2(G74), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(G288));
  INV_X1    g169(.A(G61), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n595), .B1(new_n522), .B2(new_n523), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(KEYINPUT82), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(G73), .A2(G543), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(new_n596), .B2(KEYINPUT82), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n508), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n534), .A2(G48), .ZN(new_n602));
  NAND4_X1  g177(.A1(new_n512), .A2(KEYINPUT83), .A3(G86), .A4(new_n526), .ZN(new_n603));
  OAI211_X1 g178(.A(G86), .B(new_n526), .C1(new_n516), .C2(new_n510), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT83), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g181(.A1(new_n601), .A2(new_n602), .A3(new_n603), .A4(new_n606), .ZN(G305));
  NAND2_X1  g182(.A1(G72), .A2(G543), .ZN(new_n608));
  INV_X1    g183(.A(G60), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n530), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(new_n508), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT84), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n531), .A2(G85), .B1(new_n534), .B2(G47), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(G290));
  NAND2_X1  g189(.A1(G301), .A2(G868), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n531), .A2(G92), .ZN(new_n616));
  XNOR2_X1  g191(.A(KEYINPUT85), .B(KEYINPUT10), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT86), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n534), .A2(G54), .ZN(new_n621));
  INV_X1    g196(.A(G66), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n622), .B1(new_n585), .B2(new_n577), .ZN(new_n623));
  AND2_X1   g198(.A1(G79), .A2(G543), .ZN(new_n624));
  OAI21_X1  g199(.A(G651), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n618), .A2(new_n531), .A3(G92), .ZN(new_n626));
  NAND4_X1  g201(.A1(new_n620), .A2(new_n621), .A3(new_n625), .A4(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n615), .B1(new_n628), .B2(G868), .ZN(G284));
  OAI21_X1  g204(.A(new_n615), .B1(new_n628), .B2(G868), .ZN(G321));
  NAND2_X1  g205(.A1(G286), .A2(G868), .ZN(new_n631));
  INV_X1    g206(.A(G299), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n631), .B1(new_n632), .B2(G868), .ZN(G297));
  OAI21_X1  g208(.A(new_n631), .B1(new_n632), .B2(G868), .ZN(G280));
  INV_X1    g209(.A(G559), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n628), .B1(new_n635), .B2(G860), .ZN(G148));
  INV_X1    g211(.A(G868), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n564), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n627), .A2(G559), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(G868), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT11), .Z(G282));
  INV_X1    g217(.A(new_n641), .ZN(G323));
  NAND2_X1  g218(.A1(new_n482), .A2(G2104), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT12), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT13), .ZN(new_n646));
  INV_X1    g221(.A(G2100), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n482), .A2(G135), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n481), .A2(G123), .ZN(new_n651));
  NOR2_X1   g226(.A1(G99), .A2(G2105), .ZN(new_n652));
  OAI21_X1  g227(.A(G2104), .B1(new_n459), .B2(G111), .ZN(new_n653));
  OAI211_X1 g228(.A(new_n650), .B(new_n651), .C1(new_n652), .C2(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(G2096), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n648), .A2(new_n649), .A3(new_n656), .ZN(G156));
  XOR2_X1   g232(.A(G2451), .B(G2454), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT16), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1341), .B(G1348), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2443), .B(G2446), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2427), .B(G2438), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G2430), .ZN(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT15), .B(G2435), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n665), .A2(new_n666), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n667), .A2(new_n668), .A3(KEYINPUT14), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n663), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n663), .A2(new_n670), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n671), .A2(new_n672), .A3(G14), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT87), .ZN(G401));
  XOR2_X1   g249(.A(G2072), .B(G2078), .Z(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT17), .Z(new_n676));
  XOR2_X1   g251(.A(G2084), .B(G2090), .Z(new_n677));
  XNOR2_X1  g252(.A(G2067), .B(G2678), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n676), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n677), .A2(new_n678), .ZN(new_n680));
  INV_X1    g255(.A(new_n677), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(new_n675), .ZN(new_n682));
  OAI211_X1 g257(.A(new_n679), .B(new_n680), .C1(new_n678), .C2(new_n682), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n680), .A2(new_n675), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT18), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(new_n655), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n687), .A2(G2100), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(G2100), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(G227));
  XOR2_X1   g265(.A(G1971), .B(G1976), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT19), .ZN(new_n692));
  XOR2_X1   g267(.A(G1956), .B(G2474), .Z(new_n693));
  XOR2_X1   g268(.A(G1961), .B(G1966), .Z(new_n694));
  NOR2_X1   g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  AND2_X1   g271(.A1(new_n693), .A2(new_n694), .ZN(new_n697));
  NOR3_X1   g272(.A1(new_n692), .A2(new_n697), .A3(new_n695), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n692), .A2(new_n697), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT88), .B(KEYINPUT20), .ZN(new_n700));
  AOI211_X1 g275(.A(new_n696), .B(new_n698), .C1(new_n699), .C2(new_n700), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(new_n699), .B2(new_n700), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n703));
  INV_X1    g278(.A(G1981), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n702), .B(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(G1991), .B(G1996), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT89), .B(G1986), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(G229));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G26), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT28), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n482), .A2(G140), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT96), .ZN(new_n718));
  OAI21_X1  g293(.A(G2104), .B1(new_n459), .B2(G116), .ZN(new_n719));
  INV_X1    g294(.A(G104), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(new_n459), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT97), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n481), .A2(G128), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n718), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT98), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n716), .B1(new_n726), .B2(new_n714), .ZN(new_n727));
  INV_X1    g302(.A(G2067), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(G16), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G21), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G168), .B2(new_n730), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n732), .A2(G1966), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT104), .Z(new_n734));
  NAND2_X1  g309(.A1(new_n729), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(G171), .A2(new_n730), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G5), .B2(new_n730), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT24), .ZN(new_n739));
  INV_X1    g314(.A(G34), .ZN(new_n740));
  AOI21_X1  g315(.A(G29), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(new_n739), .B2(new_n740), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G160), .B2(new_n714), .ZN(new_n743));
  AOI22_X1  g318(.A1(new_n738), .A2(G1961), .B1(G2084), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n730), .A2(G4), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n628), .B2(new_n730), .ZN(new_n746));
  INV_X1    g321(.A(G1348), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  OAI211_X1 g323(.A(new_n744), .B(new_n748), .C1(G2084), .C2(new_n743), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n735), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g325(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT26), .Z(new_n752));
  NAND2_X1  g327(.A1(new_n482), .A2(G141), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n459), .A2(G105), .A3(G2104), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT99), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n481), .A2(G129), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n754), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT100), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n760), .A2(G29), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT101), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G29), .B2(G32), .ZN(new_n763));
  XOR2_X1   g338(.A(KEYINPUT27), .B(G1996), .Z(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  XOR2_X1   g340(.A(KEYINPUT92), .B(G16), .Z(new_n766));
  NAND2_X1  g341(.A1(new_n766), .A2(G20), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT23), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n632), .B2(new_n730), .ZN(new_n769));
  INV_X1    g344(.A(G1956), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n714), .A2(G27), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G164), .B2(new_n714), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT105), .B(G2078), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n732), .A2(G1966), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n775), .B(new_n776), .C1(new_n738), .C2(G1961), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n714), .A2(G35), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G162), .B2(new_n714), .ZN(new_n779));
  XOR2_X1   g354(.A(KEYINPUT29), .B(G2090), .Z(new_n780));
  XOR2_X1   g355(.A(new_n779), .B(new_n780), .Z(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT102), .B(KEYINPUT31), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G11), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT103), .B(G28), .ZN(new_n784));
  AOI21_X1  g359(.A(G29), .B1(new_n784), .B2(KEYINPUT30), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(KEYINPUT30), .B2(new_n784), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n783), .B(new_n786), .C1(new_n654), .C2(new_n714), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n714), .A2(G33), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT25), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n460), .A2(G127), .ZN(new_n791));
  NAND2_X1  g366(.A1(G115), .A2(G2104), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n459), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  AOI211_X1 g368(.A(new_n790), .B(new_n793), .C1(G139), .C2(new_n482), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n788), .B1(new_n794), .B2(new_n714), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n787), .B1(new_n795), .B2(G2072), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G2072), .B2(new_n795), .ZN(new_n797));
  NOR3_X1   g372(.A1(new_n777), .A2(new_n781), .A3(new_n797), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n765), .A2(new_n771), .A3(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(new_n766), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n800), .A2(G19), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(new_n564), .B2(new_n800), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G1341), .ZN(new_n803));
  NOR3_X1   g378(.A1(new_n750), .A2(new_n799), .A3(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n766), .A2(G22), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT94), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G166), .B2(new_n766), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT95), .Z(new_n809));
  OR2_X1    g384(.A1(new_n809), .A2(G1971), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(G1971), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n730), .A2(G6), .ZN(new_n812));
  INV_X1    g387(.A(G305), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n812), .B1(new_n813), .B2(new_n730), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT32), .B(G1981), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n730), .A2(G23), .ZN(new_n817));
  INV_X1    g392(.A(G288), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(new_n818), .B2(new_n730), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT33), .B(G1976), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n814), .A2(new_n815), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n810), .A2(new_n811), .A3(new_n816), .A4(new_n823), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n824), .A2(KEYINPUT34), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(KEYINPUT34), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n714), .A2(G25), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n482), .A2(G131), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT90), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n481), .A2(G119), .ZN(new_n830));
  NOR2_X1   g405(.A1(G95), .A2(G2105), .ZN(new_n831));
  OAI21_X1  g406(.A(G2104), .B1(new_n459), .B2(G107), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n829), .B(new_n830), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT91), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n827), .B1(new_n835), .B2(new_n714), .ZN(new_n836));
  XOR2_X1   g411(.A(KEYINPUT35), .B(G1991), .Z(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n836), .B(new_n838), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n800), .A2(G24), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(G290), .B2(new_n766), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT93), .ZN(new_n842));
  INV_X1    g417(.A(G1986), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n842), .A2(new_n843), .ZN(new_n845));
  NOR3_X1   g420(.A1(new_n839), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n825), .A2(new_n826), .A3(new_n846), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n847), .A2(KEYINPUT36), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(KEYINPUT36), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n805), .B1(new_n849), .B2(new_n850), .ZN(G311));
  INV_X1    g426(.A(new_n850), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n804), .B1(new_n852), .B2(new_n848), .ZN(G150));
  NAND2_X1  g428(.A1(new_n628), .A2(G559), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT38), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT106), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n531), .A2(G93), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n534), .A2(G55), .ZN(new_n858));
  NAND2_X1  g433(.A1(G80), .A2(G543), .ZN(new_n859));
  INV_X1    g434(.A(G67), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n859), .B1(new_n530), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(new_n508), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n857), .A2(new_n858), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n562), .A2(new_n563), .A3(new_n863), .ZN(new_n864));
  NAND4_X1  g439(.A1(new_n560), .A2(new_n857), .A3(new_n858), .A4(new_n862), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n856), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AND3_X1   g441(.A1(new_n864), .A2(new_n856), .A3(new_n865), .ZN(new_n867));
  OR3_X1    g442(.A1(new_n855), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT39), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n855), .B1(new_n867), .B2(new_n866), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(G860), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n869), .B1(new_n868), .B2(new_n870), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT107), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n863), .A2(G860), .ZN(new_n877));
  XOR2_X1   g452(.A(KEYINPUT108), .B(KEYINPUT37), .Z(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n876), .A2(new_n879), .ZN(G145));
  INV_X1    g455(.A(KEYINPUT109), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n501), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n496), .A2(new_n500), .A3(KEYINPUT109), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n882), .A2(new_n494), .A3(new_n883), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n725), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n725), .A2(new_n884), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(new_n835), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n885), .A2(new_n834), .A3(new_n886), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n760), .A2(new_n794), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n891), .B1(new_n759), .B2(new_n794), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n482), .A2(G142), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n481), .A2(G130), .ZN(new_n894));
  NOR2_X1   g469(.A1(G106), .A2(G2105), .ZN(new_n895));
  OAI21_X1  g470(.A(G2104), .B1(new_n459), .B2(G118), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n893), .B(new_n894), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  XOR2_X1   g472(.A(new_n645), .B(new_n897), .Z(new_n898));
  XNOR2_X1  g473(.A(new_n892), .B(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n890), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(G162), .B(new_n654), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(G160), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n888), .A2(new_n899), .A3(new_n889), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n901), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(G37), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n903), .B1(new_n901), .B2(new_n904), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT40), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n909), .B(new_n910), .ZN(G395));
  NOR3_X1   g486(.A1(new_n867), .A2(new_n866), .A3(new_n639), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(G299), .A2(new_n628), .ZN(new_n914));
  OAI21_X1  g489(.A(G651), .B1(new_n586), .B2(new_n587), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(KEYINPUT81), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(new_n588), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n917), .A2(new_n627), .A3(new_n574), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n914), .A2(KEYINPUT41), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(KEYINPUT41), .B1(new_n914), .B2(new_n918), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n639), .B1(new_n867), .B2(new_n866), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n913), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n913), .A2(new_n923), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n914), .A2(new_n918), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT110), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n914), .A2(KEYINPUT110), .A3(new_n918), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n924), .B1(new_n925), .B2(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(G290), .B(new_n818), .ZN(new_n932));
  XNOR2_X1  g507(.A(G166), .B(G305), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n932), .A2(new_n933), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  XOR2_X1   g511(.A(new_n936), .B(KEYINPUT42), .Z(new_n937));
  AND2_X1   g512(.A1(new_n931), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n931), .A2(new_n937), .ZN(new_n939));
  OAI21_X1  g514(.A(G868), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n863), .A2(new_n637), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(G295));
  NAND2_X1  g517(.A1(new_n940), .A2(new_n941), .ZN(G331));
  NAND2_X1  g518(.A1(G301), .A2(KEYINPUT111), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT111), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n544), .A2(new_n545), .A3(new_n945), .A4(new_n549), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n944), .A2(G168), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(G286), .A2(G301), .A3(KEYINPUT111), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n950), .B1(new_n867), .B2(new_n866), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n864), .A2(new_n865), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT106), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n864), .A2(new_n856), .A3(new_n865), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n953), .A2(new_n954), .A3(new_n949), .ZN(new_n955));
  AND3_X1   g530(.A1(new_n951), .A2(new_n955), .A3(new_n930), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n921), .B1(new_n951), .B2(new_n955), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n936), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NOR3_X1   g533(.A1(new_n867), .A2(new_n866), .A3(new_n950), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n949), .B1(new_n953), .B2(new_n954), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n922), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n936), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n951), .A2(new_n955), .A3(new_n926), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n961), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n958), .A2(new_n964), .A3(new_n906), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT112), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT112), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n958), .A2(new_n964), .A3(new_n967), .A4(new_n906), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n966), .A2(KEYINPUT43), .A3(new_n968), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n951), .A2(new_n955), .A3(new_n926), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n936), .B1(new_n970), .B2(new_n957), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT43), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n971), .A2(new_n964), .A3(new_n972), .A4(new_n906), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n973), .A2(KEYINPUT44), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n969), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT44), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n964), .A2(new_n906), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n972), .B1(new_n977), .B2(new_n971), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n976), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n975), .A2(new_n980), .ZN(G397));
  INV_X1    g556(.A(G1384), .ZN(new_n982));
  AOI21_X1  g557(.A(KEYINPUT45), .B1(new_n884), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(G113), .A2(G2104), .ZN(new_n985));
  INV_X1    g560(.A(G125), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n986), .B1(new_n479), .B2(new_n480), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n985), .B1(new_n987), .B2(KEYINPUT69), .ZN(new_n988));
  INV_X1    g563(.A(new_n471), .ZN(new_n989));
  OAI21_X1  g564(.A(G2105), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n990), .A2(new_n463), .A3(G40), .A4(new_n466), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n984), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G1996), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n992), .A2(KEYINPUT46), .A3(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT46), .ZN(new_n995));
  INV_X1    g570(.A(new_n992), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n995), .B1(new_n996), .B2(G1996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n726), .A2(new_n728), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n725), .A2(G2067), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n998), .A2(new_n759), .A3(new_n999), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n994), .B(new_n997), .C1(new_n1000), .C2(new_n996), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT47), .ZN(new_n1002));
  OR2_X1    g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1003), .A2(KEYINPUT127), .A3(new_n1004), .ZN(new_n1005));
  NOR3_X1   g580(.A1(new_n996), .A2(G1986), .A3(G290), .ZN(new_n1006));
  XOR2_X1   g581(.A(new_n1006), .B(KEYINPUT48), .Z(new_n1007));
  NAND2_X1  g582(.A1(new_n760), .A2(new_n993), .ZN(new_n1008));
  OAI21_X1  g583(.A(G1996), .B1(new_n754), .B2(new_n758), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n998), .A2(new_n999), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n834), .B(new_n838), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n992), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n835), .A2(new_n837), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n998), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1014));
  AOI22_X1  g589(.A1(new_n1007), .A2(new_n1012), .B1(new_n992), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1005), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT127), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT62), .ZN(new_n1019));
  XOR2_X1   g594(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n1020));
  NAND3_X1  g595(.A1(new_n884), .A2(new_n982), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n991), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G2084), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n502), .A2(new_n982), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1025), .A2(KEYINPUT114), .A3(KEYINPUT50), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT114), .ZN(new_n1027));
  AOI21_X1  g602(.A(G1384), .B1(new_n494), .B2(new_n501), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT50), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1027), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1026), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1023), .A2(new_n1024), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G1966), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT45), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1034), .A2(G1384), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n502), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1022), .A2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1033), .B1(new_n1037), .B2(new_n983), .ZN(new_n1038));
  XOR2_X1   g613(.A(KEYINPUT118), .B(G8), .Z(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(G286), .A2(new_n1040), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n1032), .A2(new_n1038), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1041), .ZN(new_n1043));
  INV_X1    g618(.A(G8), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1045), .B1(new_n1032), .B2(new_n1038), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT51), .ZN(new_n1047));
  NOR3_X1   g622(.A1(new_n1042), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1032), .A2(new_n1038), .ZN(new_n1049));
  AOI211_X1 g624(.A(KEYINPUT51), .B(new_n1043), .C1(new_n1049), .C2(new_n1040), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1019), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  OAI211_X1 g626(.A(G160), .B(G40), .C1(new_n1025), .C2(KEYINPUT50), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1020), .B1(new_n884), .B2(new_n982), .ZN(new_n1053));
  NOR3_X1   g628(.A1(new_n1052), .A2(new_n1053), .A3(G2090), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n991), .B1(new_n884), .B2(new_n1035), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1025), .A2(new_n1034), .ZN(new_n1056));
  AOI21_X1  g631(.A(G1971), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1040), .B1(new_n1054), .B2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT115), .ZN(new_n1060));
  XNOR2_X1  g635(.A(new_n1059), .B(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(G303), .A2(G8), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT55), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT116), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT116), .ZN(new_n1065));
  AOI211_X1 g640(.A(new_n1065), .B(KEYINPUT55), .C1(G303), .C2(G8), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1061), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1058), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(G2090), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1023), .A2(new_n1070), .A3(new_n1031), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1072));
  INV_X1    g647(.A(G1971), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1044), .B1(new_n1071), .B2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(KEYINPUT117), .B1(new_n1061), .B2(new_n1067), .ZN(new_n1076));
  XNOR2_X1  g651(.A(new_n1059), .B(KEYINPUT115), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT117), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1077), .B(new_n1078), .C1(new_n1064), .C2(new_n1066), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1075), .A2(new_n1076), .A3(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(KEYINPUT114), .B1(new_n1025), .B2(KEYINPUT50), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n1028), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1022), .B(new_n1021), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1083));
  XOR2_X1   g658(.A(KEYINPUT122), .B(G1961), .Z(new_n1084));
  INV_X1    g659(.A(G2078), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1055), .A2(new_n1085), .A3(new_n1056), .ZN(new_n1086));
  XOR2_X1   g661(.A(KEYINPUT123), .B(KEYINPUT53), .Z(new_n1087));
  AOI22_X1  g662(.A1(new_n1083), .A2(new_n1084), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1085), .A2(KEYINPUT53), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n984), .A2(new_n1022), .A3(new_n1090), .A4(new_n1036), .ZN(new_n1091));
  AOI21_X1  g666(.A(G301), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n813), .A2(new_n704), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT82), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1094), .B1(new_n530), .B2(new_n595), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1095), .A2(new_n597), .A3(new_n599), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n1096), .A2(new_n508), .B1(G48), .B2(new_n534), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(new_n604), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(G1981), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1093), .A2(new_n1099), .A3(KEYINPUT49), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n884), .A2(new_n982), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1039), .B1(new_n1102), .B2(new_n1022), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT49), .ZN(new_n1104));
  NOR2_X1   g679(.A1(G305), .A2(G1981), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n704), .B1(new_n1097), .B2(new_n604), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1104), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1100), .A2(new_n1103), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n818), .A2(G1976), .ZN(new_n1109));
  INV_X1    g684(.A(G1976), .ZN(new_n1110));
  AOI21_X1  g685(.A(KEYINPUT52), .B1(G288), .B2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1103), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1109), .B(new_n1040), .C1(new_n1101), .C2(new_n991), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(KEYINPUT52), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n1108), .A2(new_n1112), .A3(new_n1114), .ZN(new_n1115));
  AND4_X1   g690(.A1(new_n1069), .A2(new_n1080), .A3(new_n1092), .A4(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1043), .A2(KEYINPUT51), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n1032), .A2(new_n1038), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1117), .B1(new_n1118), .B2(new_n1039), .ZN(new_n1119));
  OAI21_X1  g694(.A(KEYINPUT51), .B1(new_n1118), .B2(new_n1045), .ZN(new_n1120));
  OAI211_X1 g695(.A(KEYINPUT62), .B(new_n1119), .C1(new_n1120), .C2(new_n1042), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1051), .A2(new_n1116), .A3(new_n1121), .ZN(new_n1122));
  AOI211_X1 g697(.A(G286), .B(new_n1039), .C1(new_n1032), .C2(new_n1038), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1080), .A2(new_n1069), .A3(new_n1115), .A4(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT63), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  AND4_X1   g701(.A1(KEYINPUT63), .A2(new_n1049), .A3(G168), .A4(new_n1040), .ZN(new_n1127));
  AND2_X1   g702(.A1(new_n1071), .A2(new_n1074), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1068), .B1(new_n1128), .B2(new_n1044), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1127), .A2(new_n1129), .A3(new_n1080), .A4(new_n1115), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1126), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1080), .ZN(new_n1132));
  AND2_X1   g707(.A1(new_n1100), .A2(new_n1107), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n818), .A2(new_n1110), .ZN(new_n1134));
  XOR2_X1   g709(.A(new_n1134), .B(KEYINPUT119), .Z(new_n1135));
  OAI21_X1  g710(.A(new_n1093), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1136));
  AOI22_X1  g711(.A1(new_n1132), .A2(new_n1115), .B1(new_n1103), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1122), .A2(new_n1131), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT57), .ZN(new_n1139));
  NAND2_X1  g714(.A1(G299), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n917), .A2(KEYINPUT57), .A3(new_n574), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n770), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1143));
  XNOR2_X1  g718(.A(KEYINPUT56), .B(G2072), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1055), .A2(new_n1056), .A3(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1142), .A2(new_n1143), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(G1348), .B1(new_n1023), .B2(new_n1031), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1102), .A2(new_n728), .A3(new_n1022), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n628), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1142), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1147), .B1(new_n1151), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT121), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1146), .A2(new_n1156), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1142), .A2(new_n1143), .A3(KEYINPUT121), .A4(new_n1145), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1157), .A2(KEYINPUT61), .A3(new_n1154), .A4(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT60), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1160), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1083), .A2(new_n747), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1162), .A2(KEYINPUT60), .A3(new_n1149), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1161), .A2(new_n1163), .A3(new_n628), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1055), .A2(new_n993), .A3(new_n1056), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(KEYINPUT120), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT120), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1055), .A2(new_n1167), .A3(new_n993), .A4(new_n1056), .ZN(new_n1168));
  XOR2_X1   g743(.A(KEYINPUT58), .B(G1341), .Z(new_n1169));
  OAI21_X1  g744(.A(new_n1169), .B1(new_n1101), .B2(new_n991), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1166), .A2(new_n1168), .A3(new_n1170), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1171), .A2(KEYINPUT59), .A3(new_n564), .ZN(new_n1172));
  AND3_X1   g747(.A1(new_n1159), .A2(new_n1164), .A3(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(KEYINPUT61), .B1(new_n1154), .B2(new_n1146), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1163), .A2(new_n628), .ZN(new_n1175));
  AOI21_X1  g750(.A(KEYINPUT59), .B1(new_n1171), .B2(new_n564), .ZN(new_n1176));
  NOR3_X1   g751(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1155), .B1(new_n1173), .B2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1179));
  AND3_X1   g754(.A1(new_n1080), .A2(new_n1069), .A3(new_n1115), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n984), .A2(new_n1055), .A3(new_n1090), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1184), .A2(KEYINPUT126), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT126), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1186), .B1(new_n1088), .B2(new_n1183), .ZN(new_n1187));
  NOR3_X1   g762(.A1(new_n1185), .A2(new_n1187), .A3(G301), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1088), .A2(new_n1091), .ZN(new_n1189));
  OAI21_X1  g764(.A(KEYINPUT54), .B1(new_n1189), .B2(G171), .ZN(new_n1190));
  OAI211_X1 g765(.A(new_n1179), .B(new_n1180), .C1(new_n1188), .C2(new_n1190), .ZN(new_n1191));
  NOR2_X1   g766(.A1(new_n1178), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(new_n1092), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT124), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1194), .B1(new_n1184), .B2(G171), .ZN(new_n1195));
  NAND4_X1  g770(.A1(new_n1088), .A2(KEYINPUT124), .A3(G301), .A4(new_n1183), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1193), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT54), .ZN(new_n1198));
  AND3_X1   g773(.A1(new_n1197), .A2(KEYINPUT125), .A3(new_n1198), .ZN(new_n1199));
  AOI21_X1  g774(.A(KEYINPUT125), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1200));
  NOR2_X1   g775(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n1138), .B1(new_n1192), .B2(new_n1201), .ZN(new_n1202));
  NOR2_X1   g777(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1203));
  XNOR2_X1  g778(.A(G290), .B(new_n843), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n996), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1018), .B1(new_n1202), .B2(new_n1205), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g781(.A1(new_n978), .A2(new_n979), .ZN(new_n1208));
  NAND4_X1  g782(.A1(new_n688), .A2(new_n673), .A3(G319), .A4(new_n689), .ZN(new_n1209));
  INV_X1    g783(.A(new_n1209), .ZN(new_n1210));
  OAI211_X1 g784(.A(new_n712), .B(new_n1210), .C1(new_n907), .C2(new_n908), .ZN(new_n1211));
  NOR2_X1   g785(.A1(new_n1208), .A2(new_n1211), .ZN(G308));
  AOI21_X1  g786(.A(new_n1209), .B1(new_n710), .B2(new_n711), .ZN(new_n1213));
  OAI221_X1 g787(.A(new_n1213), .B1(new_n907), .B2(new_n908), .C1(new_n978), .C2(new_n979), .ZN(G225));
endmodule


