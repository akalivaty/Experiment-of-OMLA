//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 1 1 0 0 1 0 1 1 1 1 1 1 0 0 0 0 1 1 1 1 0 0 1 0 1 1 0 0 0 1 1 0 1 0 0 1 0 1 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:22 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n656,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937;
  XNOR2_X1  g000(.A(KEYINPUT73), .B(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT72), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT31), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT26), .B(G101), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n190), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G237), .ZN(new_n193));
  INV_X1    g007(.A(G953), .ZN(new_n194));
  AND3_X1   g008(.A1(new_n193), .A2(new_n194), .A3(G210), .ZN(new_n195));
  XOR2_X1   g009(.A(new_n192), .B(new_n195), .Z(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT11), .ZN(new_n198));
  INV_X1    g012(.A(G134), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(G137), .ZN(new_n200));
  INV_X1    g014(.A(G137), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(KEYINPUT11), .A3(G134), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n201), .A2(G134), .ZN(new_n204));
  OAI21_X1  g018(.A(G131), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(new_n204), .ZN(new_n206));
  INV_X1    g020(.A(G131), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n206), .A2(new_n207), .A3(new_n200), .A4(new_n202), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G143), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(KEYINPUT64), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G143), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n211), .B1(new_n215), .B2(G146), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(KEYINPUT0), .A3(G128), .ZN(new_n217));
  INV_X1    g031(.A(G146), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n212), .A2(new_n214), .A3(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n218), .A2(G143), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(KEYINPUT0), .A2(G128), .ZN(new_n223));
  OR2_X1    g037(.A1(KEYINPUT0), .A2(G128), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  AND3_X1   g039(.A1(new_n217), .A2(KEYINPUT66), .A3(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(KEYINPUT66), .B1(new_n217), .B2(new_n225), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n209), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  XOR2_X1   g043(.A(KEYINPUT2), .B(G113), .Z(new_n230));
  XNOR2_X1  g044(.A(G116), .B(G119), .ZN(new_n231));
  XNOR2_X1  g045(.A(new_n230), .B(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n218), .B1(new_n212), .B2(new_n214), .ZN(new_n236));
  INV_X1    g050(.A(G128), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n237), .A2(KEYINPUT1), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NOR3_X1   g053(.A1(new_n236), .A2(new_n211), .A3(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT1), .B1(new_n210), .B2(G146), .ZN(new_n241));
  AOI22_X1  g055(.A1(new_n219), .A2(new_n221), .B1(G128), .B2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n235), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n211), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT64), .B(G143), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n244), .B(new_n238), .C1(new_n245), .C2(new_n218), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n220), .B1(new_n245), .B2(new_n218), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n241), .A2(G128), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n246), .B(KEYINPUT67), .C1(new_n247), .C2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n243), .A2(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n199), .A2(G137), .ZN(new_n252));
  OAI21_X1  g066(.A(G131), .B1(new_n252), .B2(new_n204), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT65), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT65), .ZN(new_n255));
  OAI211_X1 g069(.A(new_n255), .B(G131), .C1(new_n252), .C2(new_n204), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n254), .A2(new_n208), .A3(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n234), .B1(new_n251), .B2(new_n258), .ZN(new_n259));
  AOI211_X1 g073(.A(KEYINPUT68), .B(new_n257), .C1(new_n243), .C2(new_n250), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n197), .B1(new_n233), .B2(new_n261), .ZN(new_n262));
  NOR3_X1   g076(.A1(new_n240), .A2(new_n242), .A3(new_n235), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n222), .A2(new_n248), .ZN(new_n264));
  AOI21_X1  g078(.A(KEYINPUT67), .B1(new_n264), .B2(new_n246), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n258), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(KEYINPUT68), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n251), .A2(new_n234), .A3(new_n258), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n267), .A2(KEYINPUT30), .A3(new_n228), .A4(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n269), .B(KEYINPUT69), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n217), .A2(new_n225), .ZN(new_n271));
  INV_X1    g085(.A(new_n209), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n240), .A2(new_n242), .ZN(new_n273));
  OAI22_X1  g087(.A1(new_n271), .A2(new_n272), .B1(new_n273), .B2(new_n257), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT30), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n232), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n189), .B(new_n262), .C1(new_n270), .C2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT69), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n269), .A2(new_n279), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n261), .A2(KEYINPUT69), .A3(KEYINPUT30), .A4(new_n228), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n277), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n262), .ZN(new_n283));
  OAI21_X1  g097(.A(KEYINPUT31), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT28), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n233), .A2(new_n261), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n274), .A2(new_n232), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(KEYINPUT28), .B1(new_n233), .B2(new_n266), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n197), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n278), .A2(new_n284), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT71), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n278), .A2(new_n284), .A3(new_n290), .A4(KEYINPUT71), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g109(.A1(G472), .A2(G902), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n188), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n296), .ZN(new_n298));
  AOI211_X1 g112(.A(KEYINPUT72), .B(new_n298), .C1(new_n293), .C2(new_n294), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n187), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n280), .A2(new_n281), .ZN(new_n301));
  INV_X1    g115(.A(new_n277), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n286), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n197), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT29), .ZN(new_n306));
  OR3_X1    g120(.A1(new_n288), .A2(new_n289), .A3(new_n197), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT74), .ZN(new_n309));
  INV_X1    g123(.A(G902), .ZN(new_n310));
  INV_X1    g124(.A(new_n261), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n232), .B1(new_n311), .B2(new_n229), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(new_n286), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n289), .B1(new_n313), .B2(KEYINPUT28), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n314), .A2(KEYINPUT29), .A3(new_n196), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT74), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n305), .A2(new_n316), .A3(new_n307), .A4(new_n306), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n309), .A2(new_n310), .A3(new_n315), .A4(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G472), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n298), .B1(new_n293), .B2(new_n294), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT32), .ZN(new_n322));
  OAI21_X1  g136(.A(KEYINPUT75), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT75), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n320), .A2(new_n324), .A3(KEYINPUT32), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n300), .A2(new_n319), .A3(new_n323), .A4(new_n325), .ZN(new_n326));
  XOR2_X1   g140(.A(KEYINPUT22), .B(G137), .Z(new_n327));
  NAND3_X1  g141(.A1(new_n194), .A2(G221), .A3(G234), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n327), .B(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(G125), .B(G140), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT16), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G125), .ZN(new_n333));
  OAI22_X1  g147(.A1(new_n331), .A2(new_n332), .B1(G140), .B2(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n334), .B(new_n218), .ZN(new_n335));
  INV_X1    g149(.A(G119), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n336), .A2(G128), .ZN(new_n337));
  OR2_X1    g151(.A1(new_n337), .A2(KEYINPUT23), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n336), .A2(G128), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n337), .A2(KEYINPUT23), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G110), .ZN(new_n342));
  INV_X1    g156(.A(new_n339), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n343), .A2(new_n337), .ZN(new_n344));
  XOR2_X1   g158(.A(KEYINPUT24), .B(G110), .Z(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n335), .A2(new_n342), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n330), .A2(new_n218), .ZN(new_n348));
  XOR2_X1   g162(.A(new_n348), .B(KEYINPUT77), .Z(new_n349));
  OR2_X1    g163(.A1(new_n334), .A2(new_n218), .ZN(new_n350));
  OAI22_X1  g164(.A1(new_n341), .A2(G110), .B1(new_n344), .B2(new_n345), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n329), .B1(new_n353), .B2(KEYINPUT78), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(KEYINPUT78), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n354), .B(new_n355), .ZN(new_n356));
  OR3_X1    g170(.A1(new_n356), .A2(KEYINPUT25), .A3(G902), .ZN(new_n357));
  XNOR2_X1  g171(.A(KEYINPUT76), .B(G217), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n359), .B1(G234), .B2(new_n310), .ZN(new_n360));
  OAI21_X1  g174(.A(KEYINPUT25), .B1(new_n356), .B2(G902), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n357), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n356), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n360), .A2(G902), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT6), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT86), .ZN(new_n369));
  XNOR2_X1  g183(.A(KEYINPUT80), .B(G107), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT3), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n370), .A2(new_n371), .A3(G104), .ZN(new_n372));
  INV_X1    g186(.A(G104), .ZN(new_n373));
  OAI21_X1  g187(.A(KEYINPUT3), .B1(new_n373), .B2(G107), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(G107), .ZN(new_n375));
  AND3_X1   g189(.A1(new_n372), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  XOR2_X1   g190(.A(KEYINPUT81), .B(G101), .Z(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n370), .A2(G104), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n373), .A2(G107), .ZN(new_n380));
  OAI21_X1  g194(.A(G101), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n231), .A2(KEYINPUT5), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n336), .A2(G116), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n383), .B(G113), .C1(KEYINPUT5), .C2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n230), .A2(new_n231), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n369), .B1(new_n382), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n387), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n389), .A2(new_n378), .A3(KEYINPUT86), .A4(new_n381), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(G101), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n378), .B(KEYINPUT4), .C1(new_n392), .C2(new_n376), .ZN(new_n393));
  OR3_X1    g207(.A1(new_n376), .A2(KEYINPUT4), .A3(new_n392), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n393), .A2(new_n232), .A3(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT85), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n393), .A2(KEYINPUT85), .A3(new_n232), .A4(new_n394), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n391), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  XOR2_X1   g213(.A(G110), .B(G122), .Z(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n368), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n402), .B1(new_n401), .B2(new_n399), .ZN(new_n403));
  INV_X1    g217(.A(new_n399), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n404), .A2(new_n368), .A3(new_n400), .ZN(new_n405));
  MUX2_X1   g219(.A(new_n273), .B(new_n271), .S(G125), .Z(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(G224), .A3(new_n194), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n406), .B1(G224), .B2(new_n194), .ZN(new_n409));
  OR2_X1    g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n403), .A2(new_n405), .A3(new_n410), .ZN(new_n411));
  XOR2_X1   g225(.A(new_n400), .B(KEYINPUT8), .Z(new_n412));
  NOR2_X1   g226(.A1(new_n382), .A2(new_n387), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n389), .B1(new_n378), .B2(new_n381), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n407), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n416), .B1(KEYINPUT7), .B2(new_n409), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT7), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n406), .A2(new_n418), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n417), .B(new_n419), .C1(new_n400), .C2(new_n404), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n411), .A2(new_n310), .A3(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(G210), .B1(G237), .B2(G902), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n411), .A2(new_n310), .A3(new_n420), .A4(new_n422), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(G214), .B1(G237), .B2(G902), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n427), .B(KEYINPUT84), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  XNOR2_X1  g244(.A(KEYINPUT9), .B(G234), .ZN(new_n431));
  XOR2_X1   g245(.A(new_n431), .B(KEYINPUT79), .Z(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(G221), .B1(new_n433), .B2(G902), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n393), .B(new_n394), .C1(new_n227), .C2(new_n226), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n237), .B1(new_n219), .B2(KEYINPUT1), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n246), .B1(new_n437), .B2(new_n216), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n378), .A2(new_n381), .A3(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT10), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n251), .A2(KEYINPUT10), .A3(new_n378), .A4(new_n381), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n436), .A2(new_n272), .A3(new_n441), .A4(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(G110), .B(G140), .ZN(new_n444));
  AND2_X1   g258(.A1(new_n194), .A2(G227), .ZN(new_n445));
  XOR2_X1   g259(.A(new_n444), .B(new_n445), .Z(new_n446));
  NAND2_X1  g260(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(KEYINPUT82), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n436), .A2(new_n441), .A3(new_n442), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n209), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT82), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n443), .A2(new_n451), .A3(new_n446), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n448), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n382), .A2(new_n273), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n272), .B1(new_n454), .B2(new_n439), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(KEYINPUT12), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n443), .ZN(new_n457));
  INV_X1    g271(.A(new_n446), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(G469), .B1(new_n461), .B2(G902), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n447), .A2(KEYINPUT83), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT83), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n443), .A2(new_n464), .A3(new_n446), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n463), .A2(new_n456), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n450), .A2(new_n443), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n458), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(G469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n469), .A2(new_n470), .A3(new_n310), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n435), .B1(new_n462), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(G475), .ZN(new_n474));
  XNOR2_X1  g288(.A(G113), .B(G122), .ZN(new_n475));
  XNOR2_X1  g289(.A(KEYINPUT92), .B(G104), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n475), .B(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n193), .A2(new_n194), .A3(G214), .ZN(new_n479));
  OR2_X1    g293(.A1(new_n479), .A2(G143), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n245), .A2(new_n479), .ZN(new_n481));
  AOI21_X1  g295(.A(G131), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n480), .A2(new_n481), .A3(G131), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n483), .A2(KEYINPUT88), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n480), .A2(new_n481), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT88), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n486), .A2(new_n487), .A3(new_n207), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  OR2_X1    g303(.A1(new_n489), .A2(KEYINPUT89), .ZN(new_n490));
  XNOR2_X1  g304(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n331), .A2(new_n491), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n492), .A2(KEYINPUT91), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n492), .A2(KEYINPUT91), .ZN(new_n494));
  AND2_X1   g308(.A1(new_n331), .A2(KEYINPUT19), .ZN(new_n495));
  NOR3_X1   g309(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n218), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n489), .A2(KEYINPUT89), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n490), .A2(new_n350), .A3(new_n497), .A4(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n349), .B1(new_n218), .B2(new_n330), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT18), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n486), .B1(new_n501), .B2(new_n207), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n500), .B(new_n502), .C1(new_n501), .C2(new_n484), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n478), .B1(new_n499), .B2(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n334), .B(G146), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT93), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT17), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n505), .B(new_n506), .C1(new_n507), .C2(new_n484), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n484), .A2(new_n507), .ZN(new_n509));
  OAI21_X1  g323(.A(KEYINPUT93), .B1(new_n335), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(KEYINPUT17), .B1(new_n485), .B2(new_n488), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n478), .B(new_n503), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n474), .B(new_n310), .C1(new_n504), .C2(new_n514), .ZN(new_n515));
  OR2_X1    g329(.A1(new_n515), .A2(KEYINPUT20), .ZN(new_n516));
  XOR2_X1   g330(.A(KEYINPUT87), .B(KEYINPUT20), .Z(new_n517));
  NAND2_X1  g331(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n503), .B1(new_n511), .B2(new_n512), .ZN(new_n519));
  AND2_X1   g333(.A1(new_n519), .A2(new_n477), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(KEYINPUT94), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT94), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n513), .A2(new_n522), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n521), .B(new_n310), .C1(new_n520), .C2(new_n523), .ZN(new_n524));
  AOI22_X1  g338(.A1(new_n516), .A2(new_n518), .B1(new_n524), .B2(G475), .ZN(new_n525));
  INV_X1    g339(.A(G122), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(G116), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n527), .B(KEYINPUT95), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n526), .A2(G116), .ZN(new_n529));
  OR2_X1    g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n370), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n530), .B(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n237), .A2(G143), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n533), .B1(new_n245), .B2(new_n237), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n534), .A2(G134), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT13), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n215), .A2(new_n537), .A3(G128), .ZN(new_n538));
  OAI211_X1 g352(.A(G134), .B(new_n538), .C1(new_n534), .C2(new_n537), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n532), .A2(new_n536), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n534), .A2(G134), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  OR3_X1    g356(.A1(new_n542), .A2(KEYINPUT96), .A3(new_n535), .ZN(new_n543));
  OR2_X1    g357(.A1(new_n530), .A2(new_n531), .ZN(new_n544));
  XOR2_X1   g358(.A(new_n529), .B(KEYINPUT14), .Z(new_n545));
  OAI21_X1  g359(.A(G107), .B1(new_n545), .B2(new_n528), .ZN(new_n546));
  OAI21_X1  g360(.A(KEYINPUT96), .B1(new_n542), .B2(new_n535), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n543), .A2(new_n544), .A3(new_n546), .A4(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n540), .A2(new_n548), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n433), .A2(G953), .A3(new_n359), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT97), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n540), .A2(new_n548), .A3(new_n550), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n549), .A2(KEYINPUT97), .A3(new_n551), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n555), .A2(KEYINPUT98), .A3(new_n310), .A4(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT15), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(G478), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  OR2_X1    g374(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n557), .A2(new_n560), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n194), .A2(G952), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n565), .B1(G234), .B2(G237), .ZN(new_n566));
  XOR2_X1   g380(.A(KEYINPUT21), .B(G898), .Z(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(G234), .A2(G237), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n569), .A2(G902), .A3(G953), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n566), .B1(new_n568), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n525), .A2(new_n564), .A3(new_n573), .ZN(new_n574));
  NOR3_X1   g388(.A1(new_n430), .A2(new_n473), .A3(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n326), .A2(new_n367), .A3(new_n575), .ZN(new_n576));
  XOR2_X1   g390(.A(new_n576), .B(new_n377), .Z(G3));
  INV_X1    g391(.A(G472), .ZN(new_n578));
  AOI21_X1  g392(.A(G902), .B1(new_n293), .B2(new_n294), .ZN(new_n579));
  OAI22_X1  g393(.A1(new_n297), .A2(new_n299), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n581), .A2(new_n367), .A3(new_n472), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n424), .A2(KEYINPUT99), .A3(new_n425), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT99), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n421), .A2(new_n585), .A3(new_n423), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n584), .A2(new_n429), .A3(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT33), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n555), .A2(new_n589), .A3(new_n556), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n552), .A2(KEYINPUT33), .A3(new_n554), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n590), .A2(G478), .A3(new_n310), .A4(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n555), .A2(new_n310), .A3(new_n556), .ZN(new_n593));
  XOR2_X1   g407(.A(KEYINPUT100), .B(G478), .Z(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n525), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n599), .A2(new_n572), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n583), .A2(new_n588), .A3(new_n600), .ZN(new_n601));
  XOR2_X1   g415(.A(KEYINPUT34), .B(G104), .Z(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(G6));
  OR2_X1    g417(.A1(new_n515), .A2(new_n517), .ZN(new_n604));
  AOI22_X1  g418(.A1(new_n604), .A2(new_n518), .B1(G475), .B2(new_n524), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n605), .A2(new_n563), .A3(new_n573), .ZN(new_n606));
  XOR2_X1   g420(.A(new_n606), .B(KEYINPUT101), .Z(new_n607));
  NAND3_X1  g421(.A1(new_n583), .A2(new_n588), .A3(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(G107), .ZN(new_n609));
  XNOR2_X1  g423(.A(KEYINPUT102), .B(KEYINPUT35), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(G9));
  NOR2_X1   g425(.A1(new_n329), .A2(KEYINPUT36), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n353), .B(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n364), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n362), .A2(new_n614), .ZN(new_n615));
  XOR2_X1   g429(.A(new_n615), .B(KEYINPUT103), .Z(new_n616));
  NAND3_X1  g430(.A1(new_n575), .A2(new_n581), .A3(new_n616), .ZN(new_n617));
  XOR2_X1   g431(.A(KEYINPUT37), .B(G110), .Z(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G12));
  NOR2_X1   g433(.A1(new_n587), .A2(new_n473), .ZN(new_n620));
  INV_X1    g434(.A(new_n566), .ZN(new_n621));
  OR2_X1    g435(.A1(new_n570), .A2(G900), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n605), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n624), .A2(new_n564), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n326), .A2(new_n616), .A3(new_n620), .A4(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(G128), .ZN(G30));
  XOR2_X1   g441(.A(new_n623), .B(KEYINPUT39), .Z(new_n628));
  OR2_X1    g442(.A1(new_n473), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(new_n629), .B(KEYINPUT40), .Z(new_n630));
  INV_X1    g444(.A(new_n304), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n631), .A2(new_n197), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n310), .B1(new_n313), .B2(new_n196), .ZN(new_n633));
  OAI21_X1  g447(.A(G472), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n300), .A2(new_n325), .A3(new_n323), .A4(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n636), .A2(new_n615), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n424), .A2(KEYINPUT38), .A3(new_n425), .ZN(new_n638));
  AOI21_X1  g452(.A(KEYINPUT38), .B1(new_n424), .B2(new_n425), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n525), .A2(new_n564), .A3(new_n428), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n630), .A2(new_n637), .A3(new_n640), .A4(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(new_n245), .ZN(G45));
  NAND2_X1  g457(.A1(new_n598), .A2(new_n623), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n326), .A2(new_n616), .A3(new_n620), .A4(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G146), .ZN(G48));
  INV_X1    g461(.A(new_n471), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n470), .B1(new_n469), .B2(new_n310), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n434), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n587), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n326), .A2(new_n367), .A3(new_n600), .A4(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT41), .B(G113), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G15));
  NAND4_X1  g469(.A1(new_n326), .A2(new_n607), .A3(new_n367), .A4(new_n652), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G116), .ZN(G18));
  INV_X1    g471(.A(new_n574), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n326), .A2(new_n658), .A3(new_n616), .A4(new_n652), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G119), .ZN(G21));
  AND4_X1   g474(.A1(new_n573), .A2(new_n641), .A3(new_n586), .A4(new_n584), .ZN(new_n661));
  INV_X1    g475(.A(new_n651), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n579), .A2(new_n578), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n278), .B(new_n284), .C1(new_n314), .C2(new_n196), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n663), .B1(new_n296), .B2(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n661), .A2(new_n367), .A3(new_n662), .A4(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G122), .ZN(G24));
  NAND2_X1  g481(.A1(new_n664), .A2(new_n296), .ZN(new_n668));
  OAI211_X1 g482(.A(new_n615), .B(new_n668), .C1(new_n579), .C2(new_n578), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT104), .ZN(new_n670));
  OR2_X1    g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n669), .A2(new_n670), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n673), .A2(new_n645), .A3(new_n652), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G125), .ZN(G27));
  NAND2_X1  g489(.A1(new_n320), .A2(KEYINPUT32), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n321), .A2(new_n322), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n319), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n367), .ZN(new_n679));
  AND3_X1   g493(.A1(new_n424), .A2(new_n429), .A3(new_n425), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n645), .A2(KEYINPUT42), .A3(new_n472), .A4(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT42), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n680), .A2(new_n472), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n684), .A2(new_n644), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n326), .A2(new_n367), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n682), .B1(new_n683), .B2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(new_n207), .ZN(G33));
  NOR3_X1   g502(.A1(new_n684), .A2(new_n564), .A3(new_n624), .ZN(new_n689));
  AND3_X1   g503(.A1(new_n689), .A2(new_n326), .A3(new_n367), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(new_n199), .ZN(G36));
  NAND2_X1  g505(.A1(new_n516), .A2(new_n518), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n524), .A2(G475), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n694), .A2(new_n597), .A3(KEYINPUT43), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT105), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n525), .A2(KEYINPUT105), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n697), .A2(new_n596), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n695), .B1(new_n699), .B2(KEYINPUT43), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n580), .A2(KEYINPUT106), .A3(new_n615), .ZN(new_n701));
  AOI21_X1  g515(.A(KEYINPUT106), .B1(new_n580), .B2(new_n615), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n700), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  OAI211_X1 g519(.A(KEYINPUT44), .B(new_n700), .C1(new_n701), .C2(new_n702), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n705), .A2(new_n680), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(KEYINPUT107), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT45), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n460), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n453), .A2(new_n459), .A3(KEYINPUT45), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n710), .A2(G469), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(G469), .A2(G902), .ZN(new_n713));
  AOI21_X1  g527(.A(KEYINPUT46), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n714), .A2(new_n648), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n712), .A2(KEYINPUT46), .A3(new_n713), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n434), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n718), .A2(new_n628), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT107), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n705), .A2(new_n720), .A3(new_n680), .A4(new_n706), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n708), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G137), .ZN(G39));
  INV_X1    g537(.A(KEYINPUT47), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n724), .A2(KEYINPUT108), .ZN(new_n725));
  AND2_X1   g539(.A1(new_n724), .A2(KEYINPUT108), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n725), .B1(new_n718), .B2(new_n727), .ZN(new_n728));
  AOI211_X1 g542(.A(KEYINPUT108), .B(new_n724), .C1(new_n717), .C2(new_n434), .ZN(new_n729));
  OR2_X1    g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OR2_X1    g544(.A1(new_n326), .A2(new_n367), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n645), .A2(new_n680), .ZN(new_n732));
  OAI21_X1  g546(.A(KEYINPUT109), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OR4_X1    g547(.A1(KEYINPUT109), .A2(new_n326), .A3(new_n367), .A4(new_n732), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n730), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  XOR2_X1   g549(.A(new_n735), .B(G140), .Z(G42));
  INV_X1    g550(.A(KEYINPUT52), .ZN(new_n737));
  INV_X1    g551(.A(new_n615), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n641), .A2(new_n586), .A3(new_n584), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n472), .A2(new_n623), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n635), .A2(new_n738), .A3(new_n739), .A4(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT112), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n674), .A2(new_n626), .A3(new_n646), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n737), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n742), .B(KEYINPUT112), .ZN(new_n747));
  AND3_X1   g561(.A1(new_n674), .A2(new_n626), .A3(new_n646), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n747), .A2(KEYINPUT52), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n576), .A2(new_n617), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT110), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n563), .B(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n598), .B1(new_n753), .B2(new_n525), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n754), .A2(new_n430), .A3(new_n572), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n751), .B1(new_n583), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n656), .A2(new_n659), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n653), .A2(new_n666), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  AOI211_X1 g573(.A(new_n644), .B(new_n684), .C1(new_n671), .C2(new_n672), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n684), .A2(new_n624), .A3(new_n753), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(new_n326), .A3(new_n616), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(KEYINPUT111), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT111), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n761), .A2(new_n326), .A3(new_n764), .A4(new_n616), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n760), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n686), .A2(new_n683), .ZN(new_n767));
  INV_X1    g581(.A(new_n682), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n690), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  AND4_X1   g583(.A1(new_n756), .A2(new_n759), .A3(new_n766), .A4(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n750), .A2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT53), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(KEYINPUT53), .B1(new_n750), .B2(new_n770), .ZN(new_n774));
  OAI21_X1  g588(.A(KEYINPUT54), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  XOR2_X1   g589(.A(new_n565), .B(KEYINPUT117), .Z(new_n776));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n650), .A2(new_n435), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n778), .B1(new_n728), .B2(new_n729), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n700), .A2(new_n566), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n665), .A2(new_n367), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n779), .A2(new_n680), .A3(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n779), .A2(KEYINPUT114), .A3(new_n680), .A4(new_n782), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n651), .A2(new_n428), .A3(new_n426), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n636), .A2(new_n367), .A3(new_n566), .A4(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n525), .A2(new_n597), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n700), .A2(new_n566), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n662), .B(new_n428), .C1(new_n638), .C2(new_n639), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n781), .ZN(new_n795));
  OR2_X1    g609(.A1(KEYINPUT115), .A2(KEYINPUT50), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n792), .A2(new_n794), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n780), .A2(new_n781), .A3(new_n793), .ZN(new_n798));
  XOR2_X1   g612(.A(KEYINPUT115), .B(KEYINPUT50), .Z(new_n799));
  OAI21_X1  g613(.A(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n792), .A2(new_n673), .A3(new_n788), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n791), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n777), .B1(new_n787), .B2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT116), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n791), .A2(new_n800), .A3(KEYINPUT116), .A4(new_n801), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n805), .A2(KEYINPUT51), .A3(new_n783), .A4(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n792), .A2(new_n367), .A3(new_n678), .A4(new_n788), .ZN(new_n808));
  XOR2_X1   g622(.A(new_n808), .B(KEYINPUT48), .Z(new_n809));
  NAND2_X1  g623(.A1(new_n782), .A2(new_n652), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n810), .B1(new_n789), .B2(new_n599), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  AND4_X1   g626(.A1(new_n776), .A2(new_n803), .A3(new_n807), .A4(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n771), .A2(new_n772), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT113), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n816), .B1(new_n757), .B2(new_n758), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(KEYINPUT53), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n757), .A2(new_n758), .A3(new_n816), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n756), .A2(new_n766), .A3(new_n769), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n750), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n814), .A2(new_n815), .A3(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n775), .A2(new_n813), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(KEYINPUT118), .ZN(new_n825));
  OR2_X1    g639(.A1(G952), .A2(G953), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT118), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n775), .A2(new_n813), .A3(new_n827), .A4(new_n823), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n825), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n367), .A2(new_n429), .ZN(new_n830));
  NOR4_X1   g644(.A1(new_n640), .A2(new_n699), .A3(new_n435), .A4(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n650), .B(KEYINPUT49), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n831), .A2(new_n636), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n829), .A2(new_n833), .ZN(G75));
  NOR2_X1   g648(.A1(new_n194), .A2(G952), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n750), .A2(new_n820), .A3(new_n821), .ZN(new_n836));
  OAI211_X1 g650(.A(G210), .B(G902), .C1(new_n836), .C2(new_n774), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT56), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n403), .A2(new_n405), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n840), .B(new_n410), .ZN(new_n841));
  XOR2_X1   g655(.A(new_n841), .B(KEYINPUT55), .Z(new_n842));
  AOI21_X1  g656(.A(new_n835), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  XOR2_X1   g657(.A(new_n842), .B(KEYINPUT119), .Z(new_n844));
  NAND3_X1  g658(.A1(new_n837), .A2(new_n838), .A3(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT120), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n837), .A2(KEYINPUT120), .A3(new_n838), .A4(new_n844), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n843), .A2(new_n847), .A3(new_n848), .ZN(G51));
  XOR2_X1   g663(.A(new_n713), .B(KEYINPUT57), .Z(new_n850));
  INV_X1    g664(.A(new_n823), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n815), .B1(new_n814), .B2(new_n822), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  XOR2_X1   g667(.A(new_n469), .B(KEYINPUT121), .Z(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n836), .A2(new_n774), .ZN(new_n856));
  OR3_X1    g670(.A1(new_n856), .A2(new_n310), .A3(new_n712), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n835), .B1(new_n855), .B2(new_n857), .ZN(G54));
  OAI211_X1 g672(.A(KEYINPUT58), .B(G902), .C1(new_n836), .C2(new_n774), .ZN(new_n859));
  OR2_X1    g673(.A1(new_n504), .A2(new_n514), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  OR3_X1    g675(.A1(new_n859), .A2(new_n474), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n861), .B1(new_n859), .B2(new_n474), .ZN(new_n863));
  INV_X1    g677(.A(new_n835), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(G60));
  NAND2_X1  g679(.A1(new_n590), .A2(new_n591), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n775), .A2(new_n823), .ZN(new_n868));
  NAND2_X1  g682(.A1(G478), .A2(G902), .ZN(new_n869));
  XOR2_X1   g683(.A(new_n869), .B(KEYINPUT59), .Z(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n867), .B1(new_n868), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n867), .A2(new_n871), .ZN(new_n873));
  INV_X1    g687(.A(new_n852), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n873), .B1(new_n874), .B2(new_n823), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n872), .A2(new_n875), .A3(new_n835), .ZN(G63));
  NAND2_X1  g690(.A1(G217), .A2(G902), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n877), .B(KEYINPUT60), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n878), .B1(new_n814), .B2(new_n822), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n835), .B1(new_n879), .B2(new_n613), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n356), .B1(new_n856), .B2(new_n878), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT61), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n880), .B(new_n881), .C1(KEYINPUT122), .C2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n878), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n613), .B(new_n884), .C1(new_n836), .C2(new_n774), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n885), .B(new_n864), .C1(new_n879), .C2(new_n363), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n885), .A2(KEYINPUT122), .A3(new_n864), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n886), .A2(KEYINPUT61), .A3(new_n887), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n883), .A2(new_n888), .ZN(G66));
  AOI21_X1  g703(.A(new_n194), .B1(new_n567), .B2(G224), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n756), .A2(new_n759), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n890), .B1(new_n891), .B2(new_n194), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n840), .B1(G898), .B2(new_n194), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT123), .Z(new_n894));
  XNOR2_X1  g708(.A(new_n892), .B(new_n894), .ZN(G69));
  NAND2_X1  g709(.A1(new_n301), .A2(new_n276), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n896), .B(new_n496), .Z(new_n897));
  INV_X1    g711(.A(KEYINPUT126), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n719), .A2(new_n739), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n748), .B1(new_n679), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n735), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n769), .A2(KEYINPUT125), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT125), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n903), .B1(new_n687), .B2(new_n690), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n722), .A2(new_n901), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n194), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n194), .A2(G900), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n898), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  AOI211_X1 g724(.A(KEYINPUT126), .B(new_n908), .C1(new_n906), .C2(new_n194), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n897), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n194), .B1(G227), .B2(G900), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT127), .ZN(new_n914));
  INV_X1    g728(.A(new_n735), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n642), .A2(new_n748), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(KEYINPUT62), .Z(new_n917));
  INV_X1    g731(.A(KEYINPUT124), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n326), .A2(new_n367), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n919), .A2(new_n629), .A3(new_n754), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n680), .ZN(new_n921));
  AND3_X1   g735(.A1(new_n722), .A2(new_n918), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n918), .B1(new_n722), .B2(new_n921), .ZN(new_n923));
  OAI211_X1 g737(.A(new_n915), .B(new_n917), .C1(new_n922), .C2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(new_n897), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n924), .A2(new_n194), .A3(new_n925), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n912), .A2(new_n914), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n914), .B1(new_n912), .B2(new_n926), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n927), .A2(new_n928), .ZN(G72));
  NAND2_X1  g743(.A1(G472), .A2(G902), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT63), .Z(new_n931));
  OAI21_X1  g745(.A(new_n305), .B1(new_n282), .B2(new_n283), .ZN(new_n932));
  OAI211_X1 g746(.A(new_n931), .B(new_n932), .C1(new_n773), .C2(new_n774), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n931), .B1(new_n906), .B2(new_n891), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n934), .A2(new_n197), .A3(new_n631), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n933), .A2(new_n935), .A3(new_n864), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n931), .B1(new_n924), .B2(new_n891), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n936), .B1(new_n632), .B2(new_n937), .ZN(G57));
endmodule


