//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 1 1 0 0 1 0 1 1 1 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 0 0 0 1 1 0 0 1 0 0 1 0 0 0 1 1 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:04 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n566,
    new_n567, new_n568, new_n569, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n604, new_n605,
    new_n606, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n638,
    new_n639, new_n640, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n824, new_n825, new_n826, new_n827, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916;
  XOR2_X1   g000(.A(KEYINPUT2), .B(G113), .Z(new_n187));
  XNOR2_X1  g001(.A(G116), .B(G119), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT67), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n187), .B(KEYINPUT66), .ZN(new_n192));
  INV_X1    g006(.A(new_n188), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n191), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G104), .ZN(new_n196));
  OAI21_X1  g010(.A(KEYINPUT3), .B1(new_n196), .B2(G107), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT3), .ZN(new_n198));
  INV_X1    g012(.A(G107), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n198), .A2(new_n199), .A3(G104), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n197), .B(new_n200), .C1(G104), .C2(new_n199), .ZN(new_n201));
  XNOR2_X1  g015(.A(KEYINPUT81), .B(G101), .ZN(new_n202));
  OR2_X1    g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(G101), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n203), .A2(KEYINPUT4), .A3(new_n204), .ZN(new_n205));
  OR2_X1    g019(.A1(new_n204), .A2(KEYINPUT4), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n195), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n199), .A2(G104), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n196), .A2(G107), .ZN(new_n209));
  OAI21_X1  g023(.A(G101), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  AND2_X1   g024(.A1(new_n203), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT5), .ZN(new_n212));
  INV_X1    g026(.A(G119), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(new_n213), .A3(G116), .ZN(new_n214));
  OAI211_X1 g028(.A(G113), .B(new_n214), .C1(new_n193), .C2(new_n212), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n211), .A2(new_n191), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n207), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(G110), .B(G122), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n207), .A2(new_n216), .A3(new_n218), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(KEYINPUT6), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT6), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n217), .A2(new_n223), .A3(new_n219), .ZN(new_n224));
  AND2_X1   g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G146), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G143), .ZN(new_n227));
  INV_X1    g041(.A(G143), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G146), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G128), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n226), .A2(G143), .ZN(new_n232));
  AOI22_X1  g046(.A1(new_n230), .A2(new_n231), .B1(KEYINPUT1), .B2(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(G143), .B(G146), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT1), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n234), .A2(new_n235), .A3(G128), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G125), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  XOR2_X1   g054(.A(KEYINPUT0), .B(G128), .Z(new_n241));
  OR2_X1    g055(.A1(new_n241), .A2(new_n234), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT0), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n234), .B1(new_n243), .B2(new_n231), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n240), .B1(new_n239), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G953), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G224), .ZN(new_n248));
  XOR2_X1   g062(.A(new_n246), .B(new_n248), .Z(new_n249));
  NAND3_X1  g063(.A1(new_n225), .A2(KEYINPUT85), .A3(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n222), .A2(new_n224), .A3(new_n249), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT85), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT7), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n248), .A2(KEYINPUT87), .ZN(new_n255));
  OR2_X1    g069(.A1(new_n248), .A2(KEYINPUT87), .ZN(new_n256));
  AOI211_X1 g070(.A(new_n254), .B(new_n246), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  XOR2_X1   g071(.A(new_n218), .B(KEYINPUT8), .Z(new_n258));
  INV_X1    g072(.A(new_n211), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n191), .A2(new_n215), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n258), .B1(new_n261), .B2(new_n216), .ZN(new_n262));
  AND2_X1   g076(.A1(new_n254), .A2(KEYINPUT86), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n254), .A2(KEYINPUT86), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n248), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  AND2_X1   g079(.A1(new_n246), .A2(new_n265), .ZN(new_n266));
  NOR3_X1   g080(.A1(new_n257), .A2(new_n262), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(G902), .B1(new_n267), .B2(new_n221), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n250), .A2(new_n253), .A3(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(G210), .B1(G237), .B2(G902), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n269), .B(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(G214), .B1(G237), .B2(G902), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(G122), .ZN(new_n275));
  AND2_X1   g089(.A1(new_n275), .A2(G116), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n275), .A2(G116), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n278), .B(new_n199), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n231), .A2(G143), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(KEYINPUT13), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n228), .A2(G128), .ZN(new_n282));
  MUX2_X1   g096(.A(KEYINPUT13), .B(new_n281), .S(new_n282), .Z(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G134), .ZN(new_n284));
  XNOR2_X1  g098(.A(KEYINPUT64), .B(G134), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n282), .A2(new_n280), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n279), .B(new_n284), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n278), .A2(new_n199), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n286), .B(new_n285), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n276), .A2(KEYINPUT14), .ZN(new_n290));
  MUX2_X1   g104(.A(new_n290), .B(KEYINPUT14), .S(new_n277), .Z(new_n291));
  OAI211_X1 g105(.A(new_n288), .B(new_n289), .C1(new_n291), .C2(new_n199), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n287), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g107(.A(KEYINPUT9), .B(G234), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(G217), .A3(new_n247), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n293), .B(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G902), .ZN(new_n298));
  AND2_X1   g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT92), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G478), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n302), .A2(KEYINPUT15), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n301), .B(new_n303), .ZN(new_n304));
  OR2_X1    g118(.A1(KEYINPUT93), .A2(G952), .ZN(new_n305));
  NAND2_X1  g119(.A1(KEYINPUT93), .A2(G952), .ZN(new_n306));
  AOI21_X1  g120(.A(G953), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G234), .ZN(new_n308));
  INV_X1    g122(.A(G237), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT21), .B(G898), .ZN(new_n312));
  AOI211_X1 g126(.A(new_n298), .B(new_n247), .C1(G234), .C2(G237), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n309), .A2(new_n247), .A3(G214), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n315), .B(G143), .ZN(new_n316));
  INV_X1    g130(.A(G131), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(KEYINPUT18), .A2(G131), .ZN(new_n319));
  AOI22_X1  g133(.A1(new_n318), .A2(KEYINPUT18), .B1(new_n316), .B2(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(G125), .B(G140), .ZN(new_n321));
  XNOR2_X1  g135(.A(new_n321), .B(KEYINPUT78), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n226), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT77), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n239), .A2(KEYINPUT77), .A3(G140), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n323), .B1(new_n226), .B2(new_n327), .ZN(new_n328));
  AND2_X1   g142(.A1(new_n328), .A2(KEYINPUT88), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n328), .A2(KEYINPUT88), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n320), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NOR3_X1   g145(.A1(new_n239), .A2(KEYINPUT16), .A3(G140), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n332), .B1(new_n327), .B2(KEYINPUT16), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n333), .B(new_n226), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n318), .A2(KEYINPUT17), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n316), .B(new_n317), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n334), .B(new_n335), .C1(KEYINPUT17), .C2(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(G113), .B(G122), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n338), .B(new_n196), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n331), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n339), .B1(new_n331), .B2(new_n337), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n298), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G475), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n328), .B(KEYINPUT88), .ZN(new_n345));
  XNOR2_X1  g159(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n322), .A2(new_n346), .ZN(new_n347));
  OR2_X1    g161(.A1(new_n347), .A2(KEYINPUT90), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(KEYINPUT90), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n325), .A2(KEYINPUT19), .A3(new_n326), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n348), .A2(new_n226), .A3(new_n349), .A4(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n333), .A2(G146), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n336), .A2(new_n352), .ZN(new_n353));
  AOI22_X1  g167(.A1(new_n345), .A2(new_n320), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n340), .B1(new_n354), .B2(new_n339), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT20), .ZN(new_n356));
  NOR2_X1   g170(.A1(G475), .A2(G902), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n356), .B1(new_n355), .B2(new_n357), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n344), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT91), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  OAI211_X1 g177(.A(KEYINPUT91), .B(new_n344), .C1(new_n359), .C2(new_n360), .ZN(new_n364));
  AOI211_X1 g178(.A(new_n304), .B(new_n314), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G221), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n366), .B1(new_n295), .B2(new_n298), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT10), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT82), .ZN(new_n369));
  OR2_X1    g183(.A1(new_n236), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n236), .A2(new_n369), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n370), .A2(new_n233), .A3(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT83), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n211), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n373), .B1(new_n211), .B2(new_n372), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n368), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G137), .ZN(new_n378));
  AND3_X1   g192(.A1(new_n378), .A2(KEYINPUT11), .A3(G134), .ZN(new_n379));
  AND2_X1   g193(.A1(KEYINPUT64), .A2(G134), .ZN(new_n380));
  NOR2_X1   g194(.A1(KEYINPUT64), .A2(G134), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n379), .B1(new_n382), .B2(G137), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n378), .B1(new_n380), .B2(new_n381), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT11), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n383), .A2(new_n386), .A3(new_n317), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT65), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n383), .A2(new_n386), .A3(KEYINPUT65), .A4(new_n317), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n383), .A2(new_n386), .ZN(new_n391));
  AOI22_X1  g205(.A1(new_n389), .A2(new_n390), .B1(G131), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n211), .A2(KEYINPUT10), .A3(new_n237), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n205), .A2(new_n206), .A3(new_n245), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n377), .A2(new_n392), .A3(new_n393), .A4(new_n394), .ZN(new_n395));
  OAI22_X1  g209(.A1(new_n375), .A2(new_n376), .B1(new_n211), .B2(new_n237), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n391), .A2(G131), .ZN(new_n397));
  AOI21_X1  g211(.A(KEYINPUT11), .B1(new_n285), .B2(new_n378), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT64), .ZN(new_n399));
  INV_X1    g213(.A(G134), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(KEYINPUT64), .A2(G134), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n401), .A2(G137), .A3(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n378), .A2(KEYINPUT11), .A3(G134), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n398), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(KEYINPUT65), .B1(new_n406), .B2(new_n317), .ZN(new_n407));
  INV_X1    g221(.A(new_n390), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n397), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n396), .A2(KEYINPUT12), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(KEYINPUT12), .B1(new_n396), .B2(new_n409), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n395), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(G110), .B(G140), .ZN(new_n413));
  AND2_X1   g227(.A1(new_n247), .A2(G227), .ZN(new_n414));
  XOR2_X1   g228(.A(new_n413), .B(new_n414), .Z(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n211), .A2(new_n372), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(KEYINPUT83), .ZN(new_n419));
  AOI21_X1  g233(.A(KEYINPUT10), .B1(new_n419), .B2(new_n374), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n393), .A2(new_n394), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n409), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n395), .A2(new_n422), .A3(new_n415), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n417), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n298), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(G469), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n412), .A2(new_n415), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n395), .A2(new_n422), .A3(new_n416), .ZN(new_n428));
  XNOR2_X1  g242(.A(KEYINPUT84), .B(G469), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n427), .A2(new_n298), .A3(new_n428), .A4(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n367), .B1(new_n426), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n274), .A2(new_n365), .A3(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT70), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT30), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n409), .A2(new_n245), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n389), .A2(new_n390), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n384), .B1(G134), .B2(new_n378), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G131), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n237), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n437), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n435), .B1(new_n436), .B2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n245), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n444), .B1(new_n437), .B2(new_n397), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n440), .B1(new_n389), .B2(new_n390), .ZN(new_n446));
  NOR3_X1   g260(.A1(new_n445), .A2(KEYINPUT30), .A3(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n195), .B1(new_n443), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(G210), .ZN(new_n449));
  NOR3_X1   g263(.A1(new_n449), .A2(G237), .A3(G953), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n450), .B(KEYINPUT27), .ZN(new_n451));
  XNOR2_X1  g265(.A(KEYINPUT26), .B(G101), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n451), .B(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n446), .B1(new_n409), .B2(new_n245), .ZN(new_n455));
  INV_X1    g269(.A(new_n195), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n448), .A2(new_n454), .A3(new_n457), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(KEYINPUT31), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n195), .B1(new_n445), .B2(new_n446), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NOR3_X1   g275(.A1(new_n445), .A2(new_n195), .A3(new_n446), .ZN(new_n462));
  OAI21_X1  g276(.A(KEYINPUT28), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT28), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n457), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n454), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n459), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT68), .ZN(new_n468));
  OAI21_X1  g282(.A(KEYINPUT30), .B1(new_n445), .B2(new_n446), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n442), .B(new_n435), .C1(new_n444), .C2(new_n392), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n462), .B1(new_n471), .B2(new_n195), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n468), .B1(new_n472), .B2(new_n454), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n456), .B1(new_n469), .B2(new_n470), .ZN(new_n474));
  NOR4_X1   g288(.A1(new_n474), .A2(KEYINPUT68), .A3(new_n453), .A4(new_n462), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT31), .ZN(new_n476));
  NOR3_X1   g290(.A1(new_n473), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT69), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n467), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n458), .A2(KEYINPUT68), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n472), .A2(new_n468), .A3(new_n454), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n480), .A2(new_n478), .A3(KEYINPUT31), .A4(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n434), .B1(new_n479), .B2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(G472), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n480), .A2(KEYINPUT31), .A3(new_n481), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(KEYINPUT69), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n487), .A2(KEYINPUT70), .A3(new_n482), .A4(new_n467), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n484), .A2(new_n485), .A3(new_n298), .A4(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT32), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n488), .A2(new_n298), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n492), .A2(KEYINPUT32), .A3(new_n485), .A4(new_n484), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n463), .A2(new_n454), .A3(new_n465), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT29), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n453), .B1(new_n474), .B2(new_n462), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT71), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n464), .B1(new_n457), .B2(new_n460), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n462), .A2(KEYINPUT28), .ZN(new_n501));
  NOR4_X1   g315(.A1(new_n500), .A2(new_n501), .A3(new_n495), .A4(new_n453), .ZN(new_n502));
  AOI21_X1  g316(.A(G902), .B1(new_n502), .B2(KEYINPUT72), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT72), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n504), .B1(new_n494), .B2(new_n495), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n494), .A2(KEYINPUT71), .A3(new_n495), .A4(new_n496), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n499), .A2(new_n503), .A3(new_n505), .A4(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(G472), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT73), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n508), .B(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n491), .A2(new_n493), .A3(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT23), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n512), .B1(new_n213), .B2(G128), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n231), .A2(KEYINPUT23), .A3(G119), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n513), .B(new_n514), .C1(G119), .C2(new_n231), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n515), .B(KEYINPUT75), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(G110), .ZN(new_n517));
  XOR2_X1   g331(.A(new_n517), .B(KEYINPUT76), .Z(new_n518));
  XNOR2_X1  g332(.A(G119), .B(G128), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n519), .B(KEYINPUT74), .ZN(new_n520));
  XNOR2_X1  g334(.A(KEYINPUT24), .B(G110), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n334), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n518), .A2(new_n523), .ZN(new_n524));
  OAI22_X1  g338(.A1(new_n520), .A2(new_n522), .B1(G110), .B2(new_n515), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n352), .A2(new_n323), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  XOR2_X1   g341(.A(KEYINPUT22), .B(G137), .Z(new_n528));
  NOR3_X1   g342(.A1(new_n366), .A2(new_n308), .A3(G953), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n528), .B(new_n529), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n527), .B(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(G217), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n532), .B1(G234), .B2(new_n298), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n533), .A2(G902), .ZN(new_n534));
  XOR2_X1   g348(.A(new_n534), .B(KEYINPUT79), .Z(new_n535));
  NAND2_X1  g349(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n531), .A2(new_n298), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT25), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n531), .A2(new_n538), .A3(new_n298), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n533), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n536), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n511), .A2(KEYINPUT80), .A3(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(KEYINPUT80), .B1(new_n511), .B2(new_n543), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n433), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n547), .B(new_n202), .ZN(G3));
  OR2_X1    g362(.A1(new_n271), .A2(new_n273), .ZN(new_n549));
  OR2_X1    g363(.A1(new_n549), .A2(new_n314), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n363), .A2(new_n364), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT94), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n297), .A2(new_n553), .ZN(new_n554));
  XOR2_X1   g368(.A(new_n554), .B(KEYINPUT33), .Z(new_n555));
  NAND3_X1  g369(.A1(new_n555), .A2(G478), .A3(new_n298), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n556), .B1(G478), .B2(new_n299), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n552), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n550), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n484), .A2(new_n298), .A3(new_n488), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(G472), .ZN(new_n561));
  AND4_X1   g375(.A1(new_n431), .A2(new_n561), .A3(new_n543), .A4(new_n489), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  XOR2_X1   g377(.A(KEYINPUT34), .B(G104), .Z(new_n564));
  XNOR2_X1  g378(.A(new_n563), .B(new_n564), .ZN(G6));
  INV_X1    g379(.A(new_n304), .ZN(new_n566));
  NOR3_X1   g380(.A1(new_n550), .A2(new_n361), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n562), .ZN(new_n568));
  XOR2_X1   g382(.A(KEYINPUT35), .B(G107), .Z(new_n569));
  XNOR2_X1  g383(.A(new_n568), .B(new_n569), .ZN(G9));
  INV_X1    g384(.A(KEYINPUT36), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n530), .A2(new_n571), .ZN(new_n572));
  XOR2_X1   g386(.A(new_n572), .B(KEYINPUT95), .Z(new_n573));
  XOR2_X1   g387(.A(new_n527), .B(new_n573), .Z(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n535), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n575), .B1(new_n539), .B2(new_n541), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n433), .A2(new_n489), .A3(new_n561), .A4(new_n576), .ZN(new_n577));
  XOR2_X1   g391(.A(KEYINPUT37), .B(G110), .Z(new_n578));
  XNOR2_X1  g392(.A(new_n577), .B(new_n578), .ZN(G12));
  NAND2_X1  g393(.A1(new_n274), .A2(new_n576), .ZN(new_n580));
  INV_X1    g394(.A(new_n361), .ZN(new_n581));
  INV_X1    g395(.A(G900), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n311), .B1(new_n582), .B2(new_n313), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n581), .A2(new_n304), .A3(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n511), .A2(new_n586), .A3(new_n431), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(G128), .ZN(G30));
  XNOR2_X1  g402(.A(new_n271), .B(KEYINPUT38), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n552), .A2(new_n304), .ZN(new_n590));
  NOR4_X1   g404(.A1(new_n589), .A2(new_n273), .A3(new_n576), .A4(new_n590), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n473), .A2(new_n475), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n454), .B1(new_n457), .B2(new_n460), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n298), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(G472), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n491), .A2(new_n493), .A3(new_n596), .ZN(new_n597));
  XOR2_X1   g411(.A(new_n583), .B(KEYINPUT39), .Z(new_n598));
  AOI21_X1  g412(.A(KEYINPUT40), .B1(new_n431), .B2(new_n598), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n431), .A2(KEYINPUT40), .A3(new_n598), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n591), .B(new_n597), .C1(new_n599), .C2(new_n600), .ZN(new_n601));
  XOR2_X1   g415(.A(new_n601), .B(KEYINPUT96), .Z(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(G143), .ZN(G45));
  NAND3_X1  g417(.A1(new_n552), .A2(new_n557), .A3(new_n584), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n580), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n511), .A2(new_n605), .A3(new_n431), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(G146), .ZN(G48));
  AND2_X1   g421(.A1(new_n511), .A2(new_n543), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n427), .A2(new_n298), .A3(new_n428), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(G469), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n430), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n611), .A2(new_n367), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n608), .A2(new_n559), .A3(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(KEYINPUT41), .B(G113), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G15));
  NAND3_X1  g429(.A1(new_n608), .A2(new_n567), .A3(new_n612), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(G116), .ZN(G18));
  AND4_X1   g431(.A1(new_n365), .A2(new_n274), .A3(new_n576), .A4(new_n612), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n511), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(KEYINPUT97), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT97), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n511), .A2(new_n618), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(KEYINPUT98), .B(G119), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G21));
  INV_X1    g439(.A(new_n612), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n550), .A2(new_n590), .A3(new_n626), .ZN(new_n627));
  AOI211_X1 g441(.A(G472), .B(G902), .C1(new_n467), .C2(new_n486), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n628), .B1(new_n560), .B2(G472), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n542), .A2(KEYINPUT99), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT99), .ZN(new_n631));
  OAI211_X1 g445(.A(new_n631), .B(new_n536), .C1(new_n539), .C2(new_n541), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(KEYINPUT100), .B1(new_n629), .B2(new_n633), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n629), .A2(KEYINPUT100), .A3(new_n633), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n627), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G122), .ZN(G24));
  NOR2_X1   g451(.A1(new_n549), .A2(new_n626), .ZN(new_n638));
  INV_X1    g452(.A(new_n604), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n638), .A2(new_n629), .A3(new_n576), .A4(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(G125), .ZN(G27));
  NAND2_X1  g455(.A1(new_n271), .A2(new_n272), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n423), .A2(KEYINPUT101), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT101), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n395), .A2(new_n422), .A3(new_n644), .A4(new_n415), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n417), .A2(G469), .A3(new_n643), .A4(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(G469), .A2(G902), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n430), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT102), .ZN(new_n649));
  INV_X1    g463(.A(new_n367), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n648), .A2(new_n650), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(KEYINPUT102), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n642), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n511), .A2(new_n543), .A3(new_n639), .A4(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT42), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AND3_X1   g471(.A1(new_n484), .A2(new_n298), .A3(new_n488), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT103), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n658), .A2(new_n659), .A3(KEYINPUT32), .A4(new_n485), .ZN(new_n660));
  OAI21_X1  g474(.A(KEYINPUT103), .B1(new_n489), .B2(new_n490), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n660), .A2(new_n510), .A3(new_n661), .A4(new_n491), .ZN(new_n662));
  AND3_X1   g476(.A1(new_n654), .A2(KEYINPUT42), .A3(new_n639), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n662), .A2(new_n663), .A3(new_n633), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n657), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G131), .ZN(G33));
  INV_X1    g480(.A(new_n585), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n511), .A2(new_n543), .A3(new_n667), .A4(new_n654), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G134), .ZN(G36));
  NAND2_X1  g483(.A1(new_n561), .A2(new_n489), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n551), .A2(new_n557), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n670), .A2(new_n673), .A3(new_n576), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n675));
  OAI211_X1 g489(.A(new_n272), .B(new_n271), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT105), .ZN(new_n677));
  OR2_X1    g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AOI22_X1  g492(.A1(new_n676), .A2(new_n677), .B1(new_n675), .B2(new_n674), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n680), .A2(KEYINPUT106), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n678), .A2(new_n679), .A3(KEYINPUT106), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT45), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n424), .A2(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n417), .A2(KEYINPUT45), .A3(new_n643), .A4(new_n645), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n685), .A2(G469), .A3(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n687), .A2(KEYINPUT46), .A3(new_n647), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(new_n430), .ZN(new_n689));
  AOI21_X1  g503(.A(KEYINPUT46), .B1(new_n687), .B2(new_n647), .ZN(new_n690));
  OAI211_X1 g504(.A(new_n650), .B(new_n598), .C1(new_n689), .C2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(KEYINPUT104), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n683), .A2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n682), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G137), .ZN(G39));
  OAI21_X1  g510(.A(new_n650), .B1(new_n689), .B2(new_n690), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(KEYINPUT47), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n639), .A2(new_n272), .A3(new_n271), .A4(new_n542), .ZN(new_n699));
  OR3_X1    g513(.A1(new_n698), .A2(new_n511), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G140), .ZN(G42));
  NAND3_X1  g515(.A1(new_n633), .A2(new_n272), .A3(new_n650), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n702), .A2(new_n671), .ZN(new_n703));
  INV_X1    g517(.A(new_n597), .ZN(new_n704));
  XOR2_X1   g518(.A(new_n611), .B(KEYINPUT49), .Z(new_n705));
  NAND4_X1  g519(.A1(new_n703), .A2(new_n704), .A3(new_n589), .A4(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT107), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n511), .A2(new_n543), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT80), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n432), .B1(new_n710), .B2(new_n544), .ZN(new_n711));
  INV_X1    g525(.A(new_n563), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n707), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n547), .A2(new_n563), .A3(KEYINPUT107), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n623), .A2(new_n613), .A3(new_n616), .A4(new_n636), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n629), .A2(new_n654), .A3(new_n576), .A4(new_n639), .ZN(new_n717));
  XOR2_X1   g531(.A(new_n304), .B(KEYINPUT108), .Z(new_n718));
  NAND4_X1  g532(.A1(new_n718), .A2(new_n576), .A3(new_n581), .A4(new_n584), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n719), .A2(new_n642), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n511), .A2(new_n431), .A3(new_n720), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n668), .A2(new_n717), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n665), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n716), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n718), .A2(new_n552), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n550), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n562), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n577), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  AND3_X1   g544(.A1(new_n587), .A2(new_n606), .A3(new_n640), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n549), .A2(new_n590), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n576), .A2(new_n652), .A3(new_n583), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n597), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n731), .A2(KEYINPUT52), .A3(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n587), .A2(new_n606), .A3(new_n734), .A4(new_n640), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT52), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n715), .A2(new_n724), .A3(new_n730), .A4(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT53), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT110), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n729), .B1(new_n713), .B2(new_n714), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n736), .A2(KEYINPUT109), .A3(new_n737), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n736), .A2(KEYINPUT109), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n735), .A2(new_n738), .A3(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n744), .A2(new_n724), .A3(new_n745), .A4(new_n747), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n743), .B1(new_n748), .B2(new_n741), .ZN(new_n749));
  AND3_X1   g563(.A1(new_n715), .A2(new_n724), .A3(new_n730), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n747), .A2(new_n745), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n750), .A2(KEYINPUT110), .A3(KEYINPUT53), .A4(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n742), .B1(new_n749), .B2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT54), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n748), .A2(new_n741), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n756), .B1(new_n741), .B2(new_n740), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(KEYINPUT54), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n626), .A2(new_n642), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n673), .A2(new_n311), .A3(new_n760), .ZN(new_n761));
  XOR2_X1   g575(.A(new_n761), .B(KEYINPUT114), .Z(new_n762));
  AND2_X1   g576(.A1(new_n629), .A2(new_n576), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(KEYINPUT115), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n704), .A2(new_n311), .A3(new_n543), .A4(new_n760), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n766), .A2(new_n552), .A3(new_n557), .ZN(new_n767));
  OR2_X1    g581(.A1(new_n767), .A2(KEYINPUT116), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(KEYINPUT116), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n765), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n673), .A2(new_n311), .ZN(new_n771));
  INV_X1    g585(.A(new_n635), .ZN(new_n772));
  INV_X1    g586(.A(new_n634), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n771), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT112), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n612), .A2(new_n273), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n589), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n777), .B1(new_n775), .B2(new_n776), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n774), .A2(KEYINPUT50), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(KEYINPUT50), .B1(new_n774), .B2(new_n778), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n774), .A2(new_n272), .A3(new_n271), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n610), .A2(new_n367), .A3(new_n430), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n782), .B1(new_n698), .B2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT51), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n781), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n770), .A2(new_n786), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n662), .A2(new_n633), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n762), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(KEYINPUT48), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n307), .B1(new_n766), .B2(new_n558), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n791), .B1(new_n774), .B2(new_n638), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n787), .A2(new_n790), .A3(new_n792), .ZN(new_n793));
  OR3_X1    g607(.A1(new_n779), .A2(new_n780), .A3(KEYINPUT113), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n770), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g609(.A(KEYINPUT113), .B1(new_n779), .B2(new_n780), .ZN(new_n796));
  AOI21_X1  g610(.A(KEYINPUT117), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n770), .A2(KEYINPUT117), .A3(new_n796), .A4(new_n794), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n783), .B(KEYINPUT111), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n698), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n798), .B1(new_n782), .B2(new_n800), .ZN(new_n801));
  OR2_X1    g615(.A1(new_n797), .A2(new_n801), .ZN(new_n802));
  AOI211_X1 g616(.A(new_n759), .B(new_n793), .C1(new_n802), .C2(new_n785), .ZN(new_n803));
  NOR2_X1   g617(.A1(G952), .A2(G953), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n706), .B1(new_n803), .B2(new_n804), .ZN(G75));
  INV_X1    g619(.A(KEYINPUT56), .ZN(new_n806));
  INV_X1    g620(.A(new_n753), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(G902), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n806), .B1(new_n808), .B2(new_n449), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n225), .B(new_n249), .ZN(new_n810));
  XOR2_X1   g624(.A(KEYINPUT118), .B(KEYINPUT55), .Z(new_n811));
  XNOR2_X1  g625(.A(new_n810), .B(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n809), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n809), .A2(new_n813), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n247), .A2(G952), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(G51));
  NAND2_X1  g631(.A1(new_n807), .A2(KEYINPUT54), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n818), .A2(new_n755), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n647), .B(KEYINPUT57), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n427), .B(new_n428), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  OR2_X1    g635(.A1(new_n808), .A2(new_n687), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n816), .B1(new_n821), .B2(new_n822), .ZN(G54));
  NAND4_X1  g637(.A1(new_n807), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n824));
  INV_X1    g638(.A(new_n355), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n824), .A2(new_n825), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n826), .A2(new_n827), .A3(new_n816), .ZN(G60));
  NAND2_X1  g642(.A1(G478), .A2(G902), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(KEYINPUT59), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n555), .B1(new_n759), .B2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n816), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n555), .A2(new_n830), .ZN(new_n833));
  OAI211_X1 g647(.A(KEYINPUT119), .B(new_n832), .C1(new_n819), .C2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT119), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n833), .B1(new_n818), .B2(new_n755), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n835), .B1(new_n836), .B2(new_n816), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n831), .B1(new_n834), .B2(new_n837), .ZN(G63));
  INV_X1    g652(.A(KEYINPUT61), .ZN(new_n839));
  XNOR2_X1  g653(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n840), .B(KEYINPUT121), .ZN(new_n841));
  NAND2_X1  g655(.A1(G217), .A2(G902), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n841), .B(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n749), .A2(new_n752), .ZN(new_n845));
  INV_X1    g659(.A(new_n742), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n832), .B1(new_n847), .B2(new_n531), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT124), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT124), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n850), .B(new_n832), .C1(new_n847), .C2(new_n531), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT122), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n853), .B1(new_n847), .B2(new_n574), .ZN(new_n854));
  INV_X1    g668(.A(new_n574), .ZN(new_n855));
  NOR4_X1   g669(.A1(new_n753), .A2(KEYINPUT122), .A3(new_n855), .A4(new_n844), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n854), .A2(new_n856), .A3(KEYINPUT123), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n839), .B1(new_n852), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n839), .A2(KEYINPUT123), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n859), .B1(new_n848), .B2(new_n839), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n860), .B1(new_n856), .B2(new_n854), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n858), .A2(new_n861), .ZN(G66));
  NAND2_X1  g676(.A1(G224), .A2(G953), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n312), .A2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n716), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n744), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(KEYINPUT125), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n864), .B1(new_n867), .B2(new_n247), .ZN(new_n868));
  INV_X1    g682(.A(G898), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n225), .B1(new_n869), .B2(G953), .ZN(new_n870));
  XOR2_X1   g684(.A(new_n868), .B(new_n870), .Z(G69));
  NAND3_X1  g685(.A1(new_n788), .A2(new_n692), .A3(new_n732), .ZN(new_n872));
  AND4_X1   g686(.A1(new_n668), .A2(new_n700), .A3(new_n872), .A4(new_n731), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n695), .A2(new_n665), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(new_n247), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n471), .B(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n875), .B(new_n878), .C1(new_n582), .C2(new_n247), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n602), .A2(new_n731), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT62), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n602), .A2(KEYINPUT62), .A3(new_n731), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT126), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n431), .A2(new_n598), .ZN(new_n887));
  AOI211_X1 g701(.A(new_n887), .B(new_n642), .C1(new_n726), .C2(new_n558), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n888), .B1(new_n545), .B2(new_n546), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n700), .B(new_n889), .C1(new_n681), .C2(new_n693), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n885), .A2(new_n886), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n700), .A2(new_n889), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n892), .B1(new_n682), .B2(new_n694), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT126), .B1(new_n893), .B2(new_n884), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n247), .B1(new_n891), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(KEYINPUT127), .B1(new_n895), .B2(new_n877), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n886), .B1(new_n885), .B2(new_n890), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n893), .A2(KEYINPUT126), .A3(new_n884), .ZN(new_n898));
  AOI21_X1  g712(.A(G953), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT127), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n899), .A2(new_n900), .A3(new_n878), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n879), .B1(new_n896), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n247), .B1(G227), .B2(G900), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n903), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n905), .B(new_n879), .C1(new_n896), .C2(new_n901), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n904), .A2(new_n906), .ZN(G72));
  NAND3_X1  g721(.A1(new_n897), .A2(new_n867), .A3(new_n898), .ZN(new_n908));
  NAND2_X1  g722(.A1(G472), .A2(G902), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n909), .B(KEYINPUT63), .Z(new_n910));
  AOI211_X1 g724(.A(new_n453), .B(new_n472), .C1(new_n908), .C2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(new_n910), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n912), .B1(new_n874), .B2(new_n867), .ZN(new_n913));
  NOR4_X1   g727(.A1(new_n913), .A2(new_n454), .A3(new_n462), .A4(new_n474), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n912), .B1(new_n592), .B2(new_n496), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n757), .A2(new_n915), .ZN(new_n916));
  NOR4_X1   g730(.A1(new_n911), .A2(new_n914), .A3(new_n816), .A4(new_n916), .ZN(G57));
endmodule


