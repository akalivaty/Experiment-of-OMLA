

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X2 U552 ( .A1(n521), .A2(G2104), .ZN(n522) );
  OR2_X1 U553 ( .A1(n817), .A2(n816), .ZN(n818) );
  AND2_X1 U554 ( .A1(n744), .A2(n743), .ZN(n745) );
  INV_X1 U555 ( .A(n737), .ZN(n711) );
  NOR2_X1 U556 ( .A1(n729), .A2(n727), .ZN(n717) );
  NOR2_X1 U557 ( .A1(G2105), .A2(G2104), .ZN(n524) );
  AND2_X1 U558 ( .A1(n530), .A2(n529), .ZN(G164) );
  AND2_X1 U559 ( .A1(G138), .A2(n881), .ZN(n519) );
  XOR2_X1 U560 ( .A(n720), .B(n719), .Z(n520) );
  INV_X1 U561 ( .A(KEYINPUT99), .ZN(n716) );
  NOR2_X1 U562 ( .A1(n726), .A2(n725), .ZN(n732) );
  INV_X1 U563 ( .A(KEYINPUT91), .ZN(n682) );
  XNOR2_X1 U564 ( .A(n683), .B(n682), .ZN(n792) );
  INV_X1 U565 ( .A(G2105), .ZN(n521) );
  XNOR2_X2 U566 ( .A(n522), .B(KEYINPUT66), .ZN(n883) );
  NAND2_X1 U567 ( .A1(n883), .A2(G102), .ZN(n523) );
  XOR2_X1 U568 ( .A(KEYINPUT90), .B(n523), .Z(n525) );
  XOR2_X2 U569 ( .A(KEYINPUT17), .B(n524), .Z(n881) );
  NOR2_X1 U570 ( .A1(n525), .A2(n519), .ZN(n530) );
  NOR2_X2 U571 ( .A1(G2104), .A2(n521), .ZN(n877) );
  NAND2_X1 U572 ( .A1(G126), .A2(n877), .ZN(n527) );
  AND2_X1 U573 ( .A1(G2105), .A2(G2104), .ZN(n878) );
  NAND2_X1 U574 ( .A1(G114), .A2(n878), .ZN(n526) );
  NAND2_X1 U575 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U576 ( .A(n528), .B(KEYINPUT89), .ZN(n529) );
  NOR2_X1 U577 ( .A1(G651), .A2(G543), .ZN(n639) );
  NAND2_X1 U578 ( .A1(G88), .A2(n639), .ZN(n533) );
  INV_X1 U579 ( .A(G651), .ZN(n535) );
  XOR2_X1 U580 ( .A(KEYINPUT0), .B(G543), .Z(n636) );
  OR2_X1 U581 ( .A1(n535), .A2(n636), .ZN(n531) );
  XOR2_X1 U582 ( .A(KEYINPUT68), .B(n531), .Z(n640) );
  NAND2_X1 U583 ( .A1(G75), .A2(n640), .ZN(n532) );
  NAND2_X1 U584 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U585 ( .A(KEYINPUT83), .B(n534), .ZN(n543) );
  NOR2_X1 U586 ( .A1(G543), .A2(n535), .ZN(n536) );
  XOR2_X1 U587 ( .A(KEYINPUT1), .B(n536), .Z(n643) );
  NAND2_X1 U588 ( .A1(G62), .A2(n643), .ZN(n537) );
  XNOR2_X1 U589 ( .A(n537), .B(KEYINPUT81), .ZN(n541) );
  NOR2_X1 U590 ( .A1(G651), .A2(n636), .ZN(n538) );
  XOR2_X1 U591 ( .A(KEYINPUT65), .B(n538), .Z(n644) );
  NAND2_X1 U592 ( .A1(G50), .A2(n644), .ZN(n539) );
  XOR2_X1 U593 ( .A(KEYINPUT82), .B(n539), .Z(n540) );
  NOR2_X1 U594 ( .A1(n541), .A2(n540), .ZN(n542) );
  NAND2_X1 U595 ( .A1(n543), .A2(n542), .ZN(G303) );
  INV_X1 U596 ( .A(G303), .ZN(G166) );
  NAND2_X1 U597 ( .A1(n883), .A2(G101), .ZN(n544) );
  XNOR2_X1 U598 ( .A(n544), .B(KEYINPUT23), .ZN(n545) );
  XNOR2_X1 U599 ( .A(n545), .B(KEYINPUT67), .ZN(n680) );
  NAND2_X1 U600 ( .A1(G137), .A2(n881), .ZN(n549) );
  NAND2_X1 U601 ( .A1(G125), .A2(n877), .ZN(n547) );
  NAND2_X1 U602 ( .A1(G113), .A2(n878), .ZN(n546) );
  AND2_X1 U603 ( .A1(n547), .A2(n546), .ZN(n548) );
  AND2_X1 U604 ( .A1(n549), .A2(n548), .ZN(n679) );
  AND2_X1 U605 ( .A1(n680), .A2(n679), .ZN(G160) );
  NAND2_X1 U606 ( .A1(n644), .A2(G52), .ZN(n551) );
  NAND2_X1 U607 ( .A1(n643), .A2(G64), .ZN(n550) );
  NAND2_X1 U608 ( .A1(n551), .A2(n550), .ZN(n556) );
  NAND2_X1 U609 ( .A1(G77), .A2(n640), .ZN(n553) );
  NAND2_X1 U610 ( .A1(n639), .A2(G90), .ZN(n552) );
  NAND2_X1 U611 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U612 ( .A(KEYINPUT9), .B(n554), .Z(n555) );
  NOR2_X1 U613 ( .A1(n556), .A2(n555), .ZN(G171) );
  INV_X1 U614 ( .A(G57), .ZN(G237) );
  AND2_X1 U615 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U616 ( .A1(G65), .A2(n643), .ZN(n558) );
  NAND2_X1 U617 ( .A1(G53), .A2(n644), .ZN(n557) );
  NAND2_X1 U618 ( .A1(n558), .A2(n557), .ZN(n562) );
  NAND2_X1 U619 ( .A1(G91), .A2(n639), .ZN(n560) );
  NAND2_X1 U620 ( .A1(G78), .A2(n640), .ZN(n559) );
  NAND2_X1 U621 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U622 ( .A1(n562), .A2(n561), .ZN(n920) );
  INV_X1 U623 ( .A(n920), .ZN(G299) );
  INV_X1 U624 ( .A(G108), .ZN(G238) );
  INV_X1 U625 ( .A(G120), .ZN(G236) );
  INV_X1 U626 ( .A(G132), .ZN(G219) );
  INV_X1 U627 ( .A(G82), .ZN(G220) );
  NAND2_X1 U628 ( .A1(n639), .A2(G89), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(KEYINPUT4), .ZN(n565) );
  NAND2_X1 U630 ( .A1(G76), .A2(n640), .ZN(n564) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(KEYINPUT5), .ZN(n572) );
  XNOR2_X1 U633 ( .A(KEYINPUT6), .B(KEYINPUT75), .ZN(n570) );
  NAND2_X1 U634 ( .A1(G63), .A2(n643), .ZN(n568) );
  NAND2_X1 U635 ( .A1(G51), .A2(n644), .ZN(n567) );
  NAND2_X1 U636 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(n571) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(KEYINPUT7), .B(n573), .ZN(G168) );
  XOR2_X1 U640 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U641 ( .A1(G7), .A2(G661), .ZN(n574) );
  XNOR2_X1 U642 ( .A(n574), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U643 ( .A(G223), .B(KEYINPUT70), .Z(n831) );
  NAND2_X1 U644 ( .A1(n831), .A2(G567), .ZN(n575) );
  XNOR2_X1 U645 ( .A(n575), .B(KEYINPUT71), .ZN(n576) );
  XNOR2_X1 U646 ( .A(KEYINPUT11), .B(n576), .ZN(G234) );
  NAND2_X1 U647 ( .A1(n639), .A2(G81), .ZN(n577) );
  XNOR2_X1 U648 ( .A(n577), .B(KEYINPUT12), .ZN(n579) );
  NAND2_X1 U649 ( .A1(G68), .A2(n640), .ZN(n578) );
  NAND2_X1 U650 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U651 ( .A(KEYINPUT13), .B(n580), .ZN(n586) );
  NAND2_X1 U652 ( .A1(G56), .A2(n643), .ZN(n581) );
  XOR2_X1 U653 ( .A(KEYINPUT14), .B(n581), .Z(n584) );
  NAND2_X1 U654 ( .A1(n644), .A2(G43), .ZN(n582) );
  XOR2_X1 U655 ( .A(KEYINPUT72), .B(n582), .Z(n583) );
  NOR2_X1 U656 ( .A1(n584), .A2(n583), .ZN(n585) );
  NAND2_X1 U657 ( .A1(n586), .A2(n585), .ZN(n914) );
  INV_X1 U658 ( .A(G860), .ZN(n600) );
  OR2_X1 U659 ( .A1(n914), .A2(n600), .ZN(G153) );
  INV_X1 U660 ( .A(G868), .ZN(n659) );
  NOR2_X1 U661 ( .A1(n659), .A2(G171), .ZN(n587) );
  XNOR2_X1 U662 ( .A(n587), .B(KEYINPUT73), .ZN(n596) );
  NAND2_X1 U663 ( .A1(G92), .A2(n639), .ZN(n589) );
  NAND2_X1 U664 ( .A1(G79), .A2(n640), .ZN(n588) );
  NAND2_X1 U665 ( .A1(n589), .A2(n588), .ZN(n593) );
  NAND2_X1 U666 ( .A1(G66), .A2(n643), .ZN(n591) );
  NAND2_X1 U667 ( .A1(G54), .A2(n644), .ZN(n590) );
  NAND2_X1 U668 ( .A1(n591), .A2(n590), .ZN(n592) );
  NOR2_X1 U669 ( .A1(n593), .A2(n592), .ZN(n594) );
  XOR2_X1 U670 ( .A(KEYINPUT15), .B(n594), .Z(n915) );
  OR2_X1 U671 ( .A1(G868), .A2(n915), .ZN(n595) );
  NAND2_X1 U672 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U673 ( .A(KEYINPUT74), .B(n597), .ZN(G284) );
  NOR2_X1 U674 ( .A1(G286), .A2(n659), .ZN(n599) );
  NOR2_X1 U675 ( .A1(G868), .A2(G299), .ZN(n598) );
  NOR2_X1 U676 ( .A1(n599), .A2(n598), .ZN(G297) );
  NAND2_X1 U677 ( .A1(n600), .A2(G559), .ZN(n601) );
  NAND2_X1 U678 ( .A1(n601), .A2(n915), .ZN(n602) );
  XNOR2_X1 U679 ( .A(n602), .B(KEYINPUT76), .ZN(n603) );
  XNOR2_X1 U680 ( .A(KEYINPUT16), .B(n603), .ZN(G148) );
  NOR2_X1 U681 ( .A1(G868), .A2(n914), .ZN(n606) );
  NAND2_X1 U682 ( .A1(G868), .A2(n915), .ZN(n604) );
  NOR2_X1 U683 ( .A1(G559), .A2(n604), .ZN(n605) );
  NOR2_X1 U684 ( .A1(n606), .A2(n605), .ZN(G282) );
  NAND2_X1 U685 ( .A1(G123), .A2(n877), .ZN(n607) );
  XNOR2_X1 U686 ( .A(n607), .B(KEYINPUT18), .ZN(n610) );
  NAND2_X1 U687 ( .A1(G111), .A2(n878), .ZN(n608) );
  XOR2_X1 U688 ( .A(KEYINPUT77), .B(n608), .Z(n609) );
  NAND2_X1 U689 ( .A1(n610), .A2(n609), .ZN(n614) );
  NAND2_X1 U690 ( .A1(n881), .A2(G135), .ZN(n612) );
  NAND2_X1 U691 ( .A1(G99), .A2(n883), .ZN(n611) );
  NAND2_X1 U692 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U693 ( .A1(n614), .A2(n613), .ZN(n942) );
  XNOR2_X1 U694 ( .A(G2096), .B(n942), .ZN(n616) );
  INV_X1 U695 ( .A(G2100), .ZN(n615) );
  NAND2_X1 U696 ( .A1(n616), .A2(n615), .ZN(G156) );
  NAND2_X1 U697 ( .A1(n640), .A2(G73), .ZN(n617) );
  XOR2_X1 U698 ( .A(KEYINPUT79), .B(n617), .Z(n618) );
  XNOR2_X1 U699 ( .A(n618), .B(KEYINPUT2), .ZN(n620) );
  NAND2_X1 U700 ( .A1(G86), .A2(n639), .ZN(n619) );
  NAND2_X1 U701 ( .A1(n620), .A2(n619), .ZN(n624) );
  NAND2_X1 U702 ( .A1(G61), .A2(n643), .ZN(n622) );
  NAND2_X1 U703 ( .A1(G48), .A2(n644), .ZN(n621) );
  NAND2_X1 U704 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U705 ( .A1(n624), .A2(n623), .ZN(n625) );
  XOR2_X1 U706 ( .A(KEYINPUT80), .B(n625), .Z(G305) );
  NAND2_X1 U707 ( .A1(G85), .A2(n639), .ZN(n627) );
  NAND2_X1 U708 ( .A1(G72), .A2(n640), .ZN(n626) );
  NAND2_X1 U709 ( .A1(n627), .A2(n626), .ZN(n630) );
  NAND2_X1 U710 ( .A1(G60), .A2(n643), .ZN(n628) );
  XNOR2_X1 U711 ( .A(KEYINPUT69), .B(n628), .ZN(n629) );
  NOR2_X1 U712 ( .A1(n630), .A2(n629), .ZN(n632) );
  NAND2_X1 U713 ( .A1(n644), .A2(G47), .ZN(n631) );
  NAND2_X1 U714 ( .A1(n632), .A2(n631), .ZN(G290) );
  NAND2_X1 U715 ( .A1(G49), .A2(n644), .ZN(n634) );
  NAND2_X1 U716 ( .A1(G74), .A2(G651), .ZN(n633) );
  NAND2_X1 U717 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U718 ( .A1(n643), .A2(n635), .ZN(n638) );
  NAND2_X1 U719 ( .A1(n636), .A2(G87), .ZN(n637) );
  NAND2_X1 U720 ( .A1(n638), .A2(n637), .ZN(G288) );
  XOR2_X1 U721 ( .A(KEYINPUT85), .B(KEYINPUT19), .Z(n651) );
  NAND2_X1 U722 ( .A1(G93), .A2(n639), .ZN(n642) );
  NAND2_X1 U723 ( .A1(G80), .A2(n640), .ZN(n641) );
  NAND2_X1 U724 ( .A1(n642), .A2(n641), .ZN(n648) );
  NAND2_X1 U725 ( .A1(G67), .A2(n643), .ZN(n646) );
  NAND2_X1 U726 ( .A1(G55), .A2(n644), .ZN(n645) );
  NAND2_X1 U727 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U728 ( .A1(n648), .A2(n647), .ZN(n649) );
  XOR2_X1 U729 ( .A(KEYINPUT78), .B(n649), .Z(n910) );
  XNOR2_X1 U730 ( .A(KEYINPUT84), .B(n910), .ZN(n650) );
  XNOR2_X1 U731 ( .A(n651), .B(n650), .ZN(n654) );
  XNOR2_X1 U732 ( .A(G305), .B(G299), .ZN(n652) );
  XNOR2_X1 U733 ( .A(n652), .B(G290), .ZN(n653) );
  XNOR2_X1 U734 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U735 ( .A(n655), .B(G288), .ZN(n656) );
  XNOR2_X1 U736 ( .A(G166), .B(n656), .ZN(n896) );
  NAND2_X1 U737 ( .A1(G559), .A2(n915), .ZN(n657) );
  XNOR2_X1 U738 ( .A(n657), .B(n914), .ZN(n908) );
  XNOR2_X1 U739 ( .A(n896), .B(n908), .ZN(n658) );
  NOR2_X1 U740 ( .A1(n659), .A2(n658), .ZN(n661) );
  NOR2_X1 U741 ( .A1(G868), .A2(n910), .ZN(n660) );
  NOR2_X1 U742 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U743 ( .A(KEYINPUT86), .B(n662), .ZN(G295) );
  NAND2_X1 U744 ( .A1(G2084), .A2(G2078), .ZN(n663) );
  XOR2_X1 U745 ( .A(KEYINPUT20), .B(n663), .Z(n664) );
  NAND2_X1 U746 ( .A1(G2090), .A2(n664), .ZN(n665) );
  XNOR2_X1 U747 ( .A(KEYINPUT21), .B(n665), .ZN(n666) );
  NAND2_X1 U748 ( .A1(n666), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U749 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U750 ( .A1(G220), .A2(G219), .ZN(n667) );
  XOR2_X1 U751 ( .A(KEYINPUT22), .B(n667), .Z(n668) );
  NOR2_X1 U752 ( .A1(G218), .A2(n668), .ZN(n669) );
  NAND2_X1 U753 ( .A1(G96), .A2(n669), .ZN(n911) );
  NAND2_X1 U754 ( .A1(G2106), .A2(n911), .ZN(n670) );
  XNOR2_X1 U755 ( .A(n670), .B(KEYINPUT87), .ZN(n674) );
  NOR2_X1 U756 ( .A1(G236), .A2(G238), .ZN(n671) );
  NAND2_X1 U757 ( .A1(G69), .A2(n671), .ZN(n672) );
  OR2_X1 U758 ( .A1(G237), .A2(n672), .ZN(n912) );
  AND2_X1 U759 ( .A1(G567), .A2(n912), .ZN(n673) );
  NOR2_X1 U760 ( .A1(n674), .A2(n673), .ZN(G319) );
  INV_X1 U761 ( .A(G319), .ZN(n676) );
  NAND2_X1 U762 ( .A1(G483), .A2(G661), .ZN(n675) );
  NOR2_X1 U763 ( .A1(n676), .A2(n675), .ZN(n834) );
  NAND2_X1 U764 ( .A1(n834), .A2(G36), .ZN(n677) );
  XNOR2_X1 U765 ( .A(KEYINPUT88), .B(n677), .ZN(G176) );
  INV_X1 U766 ( .A(G171), .ZN(G301) );
  NOR2_X1 U767 ( .A1(G1384), .A2(G164), .ZN(n678) );
  XNOR2_X1 U768 ( .A(n678), .B(KEYINPUT64), .ZN(n793) );
  AND2_X1 U769 ( .A1(n679), .A2(G40), .ZN(n681) );
  NAND2_X1 U770 ( .A1(n681), .A2(n680), .ZN(n683) );
  INV_X1 U771 ( .A(n792), .ZN(n684) );
  NAND2_X2 U772 ( .A1(n793), .A2(n684), .ZN(n737) );
  NAND2_X2 U773 ( .A1(G8), .A2(n737), .ZN(n806) );
  NOR2_X1 U774 ( .A1(G1976), .A2(G288), .ZN(n687) );
  NAND2_X1 U775 ( .A1(n687), .A2(KEYINPUT33), .ZN(n685) );
  NOR2_X1 U776 ( .A1(n806), .A2(n685), .ZN(n753) );
  NOR2_X1 U777 ( .A1(G1971), .A2(G303), .ZN(n686) );
  NOR2_X1 U778 ( .A1(n687), .A2(n686), .ZN(n924) );
  INV_X1 U779 ( .A(n924), .ZN(n748) );
  NOR2_X1 U780 ( .A1(G1966), .A2(n806), .ZN(n727) );
  AND2_X1 U781 ( .A1(n711), .A2(G1996), .ZN(n688) );
  XNOR2_X1 U782 ( .A(KEYINPUT26), .B(n688), .ZN(n690) );
  AND2_X1 U783 ( .A1(n737), .A2(G1341), .ZN(n689) );
  NOR2_X1 U784 ( .A1(n690), .A2(n689), .ZN(n692) );
  INV_X1 U785 ( .A(n914), .ZN(n691) );
  AND2_X1 U786 ( .A1(n692), .A2(n691), .ZN(n693) );
  OR2_X1 U787 ( .A1(n693), .A2(n915), .ZN(n699) );
  NAND2_X1 U788 ( .A1(n693), .A2(n915), .ZN(n697) );
  NAND2_X1 U789 ( .A1(G1348), .A2(n737), .ZN(n695) );
  NAND2_X1 U790 ( .A1(n711), .A2(G2067), .ZN(n694) );
  NAND2_X1 U791 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U792 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U793 ( .A1(n699), .A2(n698), .ZN(n705) );
  NAND2_X1 U794 ( .A1(G2072), .A2(n711), .ZN(n701) );
  XNOR2_X1 U795 ( .A(KEYINPUT98), .B(KEYINPUT27), .ZN(n700) );
  XNOR2_X1 U796 ( .A(n701), .B(n700), .ZN(n703) );
  INV_X1 U797 ( .A(G1956), .ZN(n988) );
  NOR2_X1 U798 ( .A1(n711), .A2(n988), .ZN(n702) );
  NOR2_X1 U799 ( .A1(n703), .A2(n702), .ZN(n706) );
  NAND2_X1 U800 ( .A1(n706), .A2(n920), .ZN(n704) );
  NAND2_X1 U801 ( .A1(n705), .A2(n704), .ZN(n709) );
  NOR2_X1 U802 ( .A1(n706), .A2(n920), .ZN(n707) );
  XOR2_X1 U803 ( .A(n707), .B(KEYINPUT28), .Z(n708) );
  NAND2_X1 U804 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U805 ( .A(n710), .B(KEYINPUT29), .ZN(n715) );
  XOR2_X1 U806 ( .A(KEYINPUT25), .B(G2078), .Z(n972) );
  NOR2_X1 U807 ( .A1(n972), .A2(n737), .ZN(n713) );
  NOR2_X1 U808 ( .A1(n711), .A2(G1961), .ZN(n712) );
  NOR2_X1 U809 ( .A1(n713), .A2(n712), .ZN(n721) );
  NOR2_X1 U810 ( .A1(G301), .A2(n721), .ZN(n714) );
  NOR2_X1 U811 ( .A1(n715), .A2(n714), .ZN(n726) );
  NOR2_X1 U812 ( .A1(G2084), .A2(n737), .ZN(n729) );
  XNOR2_X1 U813 ( .A(n717), .B(n716), .ZN(n718) );
  NAND2_X1 U814 ( .A1(n718), .A2(G8), .ZN(n720) );
  XOR2_X1 U815 ( .A(KEYINPUT100), .B(KEYINPUT30), .Z(n719) );
  NOR2_X1 U816 ( .A1(G168), .A2(n520), .ZN(n723) );
  AND2_X1 U817 ( .A1(G301), .A2(n721), .ZN(n722) );
  NOR2_X1 U818 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U819 ( .A(n724), .B(KEYINPUT31), .ZN(n725) );
  NOR2_X1 U820 ( .A1(n727), .A2(n732), .ZN(n728) );
  XNOR2_X1 U821 ( .A(n728), .B(KEYINPUT101), .ZN(n731) );
  AND2_X1 U822 ( .A1(G8), .A2(n729), .ZN(n730) );
  NOR2_X1 U823 ( .A1(n731), .A2(n730), .ZN(n747) );
  INV_X1 U824 ( .A(n732), .ZN(n734) );
  AND2_X1 U825 ( .A1(G286), .A2(G8), .ZN(n733) );
  NAND2_X1 U826 ( .A1(n734), .A2(n733), .ZN(n744) );
  INV_X1 U827 ( .A(G8), .ZN(n742) );
  NOR2_X1 U828 ( .A1(G1971), .A2(n806), .ZN(n735) );
  XNOR2_X1 U829 ( .A(n735), .B(KEYINPUT102), .ZN(n736) );
  NOR2_X1 U830 ( .A1(G166), .A2(n736), .ZN(n740) );
  NOR2_X1 U831 ( .A1(G2090), .A2(n737), .ZN(n738) );
  XNOR2_X1 U832 ( .A(n738), .B(KEYINPUT103), .ZN(n739) );
  NAND2_X1 U833 ( .A1(n740), .A2(n739), .ZN(n741) );
  OR2_X1 U834 ( .A1(n742), .A2(n741), .ZN(n743) );
  XOR2_X1 U835 ( .A(KEYINPUT32), .B(n745), .Z(n746) );
  NOR2_X1 U836 ( .A1(n747), .A2(n746), .ZN(n809) );
  OR2_X1 U837 ( .A1(n748), .A2(n809), .ZN(n749) );
  NAND2_X1 U838 ( .A1(G1976), .A2(G288), .ZN(n923) );
  NAND2_X1 U839 ( .A1(n749), .A2(n923), .ZN(n750) );
  NOR2_X1 U840 ( .A1(n806), .A2(n750), .ZN(n751) );
  NOR2_X1 U841 ( .A1(KEYINPUT33), .A2(n751), .ZN(n752) );
  NOR2_X1 U842 ( .A1(n753), .A2(n752), .ZN(n801) );
  XOR2_X1 U843 ( .A(G305), .B(G1981), .Z(n930) );
  NAND2_X1 U844 ( .A1(n881), .A2(G140), .ZN(n755) );
  NAND2_X1 U845 ( .A1(G104), .A2(n883), .ZN(n754) );
  NAND2_X1 U846 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U847 ( .A(KEYINPUT34), .B(n756), .ZN(n762) );
  NAND2_X1 U848 ( .A1(n878), .A2(G116), .ZN(n757) );
  XNOR2_X1 U849 ( .A(n757), .B(KEYINPUT92), .ZN(n759) );
  NAND2_X1 U850 ( .A1(G128), .A2(n877), .ZN(n758) );
  NAND2_X1 U851 ( .A1(n759), .A2(n758), .ZN(n760) );
  XOR2_X1 U852 ( .A(n760), .B(KEYINPUT35), .Z(n761) );
  NOR2_X1 U853 ( .A1(n762), .A2(n761), .ZN(n763) );
  XOR2_X1 U854 ( .A(KEYINPUT36), .B(n763), .Z(n764) );
  XOR2_X1 U855 ( .A(KEYINPUT93), .B(n764), .Z(n893) );
  XOR2_X1 U856 ( .A(G2067), .B(KEYINPUT37), .Z(n765) );
  NOR2_X1 U857 ( .A1(n893), .A2(n765), .ZN(n958) );
  AND2_X1 U858 ( .A1(n893), .A2(n765), .ZN(n962) );
  NAND2_X1 U859 ( .A1(n883), .A2(G105), .ZN(n766) );
  XNOR2_X1 U860 ( .A(n766), .B(KEYINPUT38), .ZN(n773) );
  NAND2_X1 U861 ( .A1(G129), .A2(n877), .ZN(n768) );
  NAND2_X1 U862 ( .A1(G141), .A2(n881), .ZN(n767) );
  NAND2_X1 U863 ( .A1(n768), .A2(n767), .ZN(n771) );
  NAND2_X1 U864 ( .A1(n878), .A2(G117), .ZN(n769) );
  XOR2_X1 U865 ( .A(KEYINPUT96), .B(n769), .Z(n770) );
  NOR2_X1 U866 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U867 ( .A1(n773), .A2(n772), .ZN(n860) );
  NOR2_X1 U868 ( .A1(G1996), .A2(n860), .ZN(n955) );
  NAND2_X1 U869 ( .A1(n881), .A2(G131), .ZN(n775) );
  NAND2_X1 U870 ( .A1(G95), .A2(n883), .ZN(n774) );
  NAND2_X1 U871 ( .A1(n775), .A2(n774), .ZN(n778) );
  NAND2_X1 U872 ( .A1(n877), .A2(G119), .ZN(n776) );
  XOR2_X1 U873 ( .A(KEYINPUT94), .B(n776), .Z(n777) );
  NOR2_X1 U874 ( .A1(n778), .A2(n777), .ZN(n780) );
  NAND2_X1 U875 ( .A1(n878), .A2(G107), .ZN(n779) );
  NAND2_X1 U876 ( .A1(n780), .A2(n779), .ZN(n861) );
  NAND2_X1 U877 ( .A1(G1991), .A2(n861), .ZN(n781) );
  XOR2_X1 U878 ( .A(KEYINPUT95), .B(n781), .Z(n783) );
  NAND2_X1 U879 ( .A1(G1996), .A2(n860), .ZN(n782) );
  NAND2_X1 U880 ( .A1(n783), .A2(n782), .ZN(n943) );
  NOR2_X1 U881 ( .A1(G1986), .A2(G290), .ZN(n784) );
  NOR2_X1 U882 ( .A1(G1991), .A2(n861), .ZN(n944) );
  NOR2_X1 U883 ( .A1(n784), .A2(n944), .ZN(n785) );
  NOR2_X1 U884 ( .A1(n943), .A2(n785), .ZN(n786) );
  NOR2_X1 U885 ( .A1(n955), .A2(n786), .ZN(n787) );
  XOR2_X1 U886 ( .A(KEYINPUT39), .B(n787), .Z(n788) );
  NOR2_X1 U887 ( .A1(n962), .A2(n788), .ZN(n789) );
  XNOR2_X1 U888 ( .A(n789), .B(KEYINPUT104), .ZN(n790) );
  NOR2_X1 U889 ( .A1(n958), .A2(n790), .ZN(n791) );
  XNOR2_X1 U890 ( .A(KEYINPUT105), .B(n791), .ZN(n794) );
  NOR2_X1 U891 ( .A1(n793), .A2(n792), .ZN(n796) );
  NAND2_X1 U892 ( .A1(n794), .A2(n796), .ZN(n814) );
  INV_X1 U893 ( .A(n814), .ZN(n799) );
  XOR2_X1 U894 ( .A(G1986), .B(G290), .Z(n935) );
  NOR2_X1 U895 ( .A1(n962), .A2(n943), .ZN(n795) );
  NAND2_X1 U896 ( .A1(n935), .A2(n795), .ZN(n797) );
  NAND2_X1 U897 ( .A1(n797), .A2(n796), .ZN(n798) );
  OR2_X1 U898 ( .A1(n799), .A2(n798), .ZN(n802) );
  AND2_X1 U899 ( .A1(n930), .A2(n802), .ZN(n800) );
  NAND2_X1 U900 ( .A1(n801), .A2(n800), .ZN(n819) );
  INV_X1 U901 ( .A(n802), .ZN(n817) );
  NOR2_X1 U902 ( .A1(G305), .A2(G1981), .ZN(n803) );
  XNOR2_X1 U903 ( .A(n803), .B(KEYINPUT24), .ZN(n804) );
  XNOR2_X1 U904 ( .A(n804), .B(KEYINPUT97), .ZN(n805) );
  NOR2_X1 U905 ( .A1(n805), .A2(n806), .ZN(n813) );
  INV_X1 U906 ( .A(n806), .ZN(n811) );
  NAND2_X1 U907 ( .A1(G166), .A2(G8), .ZN(n807) );
  NOR2_X1 U908 ( .A1(G2090), .A2(n807), .ZN(n808) );
  NOR2_X1 U909 ( .A1(n809), .A2(n808), .ZN(n810) );
  NOR2_X1 U910 ( .A1(n811), .A2(n810), .ZN(n812) );
  NOR2_X1 U911 ( .A1(n813), .A2(n812), .ZN(n815) );
  AND2_X1 U912 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U913 ( .A1(n819), .A2(n818), .ZN(n820) );
  XNOR2_X1 U914 ( .A(KEYINPUT40), .B(n820), .ZN(G329) );
  XNOR2_X1 U915 ( .A(G2454), .B(G2435), .ZN(n829) );
  XNOR2_X1 U916 ( .A(KEYINPUT106), .B(G2427), .ZN(n827) );
  XOR2_X1 U917 ( .A(G2430), .B(G2446), .Z(n822) );
  XNOR2_X1 U918 ( .A(G2443), .B(G2451), .ZN(n821) );
  XNOR2_X1 U919 ( .A(n822), .B(n821), .ZN(n823) );
  XOR2_X1 U920 ( .A(n823), .B(G2438), .Z(n825) );
  XNOR2_X1 U921 ( .A(G1348), .B(G1341), .ZN(n824) );
  XNOR2_X1 U922 ( .A(n825), .B(n824), .ZN(n826) );
  XNOR2_X1 U923 ( .A(n827), .B(n826), .ZN(n828) );
  XNOR2_X1 U924 ( .A(n829), .B(n828), .ZN(n830) );
  NAND2_X1 U925 ( .A1(n830), .A2(G14), .ZN(n902) );
  XNOR2_X1 U926 ( .A(KEYINPUT107), .B(n902), .ZN(G401) );
  NAND2_X1 U927 ( .A1(G2106), .A2(n831), .ZN(G217) );
  AND2_X1 U928 ( .A1(G15), .A2(G2), .ZN(n832) );
  NAND2_X1 U929 ( .A1(G661), .A2(n832), .ZN(G259) );
  NAND2_X1 U930 ( .A1(G3), .A2(G1), .ZN(n833) );
  NAND2_X1 U931 ( .A1(n834), .A2(n833), .ZN(G188) );
  XOR2_X1 U932 ( .A(G2096), .B(KEYINPUT43), .Z(n836) );
  XNOR2_X1 U933 ( .A(G2072), .B(G2678), .ZN(n835) );
  XNOR2_X1 U934 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U935 ( .A(n837), .B(KEYINPUT108), .Z(n839) );
  XNOR2_X1 U936 ( .A(G2067), .B(G2090), .ZN(n838) );
  XNOR2_X1 U937 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U938 ( .A(KEYINPUT42), .B(G2100), .Z(n841) );
  XNOR2_X1 U939 ( .A(G2084), .B(G2078), .ZN(n840) );
  XNOR2_X1 U940 ( .A(n841), .B(n840), .ZN(n842) );
  XNOR2_X1 U941 ( .A(n843), .B(n842), .ZN(G227) );
  XOR2_X1 U942 ( .A(G1986), .B(G1981), .Z(n845) );
  XNOR2_X1 U943 ( .A(G1966), .B(G1956), .ZN(n844) );
  XNOR2_X1 U944 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U945 ( .A(n846), .B(KEYINPUT41), .Z(n848) );
  XNOR2_X1 U946 ( .A(G1971), .B(G1976), .ZN(n847) );
  XNOR2_X1 U947 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U948 ( .A(G2474), .B(G1991), .Z(n850) );
  XNOR2_X1 U949 ( .A(G1961), .B(G1996), .ZN(n849) );
  XNOR2_X1 U950 ( .A(n850), .B(n849), .ZN(n851) );
  XNOR2_X1 U951 ( .A(n852), .B(n851), .ZN(G229) );
  NAND2_X1 U952 ( .A1(n877), .A2(G124), .ZN(n853) );
  XNOR2_X1 U953 ( .A(n853), .B(KEYINPUT44), .ZN(n855) );
  NAND2_X1 U954 ( .A1(G100), .A2(n883), .ZN(n854) );
  NAND2_X1 U955 ( .A1(n855), .A2(n854), .ZN(n859) );
  NAND2_X1 U956 ( .A1(G112), .A2(n878), .ZN(n857) );
  NAND2_X1 U957 ( .A1(G136), .A2(n881), .ZN(n856) );
  NAND2_X1 U958 ( .A1(n857), .A2(n856), .ZN(n858) );
  NOR2_X1 U959 ( .A1(n859), .A2(n858), .ZN(G162) );
  XNOR2_X1 U960 ( .A(G160), .B(n860), .ZN(n862) );
  XNOR2_X1 U961 ( .A(n862), .B(n861), .ZN(n863) );
  XNOR2_X1 U962 ( .A(G164), .B(n863), .ZN(n892) );
  XOR2_X1 U963 ( .A(KEYINPUT48), .B(KEYINPUT112), .Z(n865) );
  XNOR2_X1 U964 ( .A(KEYINPUT46), .B(KEYINPUT110), .ZN(n864) );
  XNOR2_X1 U965 ( .A(n865), .B(n864), .ZN(n866) );
  XOR2_X1 U966 ( .A(n866), .B(n942), .Z(n876) );
  NAND2_X1 U967 ( .A1(n881), .A2(G139), .ZN(n868) );
  NAND2_X1 U968 ( .A1(G103), .A2(n883), .ZN(n867) );
  NAND2_X1 U969 ( .A1(n868), .A2(n867), .ZN(n874) );
  NAND2_X1 U970 ( .A1(G127), .A2(n877), .ZN(n870) );
  NAND2_X1 U971 ( .A1(G115), .A2(n878), .ZN(n869) );
  NAND2_X1 U972 ( .A1(n870), .A2(n869), .ZN(n871) );
  XNOR2_X1 U973 ( .A(KEYINPUT111), .B(n871), .ZN(n872) );
  XNOR2_X1 U974 ( .A(KEYINPUT47), .B(n872), .ZN(n873) );
  NOR2_X1 U975 ( .A1(n874), .A2(n873), .ZN(n947) );
  XNOR2_X1 U976 ( .A(n947), .B(G162), .ZN(n875) );
  XNOR2_X1 U977 ( .A(n876), .B(n875), .ZN(n890) );
  NAND2_X1 U978 ( .A1(G130), .A2(n877), .ZN(n880) );
  NAND2_X1 U979 ( .A1(G118), .A2(n878), .ZN(n879) );
  NAND2_X1 U980 ( .A1(n880), .A2(n879), .ZN(n888) );
  NAND2_X1 U981 ( .A1(n881), .A2(G142), .ZN(n882) );
  XOR2_X1 U982 ( .A(KEYINPUT109), .B(n882), .Z(n885) );
  NAND2_X1 U983 ( .A1(G106), .A2(n883), .ZN(n884) );
  NAND2_X1 U984 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U985 ( .A(n886), .B(KEYINPUT45), .Z(n887) );
  NOR2_X1 U986 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U987 ( .A(n890), .B(n889), .Z(n891) );
  XNOR2_X1 U988 ( .A(n892), .B(n891), .ZN(n894) );
  XNOR2_X1 U989 ( .A(n894), .B(n893), .ZN(n895) );
  NOR2_X1 U990 ( .A1(G37), .A2(n895), .ZN(G395) );
  XOR2_X1 U991 ( .A(KEYINPUT113), .B(n896), .Z(n898) );
  XNOR2_X1 U992 ( .A(n915), .B(G286), .ZN(n897) );
  XNOR2_X1 U993 ( .A(n898), .B(n897), .ZN(n900) );
  XOR2_X1 U994 ( .A(n914), .B(G171), .Z(n899) );
  XNOR2_X1 U995 ( .A(n900), .B(n899), .ZN(n901) );
  NOR2_X1 U996 ( .A1(G37), .A2(n901), .ZN(G397) );
  NAND2_X1 U997 ( .A1(G319), .A2(n902), .ZN(n905) );
  NOR2_X1 U998 ( .A1(G227), .A2(G229), .ZN(n903) );
  XNOR2_X1 U999 ( .A(KEYINPUT49), .B(n903), .ZN(n904) );
  NOR2_X1 U1000 ( .A1(n905), .A2(n904), .ZN(n907) );
  NOR2_X1 U1001 ( .A1(G395), .A2(G397), .ZN(n906) );
  NAND2_X1 U1002 ( .A1(n907), .A2(n906), .ZN(G225) );
  XOR2_X1 U1003 ( .A(KEYINPUT114), .B(G225), .Z(G308) );
  NOR2_X1 U1005 ( .A1(G860), .A2(n908), .ZN(n909) );
  XOR2_X1 U1006 ( .A(n910), .B(n909), .Z(G145) );
  INV_X1 U1007 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1008 ( .A1(n912), .A2(n911), .ZN(G325) );
  INV_X1 U1009 ( .A(G325), .ZN(G261) );
  INV_X1 U1010 ( .A(G69), .ZN(G235) );
  XOR2_X1 U1011 ( .A(G16), .B(KEYINPUT56), .Z(n940) );
  XOR2_X1 U1012 ( .A(G1341), .B(KEYINPUT123), .Z(n913) );
  XNOR2_X1 U1013 ( .A(n914), .B(n913), .ZN(n938) );
  XNOR2_X1 U1014 ( .A(G171), .B(G1961), .ZN(n918) );
  XNOR2_X1 U1015 ( .A(G1348), .B(n915), .ZN(n916) );
  XNOR2_X1 U1016 ( .A(n916), .B(KEYINPUT120), .ZN(n917) );
  NAND2_X1 U1017 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1018 ( .A(n919), .B(KEYINPUT121), .ZN(n929) );
  XNOR2_X1 U1019 ( .A(n920), .B(G1956), .ZN(n922) );
  NAND2_X1 U1020 ( .A1(G1971), .A2(G303), .ZN(n921) );
  NAND2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(n926) );
  NAND2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n925) );
  NOR2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1024 ( .A(n927), .B(KEYINPUT122), .ZN(n928) );
  NAND2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n934) );
  XNOR2_X1 U1026 ( .A(G1966), .B(G168), .ZN(n931) );
  NAND2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1028 ( .A(KEYINPUT57), .B(n932), .Z(n933) );
  NOR2_X1 U1029 ( .A1(n934), .A2(n933), .ZN(n936) );
  NAND2_X1 U1030 ( .A1(n936), .A2(n935), .ZN(n937) );
  NOR2_X1 U1031 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1032 ( .A1(n940), .A2(n939), .ZN(n1025) );
  INV_X1 U1033 ( .A(KEYINPUT55), .ZN(n966) );
  XNOR2_X1 U1034 ( .A(KEYINPUT116), .B(KEYINPUT52), .ZN(n964) );
  XOR2_X1 U1035 ( .A(G2084), .B(G160), .Z(n941) );
  NOR2_X1 U1036 ( .A1(n942), .A2(n941), .ZN(n946) );
  NOR2_X1 U1037 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1038 ( .A1(n946), .A2(n945), .ZN(n953) );
  XNOR2_X1 U1039 ( .A(G2072), .B(n947), .ZN(n949) );
  XNOR2_X1 U1040 ( .A(G164), .B(G2078), .ZN(n948) );
  NAND2_X1 U1041 ( .A1(n949), .A2(n948), .ZN(n950) );
  XOR2_X1 U1042 ( .A(KEYINPUT50), .B(n950), .Z(n951) );
  XNOR2_X1 U1043 ( .A(KEYINPUT115), .B(n951), .ZN(n952) );
  NOR2_X1 U1044 ( .A1(n953), .A2(n952), .ZN(n960) );
  XOR2_X1 U1045 ( .A(G2090), .B(G162), .Z(n954) );
  NOR2_X1 U1046 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1047 ( .A(n956), .B(KEYINPUT51), .ZN(n957) );
  NOR2_X1 U1048 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1049 ( .A1(n960), .A2(n959), .ZN(n961) );
  NOR2_X1 U1050 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1051 ( .A(n964), .B(n963), .ZN(n965) );
  NAND2_X1 U1052 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1053 ( .A1(n967), .A2(G29), .ZN(n1023) );
  XNOR2_X1 U1054 ( .A(G2084), .B(G34), .ZN(n968) );
  XNOR2_X1 U1055 ( .A(n968), .B(KEYINPUT54), .ZN(n986) );
  XOR2_X1 U1056 ( .A(G2090), .B(G35), .Z(n969) );
  XNOR2_X1 U1057 ( .A(KEYINPUT117), .B(n969), .ZN(n983) );
  XNOR2_X1 U1058 ( .A(G2067), .B(G26), .ZN(n971) );
  XNOR2_X1 U1059 ( .A(G1996), .B(G32), .ZN(n970) );
  NOR2_X1 U1060 ( .A1(n971), .A2(n970), .ZN(n976) );
  XNOR2_X1 U1061 ( .A(n972), .B(G27), .ZN(n974) );
  XNOR2_X1 U1062 ( .A(G2072), .B(G33), .ZN(n973) );
  NOR2_X1 U1063 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1064 ( .A1(n976), .A2(n975), .ZN(n980) );
  XOR2_X1 U1065 ( .A(G1991), .B(G25), .Z(n977) );
  NAND2_X1 U1066 ( .A1(n977), .A2(G28), .ZN(n978) );
  XNOR2_X1 U1067 ( .A(KEYINPUT118), .B(n978), .ZN(n979) );
  NOR2_X1 U1068 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1069 ( .A(n981), .B(KEYINPUT53), .ZN(n982) );
  NOR2_X1 U1070 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1071 ( .A(n984), .B(KEYINPUT119), .ZN(n985) );
  NOR2_X1 U1072 ( .A1(n986), .A2(n985), .ZN(n1015) );
  NAND2_X1 U1073 ( .A1(KEYINPUT55), .A2(n1015), .ZN(n987) );
  NAND2_X1 U1074 ( .A1(G11), .A2(n987), .ZN(n1021) );
  XNOR2_X1 U1075 ( .A(G20), .B(n988), .ZN(n992) );
  XNOR2_X1 U1076 ( .A(G1341), .B(G19), .ZN(n990) );
  XNOR2_X1 U1077 ( .A(G1981), .B(G6), .ZN(n989) );
  NOR2_X1 U1078 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1079 ( .A1(n992), .A2(n991), .ZN(n995) );
  XOR2_X1 U1080 ( .A(KEYINPUT59), .B(G1348), .Z(n993) );
  XNOR2_X1 U1081 ( .A(G4), .B(n993), .ZN(n994) );
  NOR2_X1 U1082 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1083 ( .A(KEYINPUT60), .B(n996), .Z(n998) );
  XNOR2_X1 U1084 ( .A(G1966), .B(G21), .ZN(n997) );
  NOR2_X1 U1085 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1086 ( .A(KEYINPUT124), .B(n999), .Z(n1001) );
  XNOR2_X1 U1087 ( .A(G1961), .B(G5), .ZN(n1000) );
  NOR2_X1 U1088 ( .A1(n1001), .A2(n1000), .ZN(n1010) );
  XOR2_X1 U1089 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n1008) );
  XNOR2_X1 U1090 ( .A(G1971), .B(G22), .ZN(n1003) );
  XNOR2_X1 U1091 ( .A(G23), .B(G1976), .ZN(n1002) );
  NOR2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1006) );
  XNOR2_X1 U1093 ( .A(G1986), .B(KEYINPUT125), .ZN(n1004) );
  XNOR2_X1 U1094 ( .A(n1004), .B(G24), .ZN(n1005) );
  NAND2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1096 ( .A(n1008), .B(n1007), .ZN(n1009) );
  NAND2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1098 ( .A(n1011), .B(KEYINPUT127), .ZN(n1012) );
  XNOR2_X1 U1099 ( .A(KEYINPUT61), .B(n1012), .ZN(n1014) );
  INV_X1 U1100 ( .A(G16), .ZN(n1013) );
  NAND2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1019) );
  NOR2_X1 U1102 ( .A1(KEYINPUT55), .A2(G29), .ZN(n1017) );
  INV_X1 U1103 ( .A(n1015), .ZN(n1016) );
  NAND2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NOR2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1107 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1108 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1109 ( .A(n1026), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

