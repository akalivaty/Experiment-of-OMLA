//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 1 1 0 0 0 0 1 1 0 1 0 1 0 0 0 1 0 1 1 0 0 1 0 0 1 0 0 0 1 0 0 0 1 0 0 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n781, new_n782, new_n783, new_n784, new_n786,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n873, new_n874, new_n875, new_n876, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT27), .B(G183gat), .ZN(new_n203));
  INV_X1    g002(.A(G190gat), .ZN(new_n204));
  AND3_X1   g003(.A1(new_n203), .A2(KEYINPUT28), .A3(new_n204), .ZN(new_n205));
  AOI21_X1  g004(.A(KEYINPUT28), .B1(new_n203), .B2(new_n204), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208));
  OAI211_X1 g007(.A(KEYINPUT67), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n209), .B(new_n210), .C1(new_n212), .C2(KEYINPUT26), .ZN(new_n213));
  AOI21_X1  g012(.A(KEYINPUT67), .B1(new_n212), .B2(KEYINPUT26), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n208), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  OR2_X1    g014(.A1(new_n207), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT65), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n211), .B1(KEYINPUT23), .B2(new_n210), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT23), .ZN(new_n219));
  NOR3_X1   g018(.A1(new_n219), .A2(G169gat), .A3(G176gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n217), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  NOR2_X1   g020(.A1(G183gat), .A2(G190gat), .ZN(new_n222));
  AND2_X1   g021(.A1(G183gat), .A2(G190gat), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n222), .B1(new_n223), .B2(KEYINPUT24), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT24), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT64), .ZN(new_n227));
  AOI21_X1  g026(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT64), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n224), .A2(new_n227), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n211), .A2(KEYINPUT23), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n219), .B1(G169gat), .B2(G176gat), .ZN(new_n233));
  OAI211_X1 g032(.A(KEYINPUT65), .B(new_n232), .C1(new_n233), .C2(new_n211), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n221), .A2(new_n231), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT25), .ZN(new_n236));
  AND2_X1   g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n238));
  OAI211_X1 g037(.A(KEYINPUT25), .B(new_n232), .C1(new_n233), .C2(new_n211), .ZN(new_n239));
  NAND3_X1  g038(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  NOR3_X1   g040(.A1(new_n241), .A2(new_n228), .A3(new_n222), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n238), .B1(new_n239), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n210), .A2(KEYINPUT23), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n220), .B1(new_n212), .B2(new_n244), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n226), .B(new_n240), .C1(G183gat), .C2(G190gat), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n245), .A2(KEYINPUT66), .A3(KEYINPUT25), .A4(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n216), .B1(new_n237), .B2(new_n248), .ZN(new_n249));
  XOR2_X1   g048(.A(G113gat), .B(G120gat), .Z(new_n250));
  XNOR2_X1  g049(.A(G127gat), .B(G134gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(KEYINPUT69), .B(KEYINPUT1), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n250), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G113gat), .B(G120gat), .ZN(new_n254));
  OAI22_X1  g053(.A1(new_n254), .A2(KEYINPUT1), .B1(G127gat), .B2(G134gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(KEYINPUT68), .B(G127gat), .ZN(new_n256));
  INV_X1    g055(.A(G134gat), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n253), .B1(new_n255), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT70), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT70), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n253), .B(new_n261), .C1(new_n255), .C2(new_n258), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n249), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n207), .A2(new_n215), .ZN(new_n266));
  AND2_X1   g065(.A1(new_n243), .A2(new_n247), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n235), .A2(new_n236), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(new_n263), .ZN(new_n270));
  NAND2_X1  g069(.A1(G227gat), .A2(G233gat), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n265), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT32), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT33), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  XOR2_X1   g075(.A(G15gat), .B(G43gat), .Z(new_n277));
  XNOR2_X1  g076(.A(G71gat), .B(G99gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n274), .A2(new_n276), .A3(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n279), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n273), .B(KEYINPUT32), .C1(new_n275), .C2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT74), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n268), .A2(new_n243), .A3(new_n247), .ZN(new_n285));
  AND3_X1   g084(.A1(new_n285), .A2(new_n263), .A3(new_n216), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n263), .B1(new_n285), .B2(new_n216), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n288));
  NOR3_X1   g087(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT71), .B1(new_n265), .B2(new_n270), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n271), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n291), .A2(KEYINPUT72), .A3(KEYINPUT34), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n288), .B1(new_n286), .B2(new_n287), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n265), .A2(new_n270), .A3(KEYINPUT71), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n272), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT34), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n293), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n265), .A2(new_n270), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n299), .A2(new_n297), .A3(new_n271), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT73), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT73), .ZN(new_n302));
  NAND4_X1  g101(.A1(new_n299), .A2(new_n302), .A3(new_n297), .A4(new_n271), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n284), .A2(new_n292), .A3(new_n298), .A4(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n298), .A2(new_n292), .A3(new_n304), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT74), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n307), .B1(new_n280), .B2(new_n282), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n202), .B1(new_n305), .B2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n283), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n283), .A2(new_n298), .A3(new_n292), .A4(new_n304), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT36), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT78), .ZN(new_n316));
  XNOR2_X1  g115(.A(G197gat), .B(G204gat), .ZN(new_n317));
  INV_X1    g116(.A(G211gat), .ZN(new_n318));
  OR2_X1    g117(.A1(KEYINPUT75), .A2(G218gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(KEYINPUT75), .A2(G218gat), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n317), .B1(new_n321), .B2(KEYINPUT22), .ZN(new_n322));
  XOR2_X1   g121(.A(G211gat), .B(G218gat), .Z(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n323), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n325), .B(new_n317), .C1(KEYINPUT22), .C2(new_n321), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(G226gat), .ZN(new_n328));
  INV_X1    g127(.A(G233gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NOR3_X1   g130(.A1(new_n269), .A2(KEYINPUT77), .A3(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT29), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n249), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(KEYINPUT77), .B1(new_n335), .B2(new_n331), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n269), .A2(new_n331), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n327), .B(new_n333), .C1(new_n336), .C2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G8gat), .B(G36gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(G64gat), .B(G92gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n339), .B(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT76), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n331), .B1(new_n269), .B2(KEYINPUT29), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n249), .A2(new_n330), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n327), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n343), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  AOI211_X1 g147(.A(KEYINPUT76), .B(new_n327), .C1(new_n344), .C2(new_n345), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n338), .B(new_n342), .C1(new_n348), .C2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT30), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n316), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n330), .B1(new_n249), .B2(new_n334), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n347), .B1(new_n353), .B2(new_n337), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT76), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n346), .A2(new_n343), .A3(new_n347), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT77), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n344), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n332), .B1(new_n358), .B2(new_n345), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n355), .A2(new_n356), .B1(new_n359), .B2(new_n327), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n360), .A2(KEYINPUT78), .A3(KEYINPUT30), .A4(new_n342), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n352), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT5), .ZN(new_n363));
  XNOR2_X1  g162(.A(G155gat), .B(G162gat), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT80), .ZN(new_n366));
  XNOR2_X1  g165(.A(KEYINPUT81), .B(G155gat), .ZN(new_n367));
  INV_X1    g166(.A(G162gat), .ZN(new_n368));
  OAI21_X1  g167(.A(KEYINPUT2), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(G141gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT79), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT79), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(G141gat), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n371), .A2(new_n373), .A3(G148gat), .ZN(new_n374));
  INV_X1    g173(.A(G148gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(G141gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT80), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n364), .A2(new_n378), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n366), .A2(new_n369), .A3(new_n377), .A4(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(G141gat), .B(G148gat), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n365), .B1(KEYINPUT2), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n383), .B(new_n259), .ZN(new_n384));
  NAND2_X1  g183(.A1(G225gat), .A2(G233gat), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n363), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT3), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n388), .B1(new_n380), .B2(new_n382), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT82), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(KEYINPUT83), .B(KEYINPUT3), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n380), .A2(new_n382), .A3(new_n392), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n259), .B(new_n393), .C1(new_n389), .C2(KEYINPUT82), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n385), .B1(new_n391), .B2(new_n394), .ZN(new_n395));
  NOR3_X1   g194(.A1(new_n383), .A2(KEYINPUT4), .A3(new_n259), .ZN(new_n396));
  INV_X1    g195(.A(new_n383), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n397), .A2(new_n260), .A3(new_n262), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n396), .B1(new_n398), .B2(KEYINPUT4), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n387), .B1(new_n395), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(KEYINPUT4), .B1(new_n383), .B2(new_n259), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT85), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI211_X1 g202(.A(KEYINPUT85), .B(KEYINPUT4), .C1(new_n383), .C2(new_n259), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT4), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n397), .A2(new_n405), .A3(new_n260), .A4(new_n262), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n403), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  OR2_X1    g206(.A1(new_n389), .A2(KEYINPUT82), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n408), .A2(new_n259), .A3(new_n390), .A4(new_n393), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n386), .A2(KEYINPUT5), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n407), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n400), .A2(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(G1gat), .B(G29gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n413), .B(KEYINPUT0), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n414), .B(KEYINPUT84), .ZN(new_n415));
  XNOR2_X1  g214(.A(G57gat), .B(G85gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n415), .B(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n412), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT6), .ZN(new_n419));
  INV_X1    g218(.A(new_n417), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n400), .A2(new_n420), .A3(new_n411), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n418), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n412), .A2(KEYINPUT6), .A3(new_n417), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n355), .A2(new_n356), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n342), .B1(new_n425), .B2(new_n338), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n350), .B1(new_n426), .B2(new_n351), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n362), .A2(new_n424), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(KEYINPUT29), .B1(new_n324), .B2(new_n326), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n383), .B1(new_n429), .B2(KEYINPUT3), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT86), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT86), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n432), .B(new_n383), .C1(new_n429), .C2(KEYINPUT3), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(G228gat), .A2(G233gat), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n393), .A2(new_n334), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n435), .B1(new_n436), .B2(new_n347), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n436), .A2(new_n347), .ZN(new_n439));
  INV_X1    g238(.A(new_n392), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n383), .B1(new_n429), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(new_n435), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n438), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT87), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n444), .A2(new_n445), .A3(G22gat), .ZN(new_n446));
  AOI22_X1  g245(.A1(new_n434), .A2(new_n437), .B1(new_n435), .B2(new_n442), .ZN(new_n447));
  INV_X1    g246(.A(G22gat), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT87), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  XNOR2_X1  g248(.A(G78gat), .B(G106gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(KEYINPUT31), .B(G50gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n450), .B(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n452), .B1(new_n447), .B2(new_n448), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n446), .A2(new_n449), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT88), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n455), .B1(new_n447), .B2(new_n448), .ZN(new_n456));
  AND3_X1   g255(.A1(new_n438), .A2(new_n448), .A3(new_n443), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n452), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NOR3_X1   g257(.A1(new_n444), .A2(new_n455), .A3(G22gat), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n454), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n428), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n315), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT89), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n315), .A2(new_n461), .A3(KEYINPUT89), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT37), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n342), .B1(new_n360), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT38), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n338), .B1(new_n348), .B2(new_n349), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n468), .B1(new_n469), .B2(KEYINPUT37), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n338), .B(new_n466), .C1(new_n348), .C2(new_n349), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n466), .B1(new_n346), .B2(new_n327), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n333), .B1(new_n336), .B2(new_n337), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n473), .B1(new_n474), .B2(new_n327), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n472), .A2(new_n341), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(new_n468), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n471), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n423), .A2(KEYINPUT90), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT90), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n412), .A2(new_n480), .A3(KEYINPUT6), .A4(new_n417), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n422), .A2(new_n479), .A3(new_n350), .A4(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n460), .B1(new_n478), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n362), .A2(new_n427), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT40), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n385), .B1(new_n407), .B2(new_n409), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT39), .B1(new_n384), .B2(new_n386), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n420), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AOI211_X1 g288(.A(KEYINPUT39), .B(new_n385), .C1(new_n407), .C2(new_n409), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n486), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OR3_X1    g290(.A1(new_n489), .A2(new_n486), .A3(new_n490), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n492), .A2(new_n418), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n485), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n484), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n464), .A2(new_n465), .A3(new_n495), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n422), .A2(new_n479), .A3(new_n481), .ZN(new_n497));
  XOR2_X1   g296(.A(KEYINPUT92), .B(KEYINPUT35), .Z(new_n498));
  OAI211_X1 g297(.A(new_n454), .B(new_n498), .C1(new_n458), .C2(new_n459), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n312), .A2(new_n313), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT91), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT30), .B1(new_n360), .B2(new_n342), .ZN(new_n504));
  AOI22_X1  g303(.A1(new_n352), .A2(new_n361), .B1(new_n504), .B2(new_n350), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n312), .A2(KEYINPUT91), .A3(new_n313), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n500), .A2(new_n503), .A3(new_n505), .A4(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n452), .ZN(new_n508));
  AOI21_X1  g307(.A(KEYINPUT88), .B1(new_n444), .B2(G22gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n447), .A2(new_n448), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n459), .ZN(new_n512));
  AND2_X1   g311(.A1(new_n449), .A2(new_n453), .ZN(new_n513));
  AOI22_X1  g312(.A1(new_n511), .A2(new_n512), .B1(new_n513), .B2(new_n446), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n514), .A2(new_n305), .A3(new_n309), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT35), .B1(new_n515), .B2(new_n428), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n507), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n496), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(G15gat), .B(G22gat), .ZN(new_n519));
  OR2_X1    g318(.A1(new_n519), .A2(KEYINPUT96), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(KEYINPUT96), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT16), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n522), .B1(new_n523), .B2(G1gat), .ZN(new_n524));
  INV_X1    g323(.A(G1gat), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n520), .A2(new_n525), .A3(new_n521), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(G8gat), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n528), .B1(new_n526), .B2(KEYINPUT97), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n524), .B(new_n526), .C1(KEYINPUT97), .C2(new_n528), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(G43gat), .B(G50gat), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n533), .A2(KEYINPUT15), .ZN(new_n534));
  NOR2_X1   g333(.A1(G29gat), .A2(G36gat), .ZN(new_n535));
  AND2_X1   g334(.A1(new_n535), .A2(KEYINPUT14), .ZN(new_n536));
  NAND2_X1  g335(.A1(G29gat), .A2(G36gat), .ZN(new_n537));
  OAI211_X1 g336(.A(KEYINPUT94), .B(new_n537), .C1(new_n535), .C2(KEYINPUT14), .ZN(new_n538));
  NOR3_X1   g337(.A1(new_n534), .A2(new_n536), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n533), .A2(KEYINPUT15), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g340(.A(KEYINPUT15), .B(new_n533), .C1(new_n538), .C2(new_n536), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT95), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT95), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n541), .A2(new_n545), .A3(new_n542), .ZN(new_n546));
  AND3_X1   g345(.A1(new_n532), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n543), .A2(KEYINPUT17), .ZN(new_n548));
  AND2_X1   g347(.A1(new_n544), .A2(new_n546), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n548), .B1(new_n549), .B2(KEYINPUT17), .ZN(new_n550));
  AND2_X1   g349(.A1(new_n530), .A2(new_n531), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n547), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(G229gat), .A2(G233gat), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n552), .A2(KEYINPUT18), .A3(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n549), .B(new_n532), .ZN(new_n555));
  XOR2_X1   g354(.A(new_n553), .B(KEYINPUT13), .Z(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n549), .A2(new_n532), .ZN(new_n558));
  AOI21_X1  g357(.A(KEYINPUT17), .B1(new_n544), .B2(new_n546), .ZN(new_n559));
  INV_X1    g358(.A(new_n548), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  OAI211_X1 g360(.A(new_n553), .B(new_n558), .C1(new_n561), .C2(new_n532), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT18), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n554), .A2(new_n557), .A3(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G113gat), .B(G141gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(KEYINPUT11), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(G169gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(KEYINPUT93), .B(G197gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT12), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n565), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n554), .A2(new_n557), .A3(new_n564), .A4(new_n571), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n518), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT102), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT101), .ZN(new_n578));
  NAND2_X1  g377(.A1(G99gat), .A2(G106gat), .ZN(new_n579));
  INV_X1    g378(.A(G85gat), .ZN(new_n580));
  INV_X1    g379(.A(G92gat), .ZN(new_n581));
  AOI22_X1  g380(.A1(KEYINPUT8), .A2(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT7), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n583), .B1(new_n580), .B2(new_n581), .ZN(new_n584));
  NAND3_X1  g383(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n582), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  XOR2_X1   g385(.A(G99gat), .B(G106gat), .Z(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n586), .B(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(G232gat), .A2(G233gat), .ZN(new_n590));
  AOI22_X1  g389(.A1(new_n549), .A2(new_n589), .B1(KEYINPUT41), .B2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n586), .B(new_n587), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n592), .B1(new_n559), .B2(new_n560), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G190gat), .B(G218gat), .ZN(new_n595));
  XOR2_X1   g394(.A(new_n595), .B(KEYINPUT100), .Z(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n578), .B1(new_n594), .B2(new_n597), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n591), .A2(new_n593), .A3(KEYINPUT101), .A4(new_n596), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n590), .A2(KEYINPUT41), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n594), .A2(new_n597), .ZN(new_n603));
  AND3_X1   g402(.A1(new_n600), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n602), .B1(new_n600), .B2(new_n603), .ZN(new_n605));
  XOR2_X1   g404(.A(G134gat), .B(G162gat), .Z(new_n606));
  NOR3_X1   g405(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n606), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n600), .A2(new_n603), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(new_n601), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n600), .A2(new_n602), .A3(new_n603), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n608), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n607), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G127gat), .B(G155gat), .ZN(new_n614));
  XOR2_X1   g413(.A(new_n614), .B(KEYINPUT99), .Z(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT98), .ZN(new_n617));
  OR2_X1    g416(.A1(G57gat), .A2(G64gat), .ZN(new_n618));
  NAND2_X1  g417(.A1(G57gat), .A2(G64gat), .ZN(new_n619));
  INV_X1    g418(.A(G71gat), .ZN(new_n620));
  INV_X1    g419(.A(G78gat), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n618), .B(new_n619), .C1(new_n622), .C2(KEYINPUT9), .ZN(new_n623));
  XOR2_X1   g422(.A(G71gat), .B(G78gat), .Z(new_n624));
  OR2_X1    g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT21), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n617), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n627), .A2(new_n617), .A3(new_n628), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n630), .A2(G231gat), .A3(G233gat), .A4(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(G231gat), .A2(G233gat), .ZN(new_n633));
  INV_X1    g432(.A(new_n631), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n633), .B1(new_n634), .B2(new_n629), .ZN(new_n635));
  XOR2_X1   g434(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n636));
  NAND3_X1  g435(.A1(new_n632), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n636), .B1(new_n632), .B2(new_n635), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n616), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n639), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n641), .A2(new_n615), .A3(new_n637), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n551), .B1(new_n628), .B2(new_n627), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n640), .A2(new_n642), .A3(new_n644), .ZN(new_n647));
  XOR2_X1   g446(.A(G183gat), .B(G211gat), .Z(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  AND3_X1   g448(.A1(new_n646), .A2(new_n647), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n649), .B1(new_n646), .B2(new_n647), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n625), .A2(new_n626), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(new_n589), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT10), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n592), .A2(new_n627), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n653), .A2(new_n589), .A3(KEYINPUT10), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(G230gat), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n660), .A2(new_n329), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n654), .A2(new_n656), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(new_n661), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(G120gat), .B(G148gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(G176gat), .B(G204gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n669), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n663), .A2(new_n665), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n613), .A2(new_n652), .A3(new_n674), .ZN(new_n675));
  NOR3_X1   g474(.A1(new_n576), .A2(new_n577), .A3(new_n675), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n507), .A2(new_n516), .ZN(new_n677));
  AOI22_X1  g476(.A1(new_n462), .A2(new_n463), .B1(new_n494), .B2(new_n484), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n677), .B1(new_n678), .B2(new_n465), .ZN(new_n679));
  INV_X1    g478(.A(new_n575), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n675), .ZN(new_n682));
  AOI21_X1  g481(.A(KEYINPUT102), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  OR2_X1    g482(.A1(new_n676), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n424), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g486(.A(KEYINPUT16), .B(G8gat), .Z(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT103), .ZN(new_n689));
  OAI211_X1 g488(.A(new_n485), .B(new_n689), .C1(new_n676), .C2(new_n683), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n690), .A2(KEYINPUT42), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT42), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n485), .B1(new_n676), .B2(new_n683), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n692), .B1(new_n693), .B2(G8gat), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n691), .B1(new_n690), .B2(new_n694), .ZN(G1325gat));
  NAND2_X1  g494(.A1(new_n503), .A2(new_n506), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  AOI21_X1  g496(.A(G15gat), .B1(new_n684), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n305), .A2(new_n309), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(KEYINPUT36), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n501), .A2(new_n202), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n700), .A2(new_n701), .A3(KEYINPUT104), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT104), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n703), .B1(new_n310), .B2(new_n314), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(G15gat), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT105), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n698), .B1(new_n684), .B2(new_n707), .ZN(G1326gat));
  OAI21_X1  g507(.A(new_n460), .B1(new_n676), .B2(new_n683), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(KEYINPUT106), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT106), .ZN(new_n711));
  OAI211_X1 g510(.A(new_n711), .B(new_n460), .C1(new_n676), .C2(new_n683), .ZN(new_n712));
  XNOR2_X1  g511(.A(KEYINPUT43), .B(G22gat), .ZN(new_n713));
  AND3_X1   g512(.A1(new_n710), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n713), .B1(new_n710), .B2(new_n712), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n714), .A2(new_n715), .ZN(G1327gat));
  INV_X1    g515(.A(new_n613), .ZN(new_n717));
  INV_X1    g516(.A(new_n652), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n717), .A2(new_n718), .A3(new_n674), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n576), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n721), .A2(G29gat), .A3(new_n424), .ZN(new_n722));
  XNOR2_X1  g521(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(new_n724));
  XOR2_X1   g523(.A(new_n673), .B(KEYINPUT108), .Z(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n718), .A2(new_n575), .A3(new_n726), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT109), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  AOI22_X1  g528(.A1(new_n467), .A2(new_n470), .B1(new_n476), .B2(new_n468), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n514), .B1(new_n730), .B2(new_n482), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n492), .A2(new_n418), .A3(new_n491), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n732), .B1(new_n362), .B2(new_n427), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n461), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n517), .B1(new_n705), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(KEYINPUT110), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT110), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n517), .B(new_n737), .C1(new_n705), .C2(new_n734), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n613), .A2(KEYINPUT44), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n736), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  AND2_X1   g539(.A1(new_n740), .A2(KEYINPUT111), .ZN(new_n741));
  OAI21_X1  g540(.A(KEYINPUT44), .B1(new_n679), .B2(new_n613), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT111), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n736), .A2(new_n743), .A3(new_n738), .A4(new_n739), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n685), .B(new_n729), .C1(new_n741), .C2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(G29gat), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n724), .A2(new_n747), .ZN(G1328gat));
  INV_X1    g547(.A(G36gat), .ZN(new_n749));
  OAI211_X1 g548(.A(new_n485), .B(new_n729), .C1(new_n741), .C2(new_n745), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n749), .B1(new_n750), .B2(KEYINPUT112), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n751), .B1(KEYINPUT112), .B2(new_n750), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n720), .A2(new_n749), .A3(new_n485), .ZN(new_n753));
  XOR2_X1   g552(.A(new_n753), .B(KEYINPUT46), .Z(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(G1329gat));
  INV_X1    g554(.A(G43gat), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n756), .B1(new_n721), .B2(new_n696), .ZN(new_n757));
  INV_X1    g556(.A(new_n705), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n758), .A2(new_n756), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n729), .B(new_n759), .C1(new_n741), .C2(new_n745), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g561(.A(G50gat), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n763), .B1(new_n721), .B2(new_n514), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n514), .A2(new_n763), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n729), .B(new_n765), .C1(new_n741), .C2(new_n745), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(KEYINPUT48), .ZN(G1331gat));
  AND2_X1   g567(.A1(new_n736), .A2(new_n738), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n606), .B1(new_n604), .B2(new_n605), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n610), .A2(new_n611), .A3(new_n608), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n652), .A2(new_n770), .A3(new_n771), .A4(new_n680), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n772), .A2(new_n726), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n769), .A2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n685), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(G57gat), .ZN(G1332gat));
  AOI211_X1 g576(.A(new_n505), .B(new_n774), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n778));
  NOR2_X1   g577(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n778), .B(new_n779), .ZN(G1333gat));
  OAI21_X1  g579(.A(G71gat), .B1(new_n774), .B2(new_n758), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n697), .A2(new_n620), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n781), .B1(new_n774), .B2(new_n782), .ZN(new_n783));
  XOR2_X1   g582(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n784));
  XNOR2_X1  g583(.A(new_n783), .B(new_n784), .ZN(G1334gat));
  NOR2_X1   g584(.A1(new_n774), .A2(new_n514), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(new_n621), .ZN(G1335gat));
  NAND2_X1  g586(.A1(new_n718), .A2(new_n680), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n788), .A2(new_n613), .ZN(new_n789));
  AND3_X1   g588(.A1(new_n735), .A2(KEYINPUT51), .A3(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(KEYINPUT51), .B1(new_n735), .B2(new_n789), .ZN(new_n791));
  OR2_X1    g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n792), .A2(new_n580), .A3(new_n685), .A4(new_n673), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n788), .A2(new_n674), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n742), .A2(new_n744), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n740), .A2(KEYINPUT111), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n795), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n798), .A2(new_n685), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n793), .B1(new_n799), .B2(new_n580), .ZN(G1336gat));
  NAND3_X1  g599(.A1(new_n485), .A2(new_n581), .A3(new_n725), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(KEYINPUT114), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n802), .B1(new_n790), .B2(new_n791), .ZN(new_n803));
  NAND2_X1  g602(.A1(KEYINPUT115), .A2(KEYINPUT52), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n485), .B(new_n794), .C1(new_n741), .C2(new_n745), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n805), .B1(new_n806), .B2(G92gat), .ZN(new_n807));
  NOR2_X1   g606(.A1(KEYINPUT115), .A2(KEYINPUT52), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  AOI211_X1 g609(.A(new_n805), .B(new_n808), .C1(new_n806), .C2(G92gat), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n810), .A2(new_n811), .ZN(G1337gat));
  NAND2_X1  g611(.A1(new_n798), .A2(new_n705), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(G99gat), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n696), .A2(G99gat), .A3(new_n674), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n792), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n816), .ZN(G1338gat));
  INV_X1    g616(.A(G106gat), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n818), .B1(new_n798), .B2(new_n460), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n726), .A2(G106gat), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n792), .A2(new_n460), .A3(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(KEYINPUT53), .B1(new_n819), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n794), .B1(new_n741), .B2(new_n745), .ZN(new_n824));
  OAI21_X1  g623(.A(G106gat), .B1(new_n824), .B2(new_n514), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT53), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n825), .A2(new_n826), .A3(new_n821), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n823), .A2(new_n827), .ZN(G1339gat));
  NOR2_X1   g627(.A1(new_n552), .A2(new_n553), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n555), .A2(new_n556), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n570), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n574), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n657), .A2(new_n658), .A3(new_n661), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n663), .A2(KEYINPUT54), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n661), .B1(new_n657), .B2(new_n658), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n671), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n834), .A2(KEYINPUT55), .A3(new_n837), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n838), .A2(new_n672), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n834), .A2(new_n837), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT55), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n832), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n844), .B1(new_n607), .B2(new_n612), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n832), .A2(new_n674), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n843), .B1(new_n573), .B2(new_n574), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n770), .B(new_n771), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n652), .B1(new_n845), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n772), .A2(new_n673), .ZN(new_n850));
  OR2_X1    g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n485), .A2(new_n424), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n696), .A2(new_n460), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n855), .B(KEYINPUT116), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n856), .A2(G113gat), .A3(new_n575), .ZN(new_n857));
  INV_X1    g656(.A(G113gat), .ZN(new_n858));
  INV_X1    g657(.A(new_n515), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n853), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n858), .B1(new_n860), .B2(new_n680), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n857), .A2(new_n861), .ZN(G1340gat));
  NAND3_X1  g661(.A1(new_n856), .A2(G120gat), .A3(new_n725), .ZN(new_n863));
  INV_X1    g662(.A(G120gat), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n864), .B1(new_n860), .B2(new_n674), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n863), .A2(new_n865), .ZN(G1341gat));
  NOR2_X1   g665(.A1(new_n860), .A2(new_n718), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(KEYINPUT117), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n868), .A2(new_n256), .ZN(new_n869));
  OR2_X1    g668(.A1(new_n867), .A2(KEYINPUT117), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n718), .A2(new_n256), .ZN(new_n871));
  AOI22_X1  g670(.A1(new_n869), .A2(new_n870), .B1(new_n856), .B2(new_n871), .ZN(G1342gat));
  NAND2_X1  g671(.A1(new_n853), .A2(new_n717), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n873), .A2(G134gat), .A3(new_n515), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n874), .B(KEYINPUT56), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n856), .A2(new_n717), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n875), .B1(new_n876), .B2(new_n257), .ZN(G1343gat));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n514), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n840), .A2(KEYINPUT118), .ZN(new_n880));
  XNOR2_X1  g679(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n840), .A2(KEYINPUT118), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n839), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n884), .B1(new_n573), .B2(new_n574), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n771), .B(new_n770), .C1(new_n885), .C2(new_n846), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n652), .B1(new_n886), .B2(new_n845), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n879), .B1(new_n887), .B2(new_n850), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(KEYINPUT120), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n460), .B1(new_n849), .B2(new_n850), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n878), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT120), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n892), .B(new_n879), .C1(new_n887), .C2(new_n850), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n889), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n758), .A2(new_n852), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n894), .A2(new_n575), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n371), .A2(new_n373), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n705), .A2(new_n514), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n680), .A2(G141gat), .ZN(new_n901));
  AND4_X1   g700(.A1(new_n851), .A2(new_n852), .A3(new_n900), .A4(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n899), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(KEYINPUT58), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT58), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n899), .A2(new_n903), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n905), .A2(KEYINPUT121), .A3(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT121), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n906), .B1(new_n899), .B2(new_n903), .ZN(new_n910));
  AOI211_X1 g709(.A(KEYINPUT58), .B(new_n902), .C1(new_n897), .C2(new_n898), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n908), .A2(new_n912), .ZN(G1344gat));
  NAND2_X1  g712(.A1(new_n853), .A2(new_n900), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n915), .A2(new_n375), .A3(new_n673), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n375), .A2(KEYINPUT59), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n894), .A2(new_n896), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n917), .B1(new_n918), .B2(new_n674), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT122), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n890), .A2(KEYINPUT57), .ZN(new_n922));
  OAI211_X1 g721(.A(new_n878), .B(new_n460), .C1(new_n887), .C2(new_n850), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n896), .A2(new_n673), .ZN(new_n925));
  OAI21_X1  g724(.A(G148gat), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(KEYINPUT59), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n927), .B1(new_n919), .B2(new_n920), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n916), .B1(new_n921), .B2(new_n928), .ZN(G1345gat));
  NAND3_X1  g728(.A1(new_n915), .A2(new_n367), .A3(new_n652), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n918), .A2(new_n718), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n930), .B1(new_n931), .B2(new_n367), .ZN(G1346gat));
  INV_X1    g731(.A(new_n900), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n873), .A2(G162gat), .A3(new_n933), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT123), .ZN(new_n935));
  OAI21_X1  g734(.A(G162gat), .B1(new_n918), .B2(new_n613), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(G1347gat));
  NOR2_X1   g736(.A1(new_n505), .A2(new_n685), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n851), .A2(new_n859), .A3(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(G169gat), .B1(new_n940), .B2(new_n575), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n851), .A2(new_n938), .ZN(new_n942));
  INV_X1    g741(.A(new_n854), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n575), .A2(G169gat), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n941), .B1(new_n944), .B2(new_n945), .ZN(G1348gat));
  INV_X1    g745(.A(new_n944), .ZN(new_n947));
  OAI21_X1  g746(.A(G176gat), .B1(new_n947), .B2(new_n726), .ZN(new_n948));
  INV_X1    g747(.A(G176gat), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n940), .A2(new_n949), .A3(new_n673), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n948), .A2(new_n950), .ZN(G1349gat));
  NAND3_X1  g750(.A1(new_n940), .A2(new_n203), .A3(new_n652), .ZN(new_n952));
  OAI21_X1  g751(.A(G183gat), .B1(new_n947), .B2(new_n718), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n954), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g754(.A1(new_n940), .A2(new_n204), .A3(new_n717), .ZN(new_n956));
  OAI21_X1  g755(.A(G190gat), .B1(new_n947), .B2(new_n613), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n957), .A2(KEYINPUT61), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n957), .A2(KEYINPUT61), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(G1351gat));
  NOR2_X1   g759(.A1(new_n942), .A2(new_n933), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(KEYINPUT124), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT124), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n963), .B1(new_n942), .B2(new_n933), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  INV_X1    g764(.A(G197gat), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n965), .A2(new_n966), .A3(new_n575), .ZN(new_n967));
  INV_X1    g766(.A(new_n924), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n705), .A2(new_n685), .A3(new_n505), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g769(.A(G197gat), .B1(new_n970), .B2(new_n680), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n967), .A2(new_n971), .ZN(G1352gat));
  OAI21_X1  g771(.A(G204gat), .B1(new_n970), .B2(new_n726), .ZN(new_n973));
  INV_X1    g772(.A(G204gat), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n961), .A2(new_n974), .A3(new_n673), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(KEYINPUT125), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT125), .ZN(new_n977));
  NAND4_X1  g776(.A1(new_n961), .A2(new_n977), .A3(new_n974), .A4(new_n673), .ZN(new_n978));
  AND3_X1   g777(.A1(new_n976), .A2(KEYINPUT62), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g778(.A(KEYINPUT62), .B1(new_n976), .B2(new_n978), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n973), .B1(new_n979), .B2(new_n980), .ZN(G1353gat));
  NAND3_X1  g780(.A1(new_n965), .A2(new_n318), .A3(new_n652), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n968), .A2(new_n652), .A3(new_n969), .ZN(new_n983));
  AOI21_X1  g782(.A(KEYINPUT63), .B1(new_n983), .B2(G211gat), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT126), .ZN(new_n985));
  AND2_X1   g784(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n983), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n987), .B1(new_n984), .B2(new_n985), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n982), .B1(new_n986), .B2(new_n988), .ZN(G1354gat));
  AOI211_X1 g788(.A(new_n613), .B(new_n970), .C1(new_n319), .C2(new_n320), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n962), .A2(new_n717), .A3(new_n964), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT127), .ZN(new_n992));
  INV_X1    g791(.A(G218gat), .ZN(new_n993));
  AND3_X1   g792(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g793(.A(new_n992), .B1(new_n991), .B2(new_n993), .ZN(new_n995));
  NOR3_X1   g794(.A1(new_n990), .A2(new_n994), .A3(new_n995), .ZN(G1355gat));
endmodule


