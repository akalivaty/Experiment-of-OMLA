//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 0 0 0 1 1 1 1 1 1 0 0 1 1 0 0 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 1 1 0 1 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 0 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:50 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030;
  XNOR2_X1  g000(.A(KEYINPUT22), .B(G137), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  AND3_X1   g002(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n189));
  XOR2_X1   g003(.A(new_n187), .B(new_n189), .Z(new_n190));
  INV_X1    g004(.A(G140), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G125), .ZN(new_n192));
  INV_X1    g006(.A(G125), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G140), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT75), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT75), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n192), .A2(new_n194), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n196), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT76), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT76), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n196), .A2(new_n198), .A3(new_n202), .A4(new_n199), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n192), .A2(new_n194), .A3(KEYINPUT16), .ZN(new_n205));
  OR3_X1    g019(.A1(new_n193), .A2(KEYINPUT16), .A3(G140), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(G146), .ZN(new_n207));
  OR2_X1    g021(.A1(KEYINPUT67), .A2(G128), .ZN(new_n208));
  NAND2_X1  g022(.A1(KEYINPUT67), .A2(G128), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n208), .A2(KEYINPUT23), .A3(G119), .A4(new_n209), .ZN(new_n210));
  XOR2_X1   g024(.A(KEYINPUT74), .B(G110), .Z(new_n211));
  INV_X1    g025(.A(KEYINPUT23), .ZN(new_n212));
  INV_X1    g026(.A(G119), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n212), .B1(new_n213), .B2(G128), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT73), .ZN(new_n215));
  OAI22_X1  g029(.A1(new_n214), .A2(new_n215), .B1(new_n213), .B2(G128), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n213), .A2(G128), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n217), .A2(new_n215), .A3(KEYINPUT23), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n210), .B(new_n211), .C1(new_n216), .C2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n208), .A2(new_n209), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n217), .B1(new_n221), .B2(new_n213), .ZN(new_n222));
  XNOR2_X1  g036(.A(KEYINPUT24), .B(G110), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n220), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n204), .A2(new_n207), .A3(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n210), .B1(new_n216), .B2(new_n219), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G110), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n205), .A2(new_n206), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(new_n199), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(new_n207), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n228), .B(new_n231), .C1(new_n222), .C2(new_n223), .ZN(new_n232));
  AND3_X1   g046(.A1(new_n226), .A2(new_n232), .A3(KEYINPUT77), .ZN(new_n233));
  AOI21_X1  g047(.A(KEYINPUT77), .B1(new_n226), .B2(new_n232), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n190), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n190), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n226), .A2(new_n232), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT77), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  AND2_X1   g053(.A1(new_n235), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G217), .ZN(new_n241));
  INV_X1    g055(.A(G902), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n241), .B1(G234), .B2(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n243), .A2(G902), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n240), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT78), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n235), .A2(new_n242), .A3(new_n239), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT25), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT25), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n235), .A2(new_n250), .A3(new_n242), .A4(new_n239), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n249), .A2(new_n251), .A3(new_n243), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n240), .A2(KEYINPUT78), .A3(new_n244), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n247), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n199), .A2(G143), .ZN(new_n255));
  INV_X1    g069(.A(G143), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G146), .ZN(new_n257));
  AND2_X1   g071(.A1(KEYINPUT0), .A2(G128), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n255), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(G143), .B(G146), .ZN(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT0), .B(G128), .ZN(new_n261));
  OAI211_X1 g075(.A(new_n259), .B(KEYINPUT65), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n255), .A2(new_n257), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT65), .ZN(new_n264));
  INV_X1    g078(.A(new_n258), .ZN(new_n265));
  OR2_X1    g079(.A1(KEYINPUT0), .A2(G128), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n263), .A2(new_n264), .A3(new_n265), .A4(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n262), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT11), .ZN(new_n269));
  INV_X1    g083(.A(G134), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n269), .B1(new_n270), .B2(G137), .ZN(new_n271));
  INV_X1    g085(.A(G137), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n272), .A2(KEYINPUT11), .A3(G134), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n270), .A2(G137), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n271), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G131), .ZN(new_n276));
  INV_X1    g090(.A(G131), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n271), .A2(new_n273), .A3(new_n277), .A4(new_n274), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n268), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(KEYINPUT66), .B1(new_n270), .B2(G137), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT66), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n282), .A2(new_n272), .A3(G134), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n281), .A2(new_n283), .A3(new_n274), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(G131), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n255), .A2(KEYINPUT1), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n260), .B1(new_n221), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G128), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n288), .A2(KEYINPUT1), .ZN(new_n289));
  AND2_X1   g103(.A1(new_n260), .A2(new_n289), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n278), .B(new_n285), .C1(new_n287), .C2(new_n290), .ZN(new_n291));
  XOR2_X1   g105(.A(KEYINPUT2), .B(G113), .Z(new_n292));
  XNOR2_X1  g106(.A(G116), .B(G119), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n292), .A2(new_n293), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n280), .A2(new_n291), .A3(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(G237), .A2(G953), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G210), .ZN(new_n300));
  XNOR2_X1  g114(.A(new_n300), .B(KEYINPUT27), .ZN(new_n301));
  XNOR2_X1  g115(.A(KEYINPUT26), .B(G101), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n301), .B(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n298), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT68), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT68), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n298), .A2(new_n306), .A3(new_n303), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT30), .ZN(new_n309));
  AND2_X1   g123(.A1(new_n285), .A2(new_n278), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n260), .A2(new_n289), .ZN(new_n311));
  AND2_X1   g125(.A1(new_n221), .A2(new_n286), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n311), .B1(new_n312), .B2(new_n260), .ZN(new_n313));
  AOI22_X1  g127(.A1(new_n310), .A2(new_n313), .B1(new_n268), .B2(new_n279), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT64), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n309), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n280), .A2(new_n291), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n317), .A2(KEYINPUT64), .A3(KEYINPUT30), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n297), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(KEYINPUT31), .B1(new_n308), .B2(new_n319), .ZN(new_n320));
  AND3_X1   g134(.A1(new_n298), .A2(new_n306), .A3(new_n303), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n306), .B1(new_n298), .B2(new_n303), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OR2_X1    g137(.A1(new_n295), .A2(new_n296), .ZN(new_n324));
  AOI21_X1  g138(.A(KEYINPUT30), .B1(new_n317), .B2(KEYINPUT64), .ZN(new_n325));
  AOI211_X1 g139(.A(new_n315), .B(new_n309), .C1(new_n280), .C2(new_n291), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT31), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n323), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n303), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n324), .B1(new_n317), .B2(KEYINPUT69), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT69), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n314), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(KEYINPUT28), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT28), .ZN(new_n335));
  INV_X1    g149(.A(new_n291), .ZN(new_n336));
  AOI22_X1  g150(.A1(new_n262), .A2(new_n267), .B1(new_n276), .B2(new_n278), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n324), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n335), .B1(new_n338), .B2(new_n298), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n330), .B1(new_n334), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n320), .A2(new_n329), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G472), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n341), .A2(new_n342), .A3(new_n242), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(KEYINPUT70), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT32), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT70), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n341), .A2(new_n346), .A3(new_n342), .A4(new_n242), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n344), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n341), .A2(KEYINPUT32), .A3(new_n342), .A4(new_n242), .ZN(new_n349));
  AND2_X1   g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n298), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n319), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(KEYINPUT71), .B1(new_n352), .B2(new_n303), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n331), .A2(new_n333), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n339), .B1(new_n354), .B2(new_n335), .ZN(new_n355));
  AOI21_X1  g169(.A(KEYINPUT29), .B1(new_n355), .B2(new_n303), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT71), .ZN(new_n357));
  OAI211_X1 g171(.A(new_n357), .B(new_n330), .C1(new_n319), .C2(new_n351), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n353), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  NOR3_X1   g173(.A1(new_n334), .A2(new_n330), .A3(new_n339), .ZN(new_n360));
  AOI21_X1  g174(.A(G902), .B1(new_n360), .B2(KEYINPUT29), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(G472), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT72), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n362), .A2(KEYINPUT72), .A3(G472), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n254), .B1(new_n350), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g182(.A(G210), .B1(G237), .B2(G902), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n193), .B(new_n311), .C1(new_n312), .C2(new_n260), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n262), .A2(G125), .A3(new_n267), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G224), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n374), .A2(G953), .ZN(new_n375));
  XOR2_X1   g189(.A(new_n373), .B(new_n375), .Z(new_n376));
  INV_X1    g190(.A(G104), .ZN(new_n377));
  OAI21_X1  g191(.A(KEYINPUT3), .B1(new_n377), .B2(G107), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT3), .ZN(new_n379));
  INV_X1    g193(.A(G107), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(new_n380), .A3(G104), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n377), .A2(G107), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n378), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G101), .ZN(new_n384));
  INV_X1    g198(.A(G101), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n378), .A2(new_n381), .A3(new_n385), .A4(new_n382), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n384), .A2(KEYINPUT4), .A3(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT4), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n383), .A2(new_n388), .A3(G101), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n324), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n293), .A2(KEYINPUT5), .ZN(new_n391));
  INV_X1    g205(.A(G116), .ZN(new_n392));
  NOR3_X1   g206(.A1(new_n392), .A2(KEYINPUT5), .A3(G119), .ZN(new_n393));
  INV_X1    g207(.A(G113), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n396), .A2(new_n294), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT79), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n398), .B1(new_n377), .B2(G107), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n380), .A2(KEYINPUT79), .A3(G104), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n399), .A2(new_n382), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G101), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT80), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n403), .A3(new_n386), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n403), .B1(new_n402), .B2(new_n386), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n397), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  XNOR2_X1  g221(.A(G110), .B(G122), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n390), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT6), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n390), .A2(new_n407), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT82), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n408), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n410), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n411), .A2(KEYINPUT6), .A3(new_n413), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n376), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n402), .A2(new_n386), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n407), .B1(new_n418), .B2(new_n397), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n408), .B(KEYINPUT8), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT7), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n375), .A2(new_n423), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n371), .A2(new_n372), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n424), .B1(new_n371), .B2(new_n372), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n409), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n242), .B1(new_n422), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n370), .B1(new_n417), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n376), .ZN(new_n431));
  AOI22_X1  g245(.A1(new_n409), .A2(KEYINPUT6), .B1(new_n411), .B2(new_n413), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n411), .A2(KEYINPUT6), .A3(new_n413), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n431), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n428), .ZN(new_n435));
  AOI21_X1  g249(.A(G902), .B1(new_n435), .B2(new_n421), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n434), .A2(new_n436), .A3(new_n369), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n430), .A2(KEYINPUT83), .A3(new_n437), .ZN(new_n438));
  NOR3_X1   g252(.A1(new_n417), .A2(new_n429), .A3(new_n370), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT83), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(G214), .B1(G237), .B2(G902), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n438), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  OAI211_X1 g257(.A(KEYINPUT10), .B(new_n313), .C1(new_n405), .C2(new_n406), .ZN(new_n444));
  INV_X1    g258(.A(new_n279), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n288), .B1(new_n255), .B2(KEYINPUT1), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n311), .B1(new_n260), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n447), .A2(new_n386), .A3(new_n402), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT10), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n387), .A2(new_n268), .A3(new_n389), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n444), .A2(new_n445), .A3(new_n450), .A4(new_n451), .ZN(new_n452));
  XNOR2_X1  g266(.A(G110), .B(G140), .ZN(new_n453));
  AND2_X1   g267(.A1(new_n188), .A2(G227), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n453), .B(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n452), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT81), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n450), .A2(new_n451), .ZN(new_n460));
  OAI21_X1  g274(.A(KEYINPUT10), .B1(new_n287), .B2(new_n290), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n402), .A2(new_n386), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT80), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n461), .B1(new_n463), .B2(new_n404), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n279), .B1(new_n460), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n452), .A2(KEYINPUT81), .A3(new_n456), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n459), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n287), .A2(new_n290), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n463), .A2(new_n468), .A3(new_n404), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n448), .ZN(new_n470));
  AOI21_X1  g284(.A(KEYINPUT12), .B1(new_n470), .B2(new_n279), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT12), .ZN(new_n472));
  AOI211_X1 g286(.A(new_n472), .B(new_n445), .C1(new_n469), .C2(new_n448), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n452), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n455), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n467), .A2(new_n475), .A3(G469), .ZN(new_n476));
  INV_X1    g290(.A(G469), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n470), .A2(KEYINPUT12), .A3(new_n279), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n470), .A2(new_n279), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n472), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n457), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n456), .B1(new_n465), .B2(new_n452), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n477), .B(new_n242), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(G469), .A2(G902), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n476), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(KEYINPUT9), .B(G234), .ZN(new_n486));
  OAI21_X1  g300(.A(G221), .B1(new_n486), .B2(G902), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n443), .A2(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(G113), .B(G122), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n490), .B(new_n377), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT84), .ZN(new_n492));
  INV_X1    g306(.A(G214), .ZN(new_n493));
  NOR3_X1   g307(.A1(new_n493), .A2(G237), .A3(G953), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n492), .B1(new_n494), .B2(G143), .ZN(new_n495));
  INV_X1    g309(.A(G237), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n496), .A2(new_n188), .A3(G214), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n497), .A2(KEYINPUT84), .A3(new_n256), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n496), .A2(new_n188), .A3(G143), .A4(G214), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT85), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n299), .A2(KEYINPUT85), .A3(G143), .A4(G214), .ZN(new_n502));
  AOI22_X1  g316(.A1(new_n495), .A2(new_n498), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AND2_X1   g317(.A1(KEYINPUT18), .A2(G131), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n503), .B(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n195), .A2(G146), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n506), .B(KEYINPUT86), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n204), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  AOI211_X1 g323(.A(G143), .B(new_n492), .C1(new_n299), .C2(G214), .ZN(new_n510));
  AOI21_X1  g324(.A(KEYINPUT84), .B1(new_n497), .B2(new_n256), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AND2_X1   g326(.A1(new_n501), .A2(new_n502), .ZN(new_n513));
  OAI211_X1 g327(.A(KEYINPUT17), .B(G131), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  AND2_X1   g328(.A1(new_n230), .A2(new_n207), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n514), .A2(KEYINPUT87), .A3(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(G131), .B1(new_n512), .B2(new_n513), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n503), .A2(new_n277), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT17), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(KEYINPUT87), .B1(new_n514), .B2(new_n515), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n491), .B(new_n509), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(KEYINPUT88), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n514), .A2(new_n515), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT87), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n527), .A2(new_n520), .A3(new_n516), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT88), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n528), .A2(new_n529), .A3(new_n491), .A4(new_n509), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n524), .A2(new_n530), .ZN(new_n531));
  AND2_X1   g345(.A1(new_n528), .A2(new_n509), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n531), .B1(new_n491), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n242), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(G475), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n517), .A2(new_n518), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n195), .A2(KEYINPUT19), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n196), .A2(new_n198), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n538), .B1(new_n539), .B2(KEYINPUT19), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n537), .B(new_n207), .C1(G146), .C2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n491), .B1(new_n541), .B2(new_n509), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n531), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT89), .ZN(new_n545));
  NOR2_X1   g359(.A1(G475), .A2(G902), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT89), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n531), .A2(new_n547), .A3(new_n543), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n545), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT20), .ZN(new_n550));
  INV_X1    g364(.A(new_n546), .ZN(new_n551));
  AOI21_X1  g365(.A(KEYINPUT20), .B1(new_n551), .B2(KEYINPUT90), .ZN(new_n552));
  OR2_X1    g366(.A1(new_n551), .A2(KEYINPUT90), .ZN(new_n553));
  AND2_X1   g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n544), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n536), .B1(new_n550), .B2(new_n555), .ZN(new_n556));
  OR2_X1    g370(.A1(new_n392), .A2(G122), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n380), .B1(new_n557), .B2(KEYINPUT14), .ZN(new_n558));
  XOR2_X1   g372(.A(G116), .B(G122), .Z(new_n559));
  XOR2_X1   g373(.A(new_n558), .B(new_n559), .Z(new_n560));
  NAND3_X1  g374(.A1(new_n208), .A2(G143), .A3(new_n209), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT91), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n256), .A2(G128), .ZN(new_n563));
  AND3_X1   g377(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n562), .B1(new_n561), .B2(new_n563), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n270), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NOR3_X1   g381(.A1(new_n564), .A2(new_n565), .A3(new_n270), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n560), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  XOR2_X1   g383(.A(new_n563), .B(KEYINPUT13), .Z(new_n570));
  INV_X1    g384(.A(new_n561), .ZN(new_n571));
  OAI21_X1  g385(.A(G134), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n559), .B(G107), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n566), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n486), .A2(new_n241), .A3(G953), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n569), .A2(new_n574), .A3(new_n576), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n242), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT92), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(G478), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n584), .A2(KEYINPUT15), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n580), .A2(KEYINPUT92), .A3(new_n242), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n583), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  OR2_X1    g401(.A1(new_n581), .A2(new_n585), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n188), .A2(G952), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n590), .B1(G234), .B2(G237), .ZN(new_n591));
  AOI211_X1 g405(.A(new_n242), .B(new_n188), .C1(G234), .C2(G237), .ZN(new_n592));
  XNOR2_X1  g406(.A(KEYINPUT21), .B(G898), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n589), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(KEYINPUT93), .B1(new_n556), .B2(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n547), .B1(new_n531), .B2(new_n543), .ZN(new_n597));
  AOI211_X1 g411(.A(KEYINPUT89), .B(new_n542), .C1(new_n524), .C2(new_n530), .ZN(new_n598));
  NOR3_X1   g412(.A1(new_n597), .A2(new_n598), .A3(new_n551), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT20), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n555), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  AND4_X1   g415(.A1(KEYINPUT93), .A2(new_n601), .A3(new_n535), .A4(new_n595), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n368), .B(new_n489), .C1(new_n596), .C2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(G101), .ZN(G3));
  NAND2_X1  g418(.A1(new_n601), .A2(new_n535), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n583), .A2(new_n584), .A3(new_n586), .ZN(new_n606));
  OAI21_X1  g420(.A(KEYINPUT33), .B1(new_n576), .B2(KEYINPUT95), .ZN(new_n607));
  OR2_X1    g421(.A1(new_n580), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n580), .A2(new_n607), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n608), .A2(G478), .A3(new_n242), .A4(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n369), .B1(new_n434), .B2(new_n436), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n442), .B1(new_n439), .B2(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n613), .A2(new_n594), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n605), .A2(new_n611), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n341), .A2(new_n242), .ZN(new_n616));
  OAI21_X1  g430(.A(G472), .B1(new_n616), .B2(KEYINPUT94), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT94), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n618), .B1(new_n341), .B2(new_n242), .ZN(new_n619));
  OAI211_X1 g433(.A(new_n344), .B(new_n347), .C1(new_n617), .C2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n254), .ZN(new_n622));
  INV_X1    g436(.A(new_n488), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n615), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(KEYINPUT34), .B(G104), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G6));
  NOR2_X1   g441(.A1(new_n597), .A2(new_n598), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n600), .B1(new_n628), .B2(new_n546), .ZN(new_n629));
  NOR4_X1   g443(.A1(new_n597), .A2(new_n598), .A3(KEYINPUT20), .A4(new_n551), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n535), .B(new_n589), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n614), .ZN(new_n632));
  OR2_X1    g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n633), .A2(new_n624), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT35), .B(G107), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G9));
  NOR2_X1   g450(.A1(new_n236), .A2(KEYINPUT36), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n237), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n244), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n252), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(KEYINPUT96), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT96), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n252), .A2(new_n642), .A3(new_n639), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n644), .A2(new_n620), .ZN(new_n645));
  OAI211_X1 g459(.A(new_n489), .B(new_n645), .C1(new_n596), .C2(new_n602), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT37), .B(G110), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G12));
  NAND3_X1  g462(.A1(new_n623), .A2(new_n641), .A3(new_n643), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n649), .B1(new_n350), .B2(new_n367), .ZN(new_n650));
  INV_X1    g464(.A(G900), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n591), .B1(new_n592), .B2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n631), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n613), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n650), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G128), .ZN(G30));
  XOR2_X1   g470(.A(new_n652), .B(KEYINPUT39), .Z(new_n657));
  NAND3_X1  g471(.A1(new_n623), .A2(KEYINPUT98), .A3(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT98), .ZN(new_n659));
  INV_X1    g473(.A(new_n657), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n659), .B1(new_n488), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  OR2_X1    g476(.A1(new_n662), .A2(KEYINPUT40), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n323), .A2(new_n327), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n338), .A2(new_n298), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n342), .B1(new_n665), .B2(new_n330), .ZN(new_n666));
  AOI22_X1  g480(.A1(new_n664), .A2(new_n666), .B1(G472), .B2(G902), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT97), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n348), .A2(new_n349), .A3(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n640), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n671), .B1(KEYINPUT40), .B2(new_n662), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n589), .A2(new_n442), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n673), .B1(new_n601), .B2(new_n535), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n438), .A2(new_n441), .ZN(new_n675));
  XOR2_X1   g489(.A(new_n675), .B(KEYINPUT38), .Z(new_n676));
  NAND4_X1  g490(.A1(new_n663), .A2(new_n672), .A3(new_n674), .A4(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G143), .ZN(G45));
  INV_X1    g492(.A(new_n611), .ZN(new_n679));
  AOI211_X1 g493(.A(new_n652), .B(new_n679), .C1(new_n601), .C2(new_n535), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n650), .A2(new_n654), .A3(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT99), .B(G146), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G48));
  AOI21_X1  g497(.A(KEYINPUT72), .B1(new_n362), .B2(G472), .ZN(new_n684));
  AOI211_X1 g498(.A(new_n364), .B(new_n342), .C1(new_n359), .C2(new_n361), .ZN(new_n685));
  OAI211_X1 g499(.A(new_n348), .B(new_n349), .C1(new_n684), .C2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n480), .A2(new_n478), .ZN(new_n687));
  INV_X1    g501(.A(new_n457), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n482), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  OAI21_X1  g503(.A(G469), .B1(new_n689), .B2(G902), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n690), .A2(new_n487), .A3(new_n483), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(KEYINPUT100), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n686), .A2(new_n622), .A3(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n693), .A2(new_n615), .ZN(new_n694));
  XOR2_X1   g508(.A(KEYINPUT41), .B(G113), .Z(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G15));
  NOR2_X1   g510(.A1(new_n633), .A2(new_n693), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(new_n392), .ZN(G18));
  NOR2_X1   g512(.A1(new_n613), .A2(new_n691), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n699), .A2(new_n641), .A3(new_n643), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n700), .B1(new_n350), .B2(new_n367), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n701), .B1(new_n596), .B2(new_n602), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(KEYINPUT101), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT101), .ZN(new_n704));
  OAI211_X1 g518(.A(new_n701), .B(new_n704), .C1(new_n596), .C2(new_n602), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G119), .ZN(G21));
  XNOR2_X1  g521(.A(new_n616), .B(new_n342), .ZN(new_n708));
  AND2_X1   g522(.A1(new_n708), .A2(new_n622), .ZN(new_n709));
  INV_X1    g523(.A(new_n594), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n709), .A2(new_n710), .A3(new_n692), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n430), .A2(new_n437), .ZN(new_n712));
  AOI21_X1  g526(.A(KEYINPUT102), .B1(new_n674), .B2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(new_n673), .ZN(new_n714));
  INV_X1    g528(.A(new_n555), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n715), .B1(new_n549), .B2(KEYINPUT20), .ZN(new_n716));
  OAI211_X1 g530(.A(new_n712), .B(new_n714), .C1(new_n716), .C2(new_n536), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT102), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n711), .B1(new_n713), .B2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G122), .ZN(G24));
  AND2_X1   g535(.A1(new_n708), .A2(new_n640), .ZN(new_n722));
  AND2_X1   g536(.A1(new_n722), .A2(new_n699), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n680), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G125), .ZN(G27));
  INV_X1    g539(.A(KEYINPUT42), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n675), .A2(new_n442), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n727), .A2(new_n488), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n686), .A2(new_n728), .A3(new_n622), .ZN(new_n729));
  INV_X1    g543(.A(new_n652), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n605), .A2(new_n611), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n726), .B1(new_n729), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n343), .A2(new_n345), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n733), .A2(KEYINPUT103), .A3(new_n349), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n349), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT103), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n367), .A2(new_n734), .A3(new_n737), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n727), .A2(new_n726), .A3(new_n488), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n680), .A2(new_n738), .A3(new_n622), .A4(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n732), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G131), .ZN(G33));
  NAND3_X1  g556(.A1(new_n368), .A2(new_n653), .A3(new_n728), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G134), .ZN(G36));
  XNOR2_X1  g558(.A(new_n727), .B(KEYINPUT105), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n601), .A2(new_n535), .A3(new_n611), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT43), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n747), .B(new_n748), .C1(new_n605), .C2(KEYINPUT104), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT104), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n556), .B(new_n611), .C1(new_n750), .C2(KEYINPUT43), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n620), .A2(new_n640), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT44), .ZN(new_n756));
  OAI211_X1 g570(.A(KEYINPUT106), .B(new_n746), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n755), .A2(new_n756), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT106), .ZN(new_n760));
  AOI211_X1 g574(.A(new_n756), .B(new_n753), .C1(new_n749), .C2(new_n751), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n760), .B1(new_n761), .B2(new_n745), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g577(.A(KEYINPUT107), .B1(new_n759), .B2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n487), .ZN(new_n765));
  AOI21_X1  g579(.A(KEYINPUT45), .B1(new_n467), .B2(new_n475), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n477), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n467), .A2(new_n475), .A3(KEYINPUT45), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(KEYINPUT46), .B1(new_n769), .B2(new_n484), .ZN(new_n770));
  INV_X1    g584(.A(new_n483), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n769), .A2(KEYINPUT46), .A3(new_n484), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n765), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n657), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT107), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n762), .A2(new_n757), .A3(new_n777), .A4(new_n758), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n764), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(KEYINPUT108), .B(G137), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(KEYINPUT109), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n779), .B(new_n781), .ZN(G39));
  NOR2_X1   g596(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n774), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n784), .B1(new_n774), .B2(new_n785), .ZN(new_n786));
  NOR4_X1   g600(.A1(new_n731), .A2(new_n686), .A3(new_n622), .A4(new_n727), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G140), .ZN(G42));
  NAND3_X1  g603(.A1(new_n622), .A2(new_n487), .A3(new_n442), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(KEYINPUT111), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n791), .A2(new_n556), .A3(new_n611), .ZN(new_n792));
  OR2_X1    g606(.A1(new_n792), .A2(KEYINPUT112), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(KEYINPUT112), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n690), .A2(new_n483), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT49), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n676), .A2(new_n669), .A3(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n793), .A2(new_n794), .A3(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT54), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT53), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n589), .A2(new_n652), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n801), .B(new_n535), .C1(new_n629), .C2(new_n630), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n802), .A2(KEYINPUT113), .ZN(new_n803));
  INV_X1    g617(.A(new_n727), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n802), .A2(KEYINPUT113), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n803), .A2(new_n650), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n680), .A2(new_n722), .A3(new_n728), .ZN(new_n807));
  AND4_X1   g621(.A1(new_n741), .A2(new_n743), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n556), .A2(new_n679), .A3(new_n632), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n631), .A2(new_n632), .ZN(new_n810));
  OAI211_X1 g624(.A(new_n368), .B(new_n692), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n621), .A2(new_n622), .A3(new_n710), .A4(new_n489), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n605), .A2(new_n611), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n556), .A2(new_n589), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n811), .A2(new_n603), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n720), .A2(new_n646), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n808), .A2(new_n820), .A3(new_n706), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n655), .A2(new_n681), .A3(new_n724), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n623), .A2(new_n730), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n717), .A2(new_n718), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n605), .A2(KEYINPUT102), .A3(new_n712), .A4(new_n714), .ZN(new_n825));
  AOI211_X1 g639(.A(new_n823), .B(new_n671), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(KEYINPUT52), .B1(new_n822), .B2(new_n826), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n623), .A2(new_n641), .A3(new_n643), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n828), .A2(new_n686), .A3(new_n654), .ZN(new_n829));
  AOI22_X1  g643(.A1(new_n829), .A2(new_n653), .B1(new_n723), .B2(new_n680), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT52), .ZN(new_n831));
  OR2_X1    g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n824), .A2(new_n825), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n671), .A2(new_n823), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n830), .A2(new_n835), .A3(new_n831), .A4(new_n681), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n827), .A2(new_n832), .A3(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n800), .B1(new_n821), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n827), .A2(new_n836), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n693), .B1(new_n633), .B2(new_n615), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n812), .B1(new_n814), .B2(new_n815), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(new_n489), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n601), .A2(new_n535), .A3(new_n595), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT93), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n556), .A2(KEYINPUT93), .A3(new_n595), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n843), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  AOI22_X1  g662(.A1(new_n848), .A2(new_n645), .B1(new_n833), .B2(new_n711), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n706), .A2(new_n842), .A3(new_n849), .A4(new_n603), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n741), .A2(new_n743), .A3(new_n806), .A4(new_n807), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n839), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  AOI22_X1  g666(.A1(new_n838), .A2(KEYINPUT114), .B1(new_n852), .B2(KEYINPUT53), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT114), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n854), .B(new_n800), .C1(new_n821), .C2(new_n837), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n799), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n850), .A2(new_n851), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n827), .A2(new_n836), .A3(new_n832), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n857), .A2(new_n858), .A3(KEYINPUT53), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n800), .B1(new_n821), .B2(new_n839), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n859), .A2(new_n860), .A3(new_n799), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n774), .A2(new_n785), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n862), .B1(new_n774), .B2(new_n783), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT115), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n690), .A2(new_n765), .A3(new_n483), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n862), .B(KEYINPUT115), .C1(new_n774), .C2(new_n783), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n752), .A2(new_n591), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n869), .A2(new_n709), .A3(new_n746), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n869), .A2(new_n709), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT116), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(KEYINPUT50), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n873), .A2(KEYINPUT50), .ZN(new_n875));
  NOR4_X1   g689(.A1(new_n676), .A2(new_n442), .A3(new_n691), .A4(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n872), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n727), .A2(new_n691), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n869), .A2(new_n722), .A3(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n878), .A2(new_n622), .A3(new_n591), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n880), .A2(new_n669), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n881), .A2(new_n556), .A3(new_n679), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n869), .A2(new_n709), .A3(new_n876), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n884), .A2(new_n873), .A3(KEYINPUT50), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n871), .A2(new_n877), .A3(new_n883), .A4(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT51), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n884), .B(new_n874), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT117), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n883), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n863), .A2(new_n866), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n887), .B1(new_n870), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n879), .A2(new_n882), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(KEYINPUT117), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n889), .A2(new_n891), .A3(new_n893), .A4(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n872), .A2(new_n699), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n590), .B(KEYINPUT118), .ZN(new_n898));
  INV_X1    g712(.A(new_n814), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n898), .B1(new_n881), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n869), .A2(new_n878), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT48), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n738), .A2(new_n622), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n902), .A2(new_n904), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(KEYINPUT48), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n901), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n888), .A2(new_n896), .A3(new_n908), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n856), .A2(new_n861), .A3(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(G952), .A2(G953), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n798), .B1(new_n910), .B2(new_n911), .ZN(G75));
  NAND2_X1  g726(.A1(new_n859), .A2(new_n860), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n913), .A2(G210), .A3(G902), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT56), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n432), .A2(new_n433), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(new_n431), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT55), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n914), .A2(new_n915), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n918), .B1(new_n914), .B2(new_n915), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n188), .A2(G952), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(G51));
  XOR2_X1   g736(.A(new_n484), .B(KEYINPUT57), .Z(new_n923));
  AOI21_X1  g737(.A(new_n799), .B1(new_n859), .B2(new_n860), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n923), .B1(new_n861), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n925), .B1(new_n482), .B2(new_n481), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n913), .A2(G902), .A3(new_n768), .A4(new_n767), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n921), .B1(new_n926), .B2(new_n927), .ZN(G54));
  NAND4_X1  g742(.A1(new_n913), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n929));
  INV_X1    g743(.A(new_n628), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n929), .A2(new_n930), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n931), .A2(new_n932), .A3(new_n921), .ZN(G60));
  NAND2_X1  g747(.A1(new_n608), .A2(new_n609), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT119), .Z(new_n935));
  NAND2_X1  g749(.A1(G478), .A2(G902), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT59), .Z(new_n937));
  NOR2_X1   g751(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n938), .B1(new_n861), .B2(new_n924), .ZN(new_n939));
  INV_X1    g753(.A(new_n921), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n937), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n942), .B1(new_n856), .B2(new_n861), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n941), .B1(new_n943), .B2(new_n935), .ZN(G63));
  XNOR2_X1  g758(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  XNOR2_X1  g760(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT122), .ZN(new_n948));
  NAND2_X1  g762(.A1(G217), .A2(G902), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT121), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n948), .B(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n951), .B1(new_n859), .B2(new_n860), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n940), .B1(new_n952), .B2(new_n240), .ZN(new_n953));
  INV_X1    g767(.A(new_n638), .ZN(new_n954));
  AOI211_X1 g768(.A(new_n954), .B(new_n951), .C1(new_n859), .C2(new_n860), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n946), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(new_n240), .ZN(new_n957));
  INV_X1    g771(.A(new_n839), .ZN(new_n958));
  AOI21_X1  g772(.A(KEYINPUT53), .B1(new_n857), .B2(new_n958), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n821), .A2(new_n837), .A3(new_n800), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n957), .B1(new_n961), .B2(new_n951), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n952), .A2(new_n638), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n962), .A2(new_n940), .A3(new_n963), .A4(new_n945), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n956), .A2(new_n964), .ZN(G66));
  OAI21_X1  g779(.A(G953), .B1(new_n593), .B2(new_n374), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n850), .A2(KEYINPUT124), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT124), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n820), .A2(new_n968), .A3(new_n706), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n966), .B1(new_n970), .B2(G953), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n916), .B1(G898), .B2(new_n188), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n971), .B(new_n972), .ZN(G69));
  NOR2_X1   g787(.A1(new_n325), .A2(new_n326), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT125), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(new_n540), .Z(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  AND4_X1   g791(.A1(new_n368), .A2(new_n661), .A3(new_n658), .A4(new_n804), .ZN(new_n978));
  AOI22_X1  g792(.A1(new_n786), .A2(new_n787), .B1(new_n816), .B2(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n677), .A2(new_n681), .A3(new_n830), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(KEYINPUT62), .ZN(new_n981));
  INV_X1    g795(.A(new_n822), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT62), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n982), .A2(new_n983), .A3(new_n677), .ZN(new_n984));
  AND3_X1   g798(.A1(new_n979), .A2(new_n981), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n779), .A2(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n977), .B1(new_n987), .B2(G953), .ZN(new_n988));
  NAND2_X1  g802(.A1(G227), .A2(G900), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(G953), .ZN(new_n990));
  AND2_X1   g804(.A1(new_n741), .A2(new_n743), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n776), .A2(new_n904), .A3(new_n833), .ZN(new_n992));
  AND4_X1   g806(.A1(new_n788), .A2(new_n991), .A3(new_n982), .A4(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(G953), .B1(new_n779), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n651), .A2(G953), .ZN(new_n995));
  OR2_X1    g809(.A1(new_n995), .A2(KEYINPUT126), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(KEYINPUT126), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n976), .B1(new_n994), .B2(new_n998), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n988), .A2(new_n990), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n778), .A2(new_n776), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n753), .B1(new_n749), .B2(new_n751), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n745), .B1(new_n1002), .B2(KEYINPUT44), .ZN(new_n1003));
  AOI22_X1  g817(.A1(new_n1003), .A2(KEYINPUT106), .B1(new_n756), .B2(new_n755), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n777), .B1(new_n1004), .B2(new_n762), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n993), .B1(new_n1001), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1006), .A2(new_n188), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n1007), .A2(new_n997), .A3(new_n996), .ZN(new_n1008));
  OAI211_X1 g822(.A(G953), .B(new_n989), .C1(new_n1008), .C2(new_n977), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1000), .A2(new_n1009), .ZN(G72));
  INV_X1    g824(.A(KEYINPUT127), .ZN(new_n1011));
  OAI211_X1 g825(.A(new_n985), .B(new_n970), .C1(new_n1001), .C2(new_n1005), .ZN(new_n1012));
  NAND2_X1  g826(.A1(G472), .A2(G902), .ZN(new_n1013));
  XOR2_X1   g827(.A(new_n1013), .B(KEYINPUT63), .Z(new_n1014));
  NAND2_X1  g828(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n352), .A2(new_n330), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1011), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g831(.A(new_n1016), .ZN(new_n1018));
  AOI211_X1 g832(.A(KEYINPUT127), .B(new_n1018), .C1(new_n1012), .C2(new_n1014), .ZN(new_n1019));
  NOR2_X1   g833(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n838), .A2(KEYINPUT114), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n852), .A2(KEYINPUT53), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n1021), .A2(new_n855), .A3(new_n1022), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n353), .A2(new_n358), .A3(new_n664), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1023), .A2(new_n1014), .A3(new_n1024), .ZN(new_n1025));
  OAI211_X1 g839(.A(new_n970), .B(new_n993), .C1(new_n1001), .C2(new_n1005), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1026), .A2(new_n1014), .ZN(new_n1027));
  NOR3_X1   g841(.A1(new_n319), .A2(new_n303), .A3(new_n351), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n1025), .A2(new_n940), .A3(new_n1029), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n1020), .A2(new_n1030), .ZN(G57));
endmodule


