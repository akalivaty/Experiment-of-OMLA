

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591;

  XNOR2_X2 U326 ( .A(n478), .B(KEYINPUT121), .ZN(n479) );
  NAND2_X2 U327 ( .A1(n474), .A2(n473), .ZN(n475) );
  XNOR2_X2 U328 ( .A(n476), .B(n475), .ZN(n544) );
  XNOR2_X1 U329 ( .A(KEYINPUT102), .B(n460), .ZN(n504) );
  XOR2_X2 U330 ( .A(n400), .B(n399), .Z(n464) );
  XOR2_X1 U331 ( .A(G36GAT), .B(G190GAT), .Z(n418) );
  XNOR2_X1 U332 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U333 ( .A(n437), .B(n436), .ZN(n575) );
  XOR2_X1 U334 ( .A(G218GAT), .B(G106GAT), .Z(n294) );
  INV_X1 U335 ( .A(KEYINPUT98), .ZN(n406) );
  XNOR2_X1 U336 ( .A(n406), .B(KEYINPUT25), .ZN(n407) );
  XNOR2_X1 U337 ( .A(n408), .B(n407), .ZN(n411) );
  XNOR2_X1 U338 ( .A(n391), .B(n390), .ZN(n393) );
  XNOR2_X1 U339 ( .A(n424), .B(n294), .ZN(n425) );
  XNOR2_X1 U340 ( .A(n426), .B(n425), .ZN(n428) );
  XOR2_X1 U341 ( .A(KEYINPUT36), .B(n575), .Z(n588) );
  INV_X1 U342 ( .A(KEYINPUT124), .ZN(n484) );
  XNOR2_X1 U343 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U344 ( .A(n461), .B(G43GAT), .ZN(n462) );
  XNOR2_X1 U345 ( .A(n487), .B(n486), .ZN(G1352GAT) );
  XNOR2_X1 U346 ( .A(n463), .B(n462), .ZN(G1330GAT) );
  XOR2_X1 U347 ( .A(G190GAT), .B(G99GAT), .Z(n296) );
  XNOR2_X1 U348 ( .A(G43GAT), .B(G134GAT), .ZN(n295) );
  XNOR2_X1 U349 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U350 ( .A(G127GAT), .B(KEYINPUT83), .Z(n298) );
  XNOR2_X1 U351 ( .A(G120GAT), .B(KEYINPUT84), .ZN(n297) );
  XNOR2_X1 U352 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U353 ( .A(n300), .B(n299), .Z(n305) );
  XOR2_X1 U354 ( .A(G183GAT), .B(G176GAT), .Z(n302) );
  NAND2_X1 U355 ( .A1(G227GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U356 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U357 ( .A(KEYINPUT20), .B(n303), .ZN(n304) );
  XNOR2_X1 U358 ( .A(n305), .B(n304), .ZN(n309) );
  XOR2_X1 U359 ( .A(KEYINPUT85), .B(G71GAT), .Z(n307) );
  XNOR2_X1 U360 ( .A(G15GAT), .B(KEYINPUT65), .ZN(n306) );
  XNOR2_X1 U361 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U362 ( .A(n309), .B(n308), .Z(n315) );
  XOR2_X1 U363 ( .A(KEYINPUT82), .B(KEYINPUT0), .Z(n311) );
  XNOR2_X1 U364 ( .A(G113GAT), .B(KEYINPUT81), .ZN(n310) );
  XNOR2_X1 U365 ( .A(n311), .B(n310), .ZN(n354) );
  XOR2_X1 U366 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n313) );
  XNOR2_X1 U367 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n312) );
  XNOR2_X1 U368 ( .A(n313), .B(n312), .ZN(n389) );
  XNOR2_X1 U369 ( .A(n354), .B(n389), .ZN(n314) );
  XNOR2_X1 U370 ( .A(n315), .B(n314), .ZN(n564) );
  XOR2_X1 U371 ( .A(G106GAT), .B(G78GAT), .Z(n377) );
  XOR2_X1 U372 ( .A(G120GAT), .B(G148GAT), .Z(n353) );
  XNOR2_X1 U373 ( .A(n377), .B(n353), .ZN(n328) );
  XOR2_X1 U374 ( .A(G99GAT), .B(G85GAT), .Z(n429) );
  XOR2_X1 U375 ( .A(KEYINPUT32), .B(KEYINPUT72), .Z(n317) );
  XNOR2_X1 U376 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(n316) );
  XNOR2_X1 U377 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U378 ( .A(n429), .B(n318), .Z(n320) );
  NAND2_X1 U379 ( .A1(G230GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U380 ( .A(n320), .B(n319), .ZN(n326) );
  XOR2_X1 U381 ( .A(G57GAT), .B(KEYINPUT13), .Z(n322) );
  XNOR2_X1 U382 ( .A(G71GAT), .B(KEYINPUT71), .ZN(n321) );
  XNOR2_X1 U383 ( .A(n322), .B(n321), .ZN(n445) );
  XOR2_X1 U384 ( .A(G64GAT), .B(G92GAT), .Z(n324) );
  XNOR2_X1 U385 ( .A(G176GAT), .B(G204GAT), .ZN(n323) );
  XNOR2_X1 U386 ( .A(n324), .B(n323), .ZN(n387) );
  XOR2_X1 U387 ( .A(n445), .B(n387), .Z(n325) );
  XNOR2_X1 U388 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U389 ( .A(n328), .B(n327), .Z(n580) );
  XOR2_X1 U390 ( .A(KEYINPUT29), .B(KEYINPUT68), .Z(n330) );
  XNOR2_X1 U391 ( .A(G1GAT), .B(KEYINPUT69), .ZN(n329) );
  XNOR2_X1 U392 ( .A(n330), .B(n329), .ZN(n338) );
  NAND2_X1 U393 ( .A1(G229GAT), .A2(G233GAT), .ZN(n336) );
  XOR2_X1 U394 ( .A(G197GAT), .B(G113GAT), .Z(n332) );
  XNOR2_X1 U395 ( .A(G169GAT), .B(G50GAT), .ZN(n331) );
  XNOR2_X1 U396 ( .A(n332), .B(n331), .ZN(n334) );
  XOR2_X1 U397 ( .A(G29GAT), .B(G36GAT), .Z(n333) );
  XNOR2_X1 U398 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U399 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U400 ( .A(n338), .B(n337), .ZN(n346) );
  XNOR2_X1 U401 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n339) );
  XNOR2_X1 U402 ( .A(n339), .B(KEYINPUT7), .ZN(n430) );
  XOR2_X1 U403 ( .A(G8GAT), .B(KEYINPUT30), .Z(n341) );
  XNOR2_X1 U404 ( .A(G141GAT), .B(KEYINPUT70), .ZN(n340) );
  XNOR2_X1 U405 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U406 ( .A(n430), .B(n342), .ZN(n344) );
  XOR2_X1 U407 ( .A(G15GAT), .B(G22GAT), .Z(n343) );
  XOR2_X1 U408 ( .A(KEYINPUT67), .B(n343), .Z(n453) );
  XOR2_X1 U409 ( .A(n344), .B(n453), .Z(n345) );
  XNOR2_X1 U410 ( .A(n346), .B(n345), .ZN(n565) );
  INV_X1 U411 ( .A(n565), .ZN(n507) );
  NOR2_X1 U412 ( .A1(n580), .A2(n507), .ZN(n492) );
  XOR2_X1 U413 ( .A(KEYINPUT93), .B(KEYINPUT4), .Z(n348) );
  XNOR2_X1 U414 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n347) );
  XOR2_X1 U415 ( .A(n348), .B(n347), .Z(n349) );
  XOR2_X1 U416 ( .A(G1GAT), .B(G127GAT), .Z(n441) );
  XNOR2_X1 U417 ( .A(n349), .B(n441), .ZN(n351) );
  XNOR2_X1 U418 ( .A(G85GAT), .B(G57GAT), .ZN(n350) );
  XNOR2_X1 U419 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U420 ( .A(G29GAT), .B(G134GAT), .Z(n427) );
  XOR2_X1 U421 ( .A(n352), .B(n427), .Z(n356) );
  XNOR2_X1 U422 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U423 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U424 ( .A(KEYINPUT5), .B(KEYINPUT91), .Z(n358) );
  NAND2_X1 U425 ( .A1(G225GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U426 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U427 ( .A(n360), .B(n359), .Z(n366) );
  XNOR2_X1 U428 ( .A(G155GAT), .B(KEYINPUT89), .ZN(n361) );
  XNOR2_X1 U429 ( .A(n361), .B(KEYINPUT2), .ZN(n362) );
  XOR2_X1 U430 ( .A(n362), .B(KEYINPUT3), .Z(n364) );
  XNOR2_X1 U431 ( .A(G141GAT), .B(G162GAT), .ZN(n363) );
  XNOR2_X1 U432 ( .A(n364), .B(n363), .ZN(n370) );
  XNOR2_X1 U433 ( .A(n370), .B(KEYINPUT92), .ZN(n365) );
  XNOR2_X1 U434 ( .A(n366), .B(n365), .ZN(n412) );
  XOR2_X2 U435 ( .A(KEYINPUT94), .B(n412), .Z(n546) );
  XOR2_X1 U436 ( .A(KEYINPUT87), .B(G218GAT), .Z(n368) );
  XNOR2_X1 U437 ( .A(KEYINPUT21), .B(KEYINPUT88), .ZN(n367) );
  XNOR2_X1 U438 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U439 ( .A(n369), .B(G197GAT), .Z(n391) );
  XNOR2_X1 U440 ( .A(n391), .B(n370), .ZN(n384) );
  XOR2_X1 U441 ( .A(G148GAT), .B(G204GAT), .Z(n372) );
  XNOR2_X1 U442 ( .A(KEYINPUT86), .B(KEYINPUT90), .ZN(n371) );
  XNOR2_X1 U443 ( .A(n372), .B(n371), .ZN(n376) );
  XOR2_X1 U444 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n374) );
  XNOR2_X1 U445 ( .A(G22GAT), .B(KEYINPUT23), .ZN(n373) );
  XNOR2_X1 U446 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U447 ( .A(n376), .B(n375), .Z(n382) );
  XOR2_X1 U448 ( .A(G50GAT), .B(KEYINPUT73), .Z(n419) );
  XOR2_X1 U449 ( .A(G211GAT), .B(n377), .Z(n379) );
  NAND2_X1 U450 ( .A1(G228GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U451 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U452 ( .A(n419), .B(n380), .ZN(n381) );
  XNOR2_X1 U453 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U454 ( .A(n384), .B(n383), .ZN(n561) );
  XOR2_X1 U455 ( .A(n561), .B(KEYINPUT28), .Z(n526) );
  XOR2_X1 U456 ( .A(KEYINPUT76), .B(G211GAT), .Z(n386) );
  XNOR2_X1 U457 ( .A(G8GAT), .B(G183GAT), .ZN(n385) );
  XNOR2_X1 U458 ( .A(n386), .B(n385), .ZN(n452) );
  XNOR2_X1 U459 ( .A(n387), .B(n452), .ZN(n400) );
  XOR2_X1 U460 ( .A(KEYINPUT96), .B(KEYINPUT95), .Z(n388) );
  INV_X1 U461 ( .A(n393), .ZN(n392) );
  NAND2_X1 U462 ( .A1(n418), .A2(n392), .ZN(n396) );
  INV_X1 U463 ( .A(n418), .ZN(n394) );
  NAND2_X1 U464 ( .A1(n394), .A2(n393), .ZN(n395) );
  NAND2_X1 U465 ( .A1(n396), .A2(n395), .ZN(n398) );
  NAND2_X1 U466 ( .A1(G226GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U467 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U468 ( .A(n464), .B(KEYINPUT27), .ZN(n410) );
  INV_X1 U469 ( .A(n410), .ZN(n401) );
  NAND2_X1 U470 ( .A1(n526), .A2(n401), .ZN(n402) );
  NOR2_X1 U471 ( .A1(n546), .A2(n402), .ZN(n530) );
  XNOR2_X1 U472 ( .A(KEYINPUT97), .B(n530), .ZN(n404) );
  INV_X1 U473 ( .A(n564), .ZN(n403) );
  NOR2_X1 U474 ( .A1(n404), .A2(n403), .ZN(n415) );
  NOR2_X1 U475 ( .A1(n564), .A2(n464), .ZN(n405) );
  NOR2_X1 U476 ( .A1(n405), .A2(n561), .ZN(n408) );
  NAND2_X1 U477 ( .A1(n561), .A2(n564), .ZN(n409) );
  XNOR2_X1 U478 ( .A(n409), .B(KEYINPUT26), .ZN(n481) );
  NOR2_X1 U479 ( .A1(n481), .A2(n410), .ZN(n545) );
  NOR2_X1 U480 ( .A1(n411), .A2(n545), .ZN(n413) );
  NOR2_X1 U481 ( .A1(n413), .A2(n412), .ZN(n414) );
  NOR2_X1 U482 ( .A1(n415), .A2(n414), .ZN(n417) );
  INV_X1 U483 ( .A(KEYINPUT99), .ZN(n416) );
  XNOR2_X1 U484 ( .A(n417), .B(n416), .ZN(n491) );
  XOR2_X1 U485 ( .A(KEYINPUT64), .B(n418), .Z(n421) );
  XNOR2_X1 U486 ( .A(G162GAT), .B(n419), .ZN(n420) );
  XNOR2_X1 U487 ( .A(n421), .B(n420), .ZN(n426) );
  XOR2_X1 U488 ( .A(KEYINPUT75), .B(KEYINPUT9), .Z(n423) );
  XNOR2_X1 U489 ( .A(G92GAT), .B(KEYINPUT74), .ZN(n422) );
  XNOR2_X1 U490 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U491 ( .A(n428), .B(n427), .Z(n432) );
  XNOR2_X1 U492 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U493 ( .A(n432), .B(n431), .ZN(n437) );
  XOR2_X1 U494 ( .A(KEYINPUT66), .B(KEYINPUT11), .Z(n434) );
  NAND2_X1 U495 ( .A1(G232GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U496 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U497 ( .A(KEYINPUT10), .B(n435), .Z(n436) );
  XOR2_X1 U498 ( .A(KEYINPUT77), .B(G64GAT), .Z(n439) );
  XNOR2_X1 U499 ( .A(G155GAT), .B(G78GAT), .ZN(n438) );
  XNOR2_X1 U500 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U501 ( .A(n441), .B(n440), .Z(n443) );
  NAND2_X1 U502 ( .A1(G231GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U503 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U504 ( .A(n444), .B(KEYINPUT12), .Z(n447) );
  XNOR2_X1 U505 ( .A(n445), .B(KEYINPUT80), .ZN(n446) );
  XNOR2_X1 U506 ( .A(n447), .B(n446), .ZN(n451) );
  XOR2_X1 U507 ( .A(KEYINPUT79), .B(KEYINPUT15), .Z(n449) );
  XNOR2_X1 U508 ( .A(KEYINPUT78), .B(KEYINPUT14), .ZN(n448) );
  XNOR2_X1 U509 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U510 ( .A(n451), .B(n450), .Z(n455) );
  XNOR2_X1 U511 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U512 ( .A(n455), .B(n454), .ZN(n488) );
  INV_X1 U513 ( .A(n488), .ZN(n584) );
  OR2_X1 U514 ( .A1(n588), .A2(n584), .ZN(n456) );
  OR2_X1 U515 ( .A1(n491), .A2(n456), .ZN(n457) );
  XNOR2_X1 U516 ( .A(n457), .B(KEYINPUT101), .ZN(n458) );
  XOR2_X1 U517 ( .A(KEYINPUT37), .B(n458), .Z(n517) );
  NAND2_X1 U518 ( .A1(n492), .A2(n517), .ZN(n459) );
  XNOR2_X1 U519 ( .A(n459), .B(KEYINPUT38), .ZN(n460) );
  NOR2_X1 U520 ( .A1(n564), .A2(n504), .ZN(n463) );
  INV_X1 U521 ( .A(KEYINPUT40), .ZN(n461) );
  XOR2_X1 U522 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n483) );
  XOR2_X1 U523 ( .A(KEYINPUT120), .B(n464), .Z(n477) );
  XNOR2_X1 U524 ( .A(KEYINPUT112), .B(KEYINPUT48), .ZN(n476) );
  XOR2_X1 U525 ( .A(KEYINPUT41), .B(n580), .Z(n551) );
  NAND2_X1 U526 ( .A1(n565), .A2(n551), .ZN(n465) );
  XNOR2_X1 U527 ( .A(n465), .B(KEYINPUT46), .ZN(n466) );
  XNOR2_X1 U528 ( .A(n488), .B(KEYINPUT110), .ZN(n573) );
  NAND2_X1 U529 ( .A1(n466), .A2(n573), .ZN(n467) );
  NOR2_X1 U530 ( .A1(n575), .A2(n467), .ZN(n468) );
  XNOR2_X1 U531 ( .A(n468), .B(KEYINPUT47), .ZN(n474) );
  NOR2_X1 U532 ( .A1(n488), .A2(n588), .ZN(n470) );
  XNOR2_X1 U533 ( .A(KEYINPUT45), .B(KEYINPUT111), .ZN(n469) );
  XNOR2_X1 U534 ( .A(n470), .B(n469), .ZN(n471) );
  NOR2_X1 U535 ( .A1(n580), .A2(n471), .ZN(n472) );
  NAND2_X1 U536 ( .A1(n472), .A2(n507), .ZN(n473) );
  NAND2_X1 U537 ( .A1(n477), .A2(n544), .ZN(n478) );
  XNOR2_X1 U538 ( .A(KEYINPUT54), .B(n479), .ZN(n480) );
  NAND2_X1 U539 ( .A1(n480), .A2(n546), .ZN(n560) );
  NOR2_X1 U540 ( .A1(n560), .A2(n481), .ZN(n586) );
  NAND2_X1 U541 ( .A1(n586), .A2(n565), .ZN(n482) );
  XNOR2_X1 U542 ( .A(n483), .B(n482), .ZN(n487) );
  XNOR2_X1 U543 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n485) );
  NOR2_X1 U544 ( .A1(n488), .A2(n575), .ZN(n489) );
  XOR2_X1 U545 ( .A(KEYINPUT16), .B(n489), .Z(n490) );
  NOR2_X1 U546 ( .A1(n491), .A2(n490), .ZN(n508) );
  NAND2_X1 U547 ( .A1(n492), .A2(n508), .ZN(n499) );
  NOR2_X1 U548 ( .A1(n546), .A2(n499), .ZN(n494) );
  XNOR2_X1 U549 ( .A(KEYINPUT34), .B(KEYINPUT100), .ZN(n493) );
  XNOR2_X1 U550 ( .A(n494), .B(n493), .ZN(n495) );
  XOR2_X1 U551 ( .A(G1GAT), .B(n495), .Z(G1324GAT) );
  NOR2_X1 U552 ( .A1(n464), .A2(n499), .ZN(n496) );
  XOR2_X1 U553 ( .A(G8GAT), .B(n496), .Z(G1325GAT) );
  NOR2_X1 U554 ( .A1(n564), .A2(n499), .ZN(n498) );
  XNOR2_X1 U555 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n497) );
  XNOR2_X1 U556 ( .A(n498), .B(n497), .ZN(G1326GAT) );
  NOR2_X1 U557 ( .A1(n526), .A2(n499), .ZN(n500) );
  XOR2_X1 U558 ( .A(G22GAT), .B(n500), .Z(G1327GAT) );
  NOR2_X1 U559 ( .A1(n504), .A2(n546), .ZN(n502) );
  XNOR2_X1 U560 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n501) );
  XNOR2_X1 U561 ( .A(n502), .B(n501), .ZN(G1328GAT) );
  NOR2_X1 U562 ( .A1(n504), .A2(n464), .ZN(n503) );
  XOR2_X1 U563 ( .A(G36GAT), .B(n503), .Z(G1329GAT) );
  NOR2_X1 U564 ( .A1(n526), .A2(n504), .ZN(n506) );
  XNOR2_X1 U565 ( .A(G50GAT), .B(KEYINPUT103), .ZN(n505) );
  XNOR2_X1 U566 ( .A(n506), .B(n505), .ZN(G1331GAT) );
  XNOR2_X1 U567 ( .A(n551), .B(KEYINPUT104), .ZN(n568) );
  AND2_X1 U568 ( .A1(n507), .A2(n568), .ZN(n518) );
  NAND2_X1 U569 ( .A1(n518), .A2(n508), .ZN(n514) );
  NOR2_X1 U570 ( .A1(n546), .A2(n514), .ZN(n509) );
  XOR2_X1 U571 ( .A(G57GAT), .B(n509), .Z(n510) );
  XNOR2_X1 U572 ( .A(KEYINPUT42), .B(n510), .ZN(G1332GAT) );
  NOR2_X1 U573 ( .A1(n464), .A2(n514), .ZN(n511) );
  XOR2_X1 U574 ( .A(G64GAT), .B(n511), .Z(G1333GAT) );
  NOR2_X1 U575 ( .A1(n564), .A2(n514), .ZN(n513) );
  XNOR2_X1 U576 ( .A(G71GAT), .B(KEYINPUT105), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n513), .B(n512), .ZN(G1334GAT) );
  NOR2_X1 U578 ( .A1(n526), .A2(n514), .ZN(n516) );
  XNOR2_X1 U579 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n516), .B(n515), .ZN(G1335GAT) );
  XNOR2_X1 U581 ( .A(G85GAT), .B(KEYINPUT107), .ZN(n521) );
  NAND2_X1 U582 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U583 ( .A(n519), .B(KEYINPUT106), .ZN(n525) );
  NOR2_X1 U584 ( .A1(n546), .A2(n525), .ZN(n520) );
  XNOR2_X1 U585 ( .A(n521), .B(n520), .ZN(G1336GAT) );
  NOR2_X1 U586 ( .A1(n525), .A2(n464), .ZN(n522) );
  XOR2_X1 U587 ( .A(KEYINPUT108), .B(n522), .Z(n523) );
  XNOR2_X1 U588 ( .A(G92GAT), .B(n523), .ZN(G1337GAT) );
  NOR2_X1 U589 ( .A1(n564), .A2(n525), .ZN(n524) );
  XOR2_X1 U590 ( .A(G99GAT), .B(n524), .Z(G1338GAT) );
  XNOR2_X1 U591 ( .A(KEYINPUT44), .B(KEYINPUT109), .ZN(n528) );
  NOR2_X1 U592 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U594 ( .A(G106GAT), .B(n529), .ZN(G1339GAT) );
  NAND2_X1 U595 ( .A1(n544), .A2(n530), .ZN(n531) );
  NOR2_X1 U596 ( .A1(n564), .A2(n531), .ZN(n540) );
  NAND2_X1 U597 ( .A1(n540), .A2(n565), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n532), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT113), .B(KEYINPUT49), .Z(n534) );
  NAND2_X1 U600 ( .A1(n540), .A2(n568), .ZN(n533) );
  XNOR2_X1 U601 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U602 ( .A(G120GAT), .B(n535), .Z(G1341GAT) );
  INV_X1 U603 ( .A(n540), .ZN(n536) );
  NOR2_X1 U604 ( .A1(n573), .A2(n536), .ZN(n538) );
  XNOR2_X1 U605 ( .A(KEYINPUT50), .B(KEYINPUT114), .ZN(n537) );
  XNOR2_X1 U606 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U607 ( .A(G127GAT), .B(n539), .Z(G1342GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n542) );
  NAND2_X1 U609 ( .A1(n540), .A2(n575), .ZN(n541) );
  XNOR2_X1 U610 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U611 ( .A(G134GAT), .B(n543), .Z(G1343GAT) );
  XOR2_X1 U612 ( .A(G141GAT), .B(KEYINPUT117), .Z(n550) );
  NAND2_X1 U613 ( .A1(n545), .A2(n544), .ZN(n547) );
  NOR2_X1 U614 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n548), .B(KEYINPUT116), .ZN(n557) );
  NAND2_X1 U616 ( .A1(n565), .A2(n557), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(G1344GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n553) );
  NAND2_X1 U619 ( .A1(n551), .A2(n557), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(n554), .ZN(G1345GAT) );
  NAND2_X1 U622 ( .A1(n557), .A2(n584), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n555), .B(KEYINPUT118), .ZN(n556) );
  XNOR2_X1 U624 ( .A(G155GAT), .B(n556), .ZN(G1346GAT) );
  XOR2_X1 U625 ( .A(G162GAT), .B(KEYINPUT119), .Z(n559) );
  NAND2_X1 U626 ( .A1(n557), .A2(n575), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(G1347GAT) );
  NOR2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(KEYINPUT55), .ZN(n563) );
  NOR2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n576) );
  NAND2_X1 U631 ( .A1(n576), .A2(n565), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(KEYINPUT122), .ZN(n567) );
  XNOR2_X1 U633 ( .A(G169GAT), .B(n567), .ZN(G1348GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n570) );
  NAND2_X1 U635 ( .A1(n576), .A2(n568), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(G176GAT), .B(n571), .ZN(G1349GAT) );
  INV_X1 U638 ( .A(n576), .ZN(n572) );
  NOR2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U640 ( .A(G183GAT), .B(n574), .Z(G1350GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n578) );
  NAND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(G190GAT), .B(n579), .ZN(G1351GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n582) );
  NAND2_X1 U646 ( .A1(n586), .A2(n580), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(G204GAT), .B(n583), .ZN(G1353GAT) );
  NAND2_X1 U649 ( .A1(n586), .A2(n584), .ZN(n585) );
  XNOR2_X1 U650 ( .A(G211GAT), .B(n585), .ZN(G1354GAT) );
  INV_X1 U651 ( .A(n586), .ZN(n587) );
  NOR2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n590) );
  XNOR2_X1 U653 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

