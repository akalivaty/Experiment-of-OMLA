//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 1 1 1 1 1 0 0 0 0 1 1 1 0 1 1 0 0 0 1 0 1 1 0 0 0 0 0 1 0 1 1 1 0 1 1 0 0 1 0 1 1 0 1 1 0 1 0 1 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:28 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004;
  INV_X1    g000(.A(KEYINPUT69), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(KEYINPUT65), .ZN(new_n190));
  AND2_X1   g004(.A1(KEYINPUT64), .A2(G146), .ZN(new_n191));
  NOR2_X1   g005(.A1(KEYINPUT64), .A2(G146), .ZN(new_n192));
  OAI21_X1  g006(.A(G143), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(new_n189), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n190), .B1(new_n195), .B2(KEYINPUT65), .ZN(new_n196));
  INV_X1    g010(.A(G128), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(KEYINPUT1), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n193), .A2(KEYINPUT1), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G128), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n188), .A2(G143), .ZN(new_n201));
  XNOR2_X1  g015(.A(KEYINPUT64), .B(G146), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n201), .B1(new_n202), .B2(G143), .ZN(new_n203));
  AOI22_X1  g017(.A1(new_n196), .A2(new_n198), .B1(new_n200), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G137), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G134), .ZN(new_n206));
  NAND2_X1  g020(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n207), .B1(new_n205), .B2(G134), .ZN(new_n208));
  NOR2_X1   g022(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n206), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G131), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT67), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT11), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n212), .B1(new_n206), .B2(new_n213), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n205), .A2(KEYINPUT67), .A3(KEYINPUT11), .A4(G134), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n210), .A2(new_n211), .A3(new_n214), .A4(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G134), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G137), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n206), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G131), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n216), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n187), .B1(new_n204), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(KEYINPUT68), .A2(G131), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n214), .A2(new_n215), .ZN(new_n225));
  AOI22_X1  g039(.A1(new_n217), .A2(G137), .B1(KEYINPUT66), .B2(KEYINPUT11), .ZN(new_n226));
  INV_X1    g040(.A(new_n209), .ZN(new_n227));
  AOI22_X1  g041(.A1(new_n226), .A2(new_n227), .B1(G134), .B2(new_n205), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n224), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n210), .A2(new_n223), .A3(new_n214), .A4(new_n215), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(KEYINPUT0), .A2(G128), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n196), .A2(new_n233), .ZN(new_n234));
  OR2_X1    g048(.A1(KEYINPUT0), .A2(G128), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n203), .A2(new_n232), .A3(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n231), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n190), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n189), .B1(new_n202), .B2(G143), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT65), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n238), .B(new_n198), .C1(new_n239), .C2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT1), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n242), .B1(new_n202), .B2(G143), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n203), .B1(new_n243), .B2(new_n197), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n245), .A2(KEYINPUT69), .A3(new_n220), .A4(new_n216), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n222), .A2(new_n237), .A3(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT30), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XOR2_X1   g063(.A(KEYINPUT2), .B(G113), .Z(new_n250));
  XNOR2_X1  g064(.A(G116), .B(G119), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G119), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G116), .ZN(new_n254));
  INV_X1    g068(.A(G116), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G119), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT2), .B(G113), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n252), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n216), .A2(KEYINPUT70), .A3(new_n220), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n245), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(KEYINPUT70), .B1(new_n216), .B2(new_n220), .ZN(new_n263));
  OAI211_X1 g077(.A(KEYINPUT30), .B(new_n237), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n249), .A2(new_n260), .A3(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT71), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n260), .B(new_n266), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n267), .B(new_n237), .C1(new_n262), .C2(new_n263), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n269), .B(G101), .ZN(new_n270));
  INV_X1    g084(.A(G210), .ZN(new_n271));
  NOR3_X1   g085(.A1(new_n271), .A2(G237), .A3(G953), .ZN(new_n272));
  XOR2_X1   g086(.A(new_n270), .B(new_n272), .Z(new_n273));
  NAND3_X1  g087(.A1(new_n265), .A2(new_n268), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT31), .ZN(new_n275));
  INV_X1    g089(.A(new_n273), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT28), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n268), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT72), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n268), .A2(KEYINPUT72), .A3(new_n277), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n247), .A2(new_n260), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n277), .B1(new_n283), .B2(new_n268), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n276), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT31), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n265), .A2(new_n286), .A3(new_n268), .A4(new_n273), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n275), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G472), .ZN(new_n289));
  INV_X1    g103(.A(G902), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT32), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n265), .A2(new_n268), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(new_n276), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n283), .A2(new_n268), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(KEYINPUT28), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n268), .A2(KEYINPUT72), .A3(new_n277), .ZN(new_n298));
  AOI21_X1  g112(.A(KEYINPUT72), .B1(new_n268), .B2(new_n277), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n297), .A2(new_n300), .A3(new_n273), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT29), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n295), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT73), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n304), .B1(new_n298), .B2(new_n299), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n280), .A2(KEYINPUT73), .A3(new_n281), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n237), .B1(new_n262), .B2(new_n263), .ZN(new_n308));
  INV_X1    g122(.A(new_n267), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n277), .B1(new_n310), .B2(new_n268), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n307), .A2(KEYINPUT29), .A3(new_n273), .A4(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n303), .A2(new_n313), .A3(new_n290), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G472), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n288), .A2(KEYINPUT32), .A3(new_n289), .A4(new_n290), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n293), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G953), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n318), .A2(G221), .A3(G234), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n319), .B(KEYINPUT22), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n320), .B(new_n205), .ZN(new_n321));
  INV_X1    g135(.A(G125), .ZN(new_n322));
  OR3_X1    g136(.A1(new_n322), .A2(KEYINPUT16), .A3(G140), .ZN(new_n323));
  XOR2_X1   g137(.A(G125), .B(G140), .Z(new_n324));
  INV_X1    g138(.A(KEYINPUT16), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n323), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n188), .ZN(new_n327));
  OAI211_X1 g141(.A(G146), .B(new_n323), .C1(new_n324), .C2(new_n325), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT23), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n330), .B1(new_n253), .B2(G128), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n197), .A2(KEYINPUT23), .A3(G119), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n331), .B(new_n332), .C1(G119), .C2(new_n197), .ZN(new_n333));
  XNOR2_X1  g147(.A(G119), .B(G128), .ZN(new_n334));
  XOR2_X1   g148(.A(KEYINPUT24), .B(G110), .Z(new_n335));
  AOI22_X1  g149(.A1(new_n333), .A2(G110), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n329), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(G125), .B(G140), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n202), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n339), .B(KEYINPUT74), .ZN(new_n340));
  OAI22_X1  g154(.A1(new_n333), .A2(G110), .B1(new_n334), .B2(new_n335), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(new_n328), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n337), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n321), .B1(new_n343), .B2(KEYINPUT75), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(KEYINPUT75), .ZN(new_n345));
  XOR2_X1   g159(.A(new_n344), .B(new_n345), .Z(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  OAI211_X1 g161(.A(KEYINPUT76), .B(KEYINPUT25), .C1(new_n347), .C2(G902), .ZN(new_n348));
  INV_X1    g162(.A(G217), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n349), .B1(G234), .B2(new_n290), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT76), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT25), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n351), .A2(new_n352), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n346), .A2(new_n290), .A3(new_n354), .A4(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n348), .A2(new_n350), .A3(new_n356), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n350), .A2(G902), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n346), .A2(new_n358), .ZN(new_n359));
  AND2_X1   g173(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n317), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G237), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n363), .A2(new_n318), .A3(G214), .ZN(new_n364));
  INV_X1    g178(.A(G143), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n364), .B(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G131), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n364), .B(G143), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n211), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT17), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n367), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT86), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n366), .A2(KEYINPUT17), .A3(G131), .ZN(new_n374));
  AND3_X1   g188(.A1(new_n374), .A2(new_n327), .A3(new_n328), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n367), .A2(new_n369), .A3(KEYINPUT86), .A4(new_n370), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n373), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n324), .A2(G146), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT18), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n366), .B1(new_n379), .B2(new_n211), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n368), .A2(KEYINPUT18), .A3(G131), .ZN(new_n381));
  AOI22_X1  g195(.A1(new_n340), .A2(new_n378), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(G113), .B(G122), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n384), .B(G104), .ZN(new_n385));
  XOR2_X1   g199(.A(new_n385), .B(KEYINPUT85), .Z(new_n386));
  NAND3_X1  g200(.A1(new_n377), .A2(new_n383), .A3(new_n386), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n324), .B(KEYINPUT19), .ZN(new_n388));
  INV_X1    g202(.A(new_n202), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n328), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n390), .B1(new_n367), .B2(new_n369), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n385), .B1(new_n391), .B2(new_n382), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n387), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G475), .ZN(new_n394));
  AND4_X1   g208(.A1(KEYINPUT20), .A2(new_n393), .A3(new_n394), .A4(new_n290), .ZN(new_n395));
  AOI21_X1  g209(.A(G475), .B1(new_n387), .B2(new_n392), .ZN(new_n396));
  AOI21_X1  g210(.A(KEYINPUT20), .B1(new_n396), .B2(new_n290), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  XOR2_X1   g212(.A(KEYINPUT87), .B(G475), .Z(new_n399));
  INV_X1    g213(.A(new_n387), .ZN(new_n400));
  INV_X1    g214(.A(new_n385), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n377), .A2(new_n383), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n401), .B1(new_n402), .B2(KEYINPUT88), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT88), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n377), .A2(new_n404), .A3(new_n383), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n400), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n399), .B1(new_n406), .B2(G902), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n398), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n197), .A2(G143), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT89), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n409), .B(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT90), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n365), .A2(G128), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n412), .B1(new_n411), .B2(new_n413), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n217), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n411), .A2(new_n413), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(KEYINPUT90), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n419), .A2(G134), .A3(new_n414), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n255), .A2(KEYINPUT14), .A3(G122), .ZN(new_n421));
  XNOR2_X1  g235(.A(G116), .B(G122), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT14), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n421), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(KEYINPUT78), .B(G107), .ZN(new_n425));
  AOI22_X1  g239(.A1(new_n424), .A2(G107), .B1(new_n425), .B2(new_n422), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n417), .A2(new_n420), .A3(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT13), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n411), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n418), .A2(new_n429), .A3(G134), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n425), .B(new_n422), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n411), .B(new_n413), .C1(new_n428), .C2(new_n217), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n427), .A2(new_n433), .ZN(new_n434));
  XOR2_X1   g248(.A(KEYINPUT9), .B(G234), .Z(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  NOR3_X1   g250(.A1(new_n436), .A2(new_n349), .A3(G953), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n427), .A2(new_n433), .A3(new_n437), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT91), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n441), .A2(new_n442), .A3(new_n290), .ZN(new_n443));
  INV_X1    g257(.A(G478), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n444), .A2(KEYINPUT15), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n445), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n441), .A2(new_n442), .A3(new_n290), .A4(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  OR2_X1    g263(.A1(new_n408), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n318), .A2(G952), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n451), .B1(G234), .B2(G237), .ZN(new_n452));
  XOR2_X1   g266(.A(KEYINPUT21), .B(G898), .Z(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  AOI211_X1 g268(.A(new_n290), .B(new_n318), .C1(G234), .C2(G237), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n452), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n450), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(G469), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT12), .ZN(new_n459));
  INV_X1    g273(.A(G104), .ZN(new_n460));
  OAI21_X1  g274(.A(KEYINPUT3), .B1(new_n460), .B2(G107), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT77), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OAI211_X1 g277(.A(KEYINPUT77), .B(KEYINPUT3), .C1(new_n460), .C2(G107), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(G101), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n460), .A2(G107), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT3), .ZN(new_n468));
  AND2_X1   g282(.A1(KEYINPUT78), .A2(G107), .ZN(new_n469));
  NOR2_X1   g283(.A1(KEYINPUT78), .A2(G107), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n468), .B(G104), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n465), .A2(new_n466), .A3(new_n467), .A4(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(G107), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(G104), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n474), .B1(new_n425), .B2(G104), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(G101), .ZN(new_n476));
  AND2_X1   g290(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n477), .A2(new_n245), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n201), .A2(KEYINPUT1), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(G128), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n240), .B1(new_n193), .B2(new_n194), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n480), .B1(new_n481), .B2(new_n190), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT81), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  OAI211_X1 g298(.A(KEYINPUT81), .B(new_n480), .C1(new_n481), .C2(new_n190), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(new_n241), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n478), .B1(new_n477), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n231), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n459), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n486), .A2(new_n477), .ZN(new_n490));
  INV_X1    g304(.A(new_n478), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(KEYINPUT12), .A3(new_n231), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT10), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  AND2_X1   g310(.A1(new_n234), .A2(new_n236), .ZN(new_n497));
  INV_X1    g311(.A(new_n464), .ZN(new_n498));
  AOI21_X1  g312(.A(KEYINPUT77), .B1(new_n474), .B2(KEYINPUT3), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n467), .B(new_n471), .C1(new_n498), .C2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT79), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n465), .A2(KEYINPUT79), .A3(new_n467), .A4(new_n471), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n466), .A2(KEYINPUT80), .ZN(new_n505));
  AOI22_X1  g319(.A1(new_n504), .A2(new_n505), .B1(KEYINPUT4), .B2(new_n472), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT4), .ZN(new_n507));
  INV_X1    g321(.A(new_n505), .ZN(new_n508));
  AOI211_X1 g322(.A(new_n507), .B(new_n508), .C1(new_n502), .C2(new_n503), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n497), .B1(new_n506), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n472), .A2(new_n476), .ZN(new_n511));
  NOR3_X1   g325(.A1(new_n204), .A2(new_n495), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n496), .A2(new_n510), .A3(new_n488), .A4(new_n513), .ZN(new_n514));
  XOR2_X1   g328(.A(G110), .B(G140), .Z(new_n515));
  AND2_X1   g329(.A1(new_n318), .A2(G227), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n515), .B(new_n516), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n494), .A2(new_n514), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n496), .A2(new_n510), .A3(new_n513), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(new_n231), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n517), .B1(new_n520), .B2(new_n514), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n458), .B(new_n290), .C1(new_n518), .C2(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n458), .A2(new_n290), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n520), .A2(new_n514), .A3(new_n517), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n496), .A2(new_n510), .A3(new_n513), .ZN(new_n526));
  AOI22_X1  g340(.A1(new_n526), .A2(new_n488), .B1(new_n489), .B2(new_n493), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n525), .B(G469), .C1(new_n527), .C2(new_n517), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n522), .A2(new_n524), .A3(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(G221), .B1(new_n436), .B2(G902), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g345(.A(G110), .B(G122), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n260), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n504), .A2(new_n505), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n472), .A2(KEYINPUT4), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n504), .A2(KEYINPUT4), .A3(new_n505), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n534), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n254), .A2(KEYINPUT5), .ZN(new_n540));
  INV_X1    g354(.A(G113), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n254), .A2(new_n256), .A3(KEYINPUT5), .ZN(new_n543));
  AOI22_X1  g357(.A1(new_n542), .A2(new_n543), .B1(new_n251), .B2(new_n250), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n477), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n533), .B1(new_n539), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n508), .B1(new_n502), .B2(new_n503), .ZN(new_n548));
  INV_X1    g362(.A(new_n536), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n538), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n260), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n551), .A2(new_n532), .A3(new_n545), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n547), .A2(new_n552), .A3(KEYINPUT6), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n245), .A2(new_n322), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n234), .A2(G125), .A3(new_n236), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(G224), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n557), .A2(G953), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n554), .A2(new_n555), .A3(new_n558), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT6), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n563), .B(new_n533), .C1(new_n539), .C2(new_n546), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n553), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(G210), .B1(G237), .B2(G902), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n566), .A2(KEYINPUT84), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT82), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n543), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n251), .A2(KEYINPUT82), .A3(KEYINPUT5), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n542), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n252), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n572), .A2(new_n472), .A3(new_n476), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n511), .A2(new_n544), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n532), .B(KEYINPUT8), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  AND2_X1   g390(.A1(new_n561), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n556), .A2(KEYINPUT7), .A3(new_n559), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT83), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT7), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n554), .A2(new_n555), .A3(new_n580), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n577), .A2(new_n578), .A3(new_n579), .A4(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n561), .A2(new_n581), .A3(new_n576), .ZN(new_n583));
  AOI211_X1 g397(.A(new_n580), .B(new_n558), .C1(new_n554), .C2(new_n555), .ZN(new_n584));
  OAI21_X1  g398(.A(KEYINPUT83), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n582), .A2(new_n585), .A3(new_n552), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n290), .ZN(new_n587));
  NOR3_X1   g401(.A1(new_n565), .A2(new_n567), .A3(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n567), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n586), .A2(new_n290), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n553), .A2(new_n562), .A3(new_n564), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(G214), .B1(G237), .B2(G902), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NOR3_X1   g409(.A1(new_n531), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n362), .A2(new_n457), .A3(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(KEYINPUT92), .B(G101), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n597), .B(new_n598), .ZN(G3));
  AOI21_X1  g413(.A(new_n289), .B1(new_n288), .B2(new_n290), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  AND2_X1   g415(.A1(new_n601), .A2(new_n291), .ZN(new_n602));
  AND2_X1   g416(.A1(new_n529), .A2(new_n530), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n602), .A2(new_n603), .A3(new_n360), .ZN(new_n604));
  INV_X1    g418(.A(new_n566), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n605), .B1(new_n565), .B2(new_n587), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n590), .A2(new_n566), .A3(new_n591), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n456), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n608), .A2(new_n609), .A3(new_n594), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n441), .A2(KEYINPUT33), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT33), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n439), .A2(new_n612), .A3(new_n440), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n611), .A2(G478), .A3(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n441), .A2(new_n444), .A3(new_n290), .ZN(new_n615));
  NAND2_X1  g429(.A1(G478), .A2(G902), .ZN(new_n616));
  AND3_X1   g430(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n408), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n610), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n604), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g434(.A(KEYINPUT34), .B(G104), .Z(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G6));
  INV_X1    g436(.A(new_n408), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n449), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n610), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n604), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT35), .B(G107), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G9));
  NOR2_X1   g442(.A1(new_n321), .A2(KEYINPUT36), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n343), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n358), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n357), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n596), .A2(new_n457), .A3(new_n602), .A4(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT93), .B(KEYINPUT37), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(G110), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n633), .B(new_n635), .ZN(G12));
  AND3_X1   g450(.A1(new_n317), .A2(new_n603), .A3(new_n632), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n565), .A2(new_n605), .A3(new_n587), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n566), .B1(new_n590), .B2(new_n591), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n594), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(G900), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n452), .B1(new_n455), .B2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  AND4_X1   g457(.A1(new_n449), .A2(new_n398), .A3(new_n407), .A4(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g459(.A(KEYINPUT94), .B1(new_n640), .B2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT94), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n608), .A2(new_n647), .A3(new_n594), .A4(new_n644), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n637), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(G128), .ZN(G30));
  XOR2_X1   g465(.A(new_n642), .B(KEYINPUT39), .Z(new_n652));
  NAND2_X1  g466(.A1(new_n603), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT96), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT40), .ZN(new_n655));
  OR2_X1    g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(new_n593), .B(KEYINPUT38), .Z(new_n657));
  INV_X1    g471(.A(KEYINPUT95), .ZN(new_n658));
  AOI22_X1  g472(.A1(new_n398), .A2(new_n407), .B1(new_n448), .B2(new_n446), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n357), .A2(new_n594), .A3(new_n631), .A4(new_n659), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n657), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n660), .A2(new_n658), .ZN(new_n662));
  INV_X1    g476(.A(new_n294), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n663), .A2(new_n276), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n310), .A2(new_n268), .A3(new_n276), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n290), .ZN(new_n666));
  OAI21_X1  g480(.A(G472), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n293), .A2(new_n316), .A3(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n661), .A2(new_n662), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n654), .A2(new_n655), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n656), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G143), .ZN(G45));
  NAND3_X1  g487(.A1(new_n408), .A2(new_n617), .A3(new_n643), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n640), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n637), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(KEYINPUT97), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(new_n188), .ZN(G48));
  OAI21_X1  g492(.A(new_n290), .B1(new_n518), .B2(new_n521), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(G469), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n680), .A2(new_n530), .A3(new_n522), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n362), .A2(new_n619), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(KEYINPUT41), .B(G113), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G15));
  NAND3_X1  g499(.A1(new_n362), .A2(new_n625), .A3(new_n682), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G116), .ZN(G18));
  AND2_X1   g501(.A1(new_n317), .A2(new_n632), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n640), .A2(new_n681), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n688), .A2(new_n457), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G119), .ZN(G21));
  AOI21_X1  g505(.A(new_n311), .B1(new_n305), .B2(new_n306), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT98), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n276), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  AOI211_X1 g508(.A(KEYINPUT98), .B(new_n311), .C1(new_n305), .C2(new_n306), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n275), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(KEYINPUT99), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT99), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n698), .B(new_n275), .C1(new_n694), .C2(new_n695), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n697), .A2(new_n287), .A3(new_n699), .ZN(new_n700));
  NOR2_X1   g514(.A1(G472), .A2(G902), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n600), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n357), .A2(KEYINPUT100), .A3(new_n359), .ZN(new_n703));
  AOI21_X1  g517(.A(KEYINPUT100), .B1(new_n357), .B2(new_n359), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  OAI211_X1 g519(.A(new_n594), .B(new_n659), .C1(new_n638), .C2(new_n639), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT101), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n608), .A2(KEYINPUT101), .A3(new_n594), .A4(new_n659), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n681), .A2(new_n456), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n702), .A2(new_n705), .A3(new_n710), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G122), .ZN(G24));
  NAND2_X1  g527(.A1(new_n700), .A2(new_n701), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n640), .A2(new_n681), .A3(new_n674), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n714), .A2(new_n601), .A3(new_n632), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G125), .ZN(G27));
  OAI21_X1  g531(.A(new_n567), .B1(new_n565), .B2(new_n587), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n590), .A2(new_n589), .A3(new_n591), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n718), .A2(new_n594), .A3(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT42), .ZN(new_n721));
  NOR4_X1   g535(.A1(new_n531), .A2(new_n720), .A3(new_n721), .A4(new_n674), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT103), .ZN(new_n723));
  OR2_X1    g537(.A1(new_n316), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n316), .A2(new_n723), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n724), .A2(new_n315), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n293), .A2(KEYINPUT104), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT104), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n291), .A2(new_n728), .A3(new_n292), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n722), .B(new_n705), .C1(new_n726), .C2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(KEYINPUT102), .A2(KEYINPUT42), .ZN(new_n732));
  OR2_X1    g546(.A1(KEYINPUT102), .A2(KEYINPUT42), .ZN(new_n733));
  INV_X1    g547(.A(new_n720), .ZN(new_n734));
  INV_X1    g548(.A(new_n674), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n734), .A2(new_n530), .A3(new_n735), .A4(new_n529), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n732), .B(new_n733), .C1(new_n361), .C2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n731), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G131), .ZN(G33));
  NOR2_X1   g553(.A1(new_n531), .A2(new_n720), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n362), .A2(new_n644), .A3(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G134), .ZN(G36));
  INV_X1    g556(.A(KEYINPUT108), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(KEYINPUT43), .ZN(new_n744));
  XOR2_X1   g558(.A(KEYINPUT108), .B(KEYINPUT43), .Z(new_n745));
  NAND3_X1  g559(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n408), .A2(new_n746), .ZN(new_n747));
  MUX2_X1   g561(.A(new_n744), .B(new_n745), .S(new_n747), .Z(new_n748));
  INV_X1    g562(.A(new_n602), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n748), .A2(new_n749), .A3(new_n632), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT44), .ZN(new_n751));
  OR2_X1    g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n750), .A2(new_n751), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n752), .A2(new_n734), .A3(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT46), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT45), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n517), .B1(new_n494), .B2(new_n514), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n514), .A2(new_n517), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n512), .B1(new_n550), .B2(new_n497), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n488), .B1(new_n759), .B2(new_n496), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n756), .B1(new_n757), .B2(new_n761), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n525), .B(KEYINPUT45), .C1(new_n527), .C2(new_n517), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(G469), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(KEYINPUT105), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT105), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n762), .A2(new_n766), .A3(new_n763), .A4(G469), .ZN(new_n767));
  AOI211_X1 g581(.A(new_n755), .B(new_n523), .C1(new_n765), .C2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n522), .ZN(new_n769));
  OAI21_X1  g583(.A(KEYINPUT106), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n765), .A2(new_n767), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n755), .B1(new_n772), .B2(new_n523), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n771), .A2(KEYINPUT46), .A3(new_n524), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT106), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n774), .A2(new_n775), .A3(new_n522), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n770), .A2(new_n773), .A3(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n777), .A2(new_n530), .A3(new_n652), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(KEYINPUT107), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT107), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n777), .A2(new_n780), .A3(new_n530), .A4(new_n652), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n754), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(new_n205), .ZN(G39));
  NAND2_X1  g597(.A1(new_n734), .A2(new_n735), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n784), .A2(new_n317), .A3(new_n360), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n777), .A2(KEYINPUT47), .A3(new_n530), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(KEYINPUT47), .B1(new_n777), .B2(new_n530), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n785), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G140), .ZN(G42));
  NAND3_X1  g604(.A1(new_n705), .A2(new_n594), .A3(new_n530), .ZN(new_n791));
  XOR2_X1   g605(.A(new_n791), .B(KEYINPUT109), .Z(new_n792));
  NAND2_X1  g606(.A1(new_n680), .A2(new_n522), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(KEYINPUT49), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(KEYINPUT110), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n680), .A2(new_n522), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT49), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n747), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n657), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n792), .A2(new_n795), .A3(new_n669), .A4(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n788), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n801), .B(new_n786), .C1(new_n530), .C2(new_n793), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n748), .A2(new_n452), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n803), .A2(new_n702), .A3(new_n705), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n802), .A2(new_n734), .A3(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n657), .A2(new_n594), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n804), .A2(new_n682), .A3(new_n806), .ZN(new_n807));
  XOR2_X1   g621(.A(new_n807), .B(KEYINPUT50), .Z(new_n808));
  NOR2_X1   g622(.A1(new_n681), .A2(new_n720), .ZN(new_n809));
  AND4_X1   g623(.A1(new_n360), .A2(new_n669), .A3(new_n452), .A4(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n810), .A2(new_n623), .A3(new_n746), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n803), .A2(new_n809), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n812), .A2(new_n632), .A3(new_n702), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n805), .A2(new_n808), .A3(new_n811), .A4(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT51), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n451), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n804), .A2(new_n689), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n816), .B(new_n817), .C1(new_n815), .C2(new_n814), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n637), .B1(new_n649), .B2(new_n675), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n632), .A2(new_n642), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n710), .A2(new_n603), .A3(new_n668), .A4(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n819), .A2(new_n716), .A3(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT112), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT52), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n819), .A2(new_n716), .A3(new_n821), .A4(KEYINPUT112), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n827), .B1(new_n825), .B2(new_n822), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT53), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT111), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n450), .A2(new_n642), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n688), .A2(new_n830), .A3(new_n740), .A4(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n740), .A2(new_n317), .A3(new_n632), .A4(new_n831), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(KEYINPUT111), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n702), .A2(new_n632), .A3(new_n735), .A4(new_n740), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n835), .A2(new_n738), .A3(new_n741), .A4(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n712), .A2(new_n683), .A3(new_n686), .A4(new_n690), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n593), .A2(new_n595), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n624), .A2(new_n618), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n604), .A2(new_n609), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n841), .A2(new_n597), .A3(new_n633), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n837), .A2(new_n838), .A3(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n828), .A2(new_n829), .A3(new_n843), .ZN(new_n844));
  AND4_X1   g658(.A1(new_n738), .A2(new_n835), .A3(new_n741), .A4(new_n836), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n838), .A2(new_n842), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n824), .A2(new_n826), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT52), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n847), .B1(new_n849), .B2(new_n827), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n844), .B1(new_n850), .B2(new_n829), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n852));
  OR2_X1    g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g667(.A(KEYINPUT113), .B1(new_n850), .B2(KEYINPUT53), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n842), .B1(new_n838), .B2(KEYINPUT114), .ZN(new_n855));
  OAI21_X1  g669(.A(KEYINPUT53), .B1(new_n838), .B2(KEYINPUT114), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n856), .A2(new_n837), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n828), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n825), .B1(new_n824), .B2(new_n826), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n843), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT113), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n861), .A2(new_n862), .A3(new_n829), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n854), .A2(new_n852), .A3(new_n858), .A4(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n853), .A2(new_n864), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n810), .A2(new_n408), .A3(new_n617), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n726), .A2(new_n730), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n867), .A2(new_n704), .A3(new_n703), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n812), .A2(new_n868), .ZN(new_n869));
  XOR2_X1   g683(.A(new_n869), .B(KEYINPUT48), .Z(new_n870));
  NOR4_X1   g684(.A1(new_n818), .A2(new_n865), .A3(new_n866), .A4(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(G952), .A2(G953), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n800), .B1(new_n871), .B2(new_n872), .ZN(G75));
  AND3_X1   g687(.A1(new_n861), .A2(new_n862), .A3(new_n829), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n862), .B1(new_n861), .B2(new_n829), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n290), .B1(new_n876), .B2(new_n858), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(G210), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT56), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n553), .A2(new_n564), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(new_n562), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n881), .B(KEYINPUT55), .Z(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n878), .A2(KEYINPUT115), .A3(new_n879), .A4(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n854), .A2(new_n858), .A3(new_n863), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(G902), .ZN(new_n886));
  OAI211_X1 g700(.A(KEYINPUT115), .B(new_n879), .C1(new_n886), .C2(new_n271), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(new_n882), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n318), .A2(G952), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n884), .A2(new_n888), .A3(new_n890), .ZN(G51));
  OR2_X1    g705(.A1(new_n518), .A2(new_n521), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n524), .A2(KEYINPUT57), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n852), .B1(new_n876), .B2(new_n858), .ZN(new_n894));
  INV_X1    g708(.A(new_n864), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n524), .A2(KEYINPUT57), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n892), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n877), .A2(new_n772), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n889), .B1(new_n898), .B2(new_n899), .ZN(G54));
  NAND4_X1  g714(.A1(new_n885), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n901));
  INV_X1    g715(.A(new_n393), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(new_n890), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT116), .ZN(new_n905));
  OR3_X1    g719(.A1(new_n901), .A2(new_n905), .A3(new_n902), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n905), .B1(new_n901), .B2(new_n902), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n904), .B1(new_n906), .B2(new_n907), .ZN(G60));
  NAND2_X1  g722(.A1(new_n611), .A2(new_n613), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT117), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n616), .B(KEYINPUT59), .Z(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n910), .B(new_n912), .C1(new_n894), .C2(new_n895), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n890), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT118), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n911), .B1(new_n853), .B2(new_n864), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n915), .B1(new_n916), .B2(new_n910), .ZN(new_n917));
  OR3_X1    g731(.A1(new_n916), .A2(new_n915), .A3(new_n910), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n914), .B1(new_n917), .B2(new_n918), .ZN(G63));
  XNOR2_X1  g733(.A(KEYINPUT119), .B(KEYINPUT60), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n349), .A2(new_n290), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n920), .B(new_n921), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n630), .B(KEYINPUT120), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n885), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n885), .A2(new_n922), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n890), .B(new_n924), .C1(new_n925), .C2(new_n346), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT61), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n926), .B(new_n927), .ZN(G66));
  OAI21_X1  g742(.A(G953), .B1(new_n454), .B2(new_n557), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n929), .B1(new_n846), .B2(G953), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n880), .B1(G898), .B2(new_n318), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n930), .B(new_n931), .ZN(G69));
  NAND2_X1  g746(.A1(new_n738), .A2(new_n741), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n779), .A2(new_n781), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n868), .A2(new_n710), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT124), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n934), .A2(KEYINPUT124), .A3(new_n936), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n933), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n785), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n942), .B1(new_n801), .B2(new_n786), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n819), .A2(new_n716), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(KEYINPUT121), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT121), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n819), .A2(new_n716), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n782), .A2(new_n943), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(KEYINPUT125), .B1(new_n941), .B2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n933), .ZN(new_n951));
  AOI21_X1  g765(.A(KEYINPUT124), .B1(new_n934), .B2(new_n936), .ZN(new_n952));
  AOI211_X1 g766(.A(new_n938), .B(new_n935), .C1(new_n779), .C2(new_n781), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n951), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT125), .ZN(new_n955));
  INV_X1    g769(.A(new_n948), .ZN(new_n956));
  INV_X1    g770(.A(new_n934), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n789), .B(new_n956), .C1(new_n957), .C2(new_n754), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n954), .A2(new_n955), .A3(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n318), .B1(new_n950), .B2(new_n959), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n249), .A2(new_n264), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(new_n388), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n962), .B1(new_n641), .B2(G953), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n318), .B1(G227), .B2(G900), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT123), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT122), .ZN(new_n967));
  OAI211_X1 g781(.A(new_n362), .B(new_n734), .C1(new_n967), .C2(new_n840), .ZN(new_n968));
  AOI211_X1 g782(.A(new_n653), .B(new_n968), .C1(new_n967), .C2(new_n840), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n672), .A2(new_n947), .A3(new_n945), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT62), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n956), .A2(KEYINPUT62), .A3(new_n672), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n969), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n782), .A2(new_n943), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n976), .A2(new_n318), .A3(new_n962), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n964), .A2(KEYINPUT126), .A3(new_n966), .A4(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n966), .A2(KEYINPUT126), .ZN(new_n979));
  OR2_X1    g793(.A1(new_n966), .A2(KEYINPUT126), .ZN(new_n980));
  INV_X1    g794(.A(new_n963), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n955), .B1(new_n954), .B2(new_n958), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n939), .A2(new_n940), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n983), .A2(KEYINPUT125), .A3(new_n951), .A4(new_n949), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n981), .B1(new_n985), .B2(new_n318), .ZN(new_n986));
  INV_X1    g800(.A(new_n977), .ZN(new_n987));
  OAI211_X1 g801(.A(new_n979), .B(new_n980), .C1(new_n986), .C2(new_n987), .ZN(new_n988));
  AND2_X1   g802(.A1(new_n978), .A2(new_n988), .ZN(G72));
  NAND2_X1  g803(.A1(G472), .A2(G902), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT63), .Z(new_n991));
  INV_X1    g805(.A(new_n846), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n991), .B1(new_n985), .B2(new_n992), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n993), .A2(new_n663), .A3(new_n276), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n974), .A2(new_n975), .A3(new_n846), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n995), .A2(new_n991), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(new_n664), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT127), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n996), .A2(KEYINPUT127), .A3(new_n664), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n991), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n295), .A2(new_n274), .ZN(new_n1003));
  OR3_X1    g817(.A1(new_n851), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  AND4_X1   g818(.A1(new_n890), .A2(new_n994), .A3(new_n1001), .A4(new_n1004), .ZN(G57));
endmodule


