

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593;

  XOR2_X1 U324 ( .A(n585), .B(KEYINPUT41), .Z(n565) );
  XOR2_X1 U325 ( .A(n369), .B(n368), .Z(n292) );
  NAND2_X1 U326 ( .A1(n477), .A2(n573), .ZN(n293) );
  AND2_X1 U327 ( .A1(n461), .A2(n534), .ZN(n294) );
  AND2_X1 U328 ( .A1(n565), .A2(n563), .ZN(n424) );
  XNOR2_X1 U329 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U330 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U331 ( .A(n370), .B(n292), .ZN(n371) );
  XNOR2_X1 U332 ( .A(n372), .B(n371), .ZN(n373) );
  AND2_X1 U333 ( .A1(n483), .A2(n294), .ZN(n462) );
  XNOR2_X1 U334 ( .A(n414), .B(n413), .ZN(n573) );
  XNOR2_X1 U335 ( .A(n472), .B(G190GAT), .ZN(n473) );
  XNOR2_X1 U336 ( .A(n474), .B(n473), .ZN(G1351GAT) );
  XOR2_X1 U337 ( .A(G43GAT), .B(G134GAT), .Z(n404) );
  XNOR2_X1 U338 ( .A(G99GAT), .B(G71GAT), .ZN(n295) );
  XNOR2_X1 U339 ( .A(n295), .B(G120GAT), .ZN(n367) );
  XOR2_X1 U340 ( .A(n404), .B(n367), .Z(n297) );
  NAND2_X1 U341 ( .A1(G227GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U342 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U343 ( .A(KEYINPUT87), .B(KEYINPUT65), .Z(n299) );
  XNOR2_X1 U344 ( .A(KEYINPUT84), .B(KEYINPUT20), .ZN(n298) );
  XNOR2_X1 U345 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U346 ( .A(n301), .B(n300), .Z(n303) );
  XOR2_X1 U347 ( .A(G15GAT), .B(G127GAT), .Z(n388) );
  XOR2_X1 U348 ( .A(G113GAT), .B(KEYINPUT0), .Z(n445) );
  XNOR2_X1 U349 ( .A(n388), .B(n445), .ZN(n302) );
  XNOR2_X1 U350 ( .A(n303), .B(n302), .ZN(n311) );
  XOR2_X1 U351 ( .A(KEYINPUT85), .B(KEYINPUT18), .Z(n305) );
  XNOR2_X1 U352 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n304) );
  XNOR2_X1 U353 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U354 ( .A(n306), .B(KEYINPUT19), .Z(n308) );
  XNOR2_X1 U355 ( .A(G190GAT), .B(KEYINPUT86), .ZN(n307) );
  XNOR2_X1 U356 ( .A(n308), .B(n307), .ZN(n310) );
  XOR2_X1 U357 ( .A(G183GAT), .B(G176GAT), .Z(n309) );
  XNOR2_X1 U358 ( .A(n310), .B(n309), .ZN(n356) );
  XOR2_X1 U359 ( .A(n311), .B(n356), .Z(n477) );
  XOR2_X1 U360 ( .A(G22GAT), .B(G197GAT), .Z(n313) );
  XNOR2_X1 U361 ( .A(G36GAT), .B(G141GAT), .ZN(n312) );
  XNOR2_X1 U362 ( .A(n313), .B(n312), .ZN(n317) );
  XOR2_X1 U363 ( .A(KEYINPUT30), .B(G113GAT), .Z(n315) );
  XNOR2_X1 U364 ( .A(G169GAT), .B(G15GAT), .ZN(n314) );
  XNOR2_X1 U365 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U366 ( .A(n317), .B(n316), .Z(n322) );
  XOR2_X1 U367 ( .A(KEYINPUT71), .B(KEYINPUT70), .Z(n319) );
  NAND2_X1 U368 ( .A1(G229GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U369 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U370 ( .A(KEYINPUT69), .B(n320), .ZN(n321) );
  XNOR2_X1 U371 ( .A(n322), .B(n321), .ZN(n331) );
  XOR2_X1 U372 ( .A(KEYINPUT74), .B(KEYINPUT73), .Z(n324) );
  XNOR2_X1 U373 ( .A(KEYINPUT29), .B(KEYINPUT72), .ZN(n323) );
  XNOR2_X1 U374 ( .A(n324), .B(n323), .ZN(n329) );
  XOR2_X1 U375 ( .A(G8GAT), .B(G1GAT), .Z(n376) );
  XNOR2_X1 U376 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n325) );
  XNOR2_X1 U377 ( .A(n325), .B(KEYINPUT7), .ZN(n410) );
  XOR2_X1 U378 ( .A(n376), .B(n410), .Z(n327) );
  XNOR2_X1 U379 ( .A(G50GAT), .B(G43GAT), .ZN(n326) );
  XNOR2_X1 U380 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U381 ( .A(n329), .B(n328), .Z(n330) );
  XOR2_X1 U382 ( .A(n331), .B(n330), .Z(n580) );
  INV_X1 U383 ( .A(n580), .ZN(n563) );
  NAND2_X1 U384 ( .A1(n477), .A2(n563), .ZN(n463) );
  XOR2_X1 U385 ( .A(KEYINPUT24), .B(KEYINPUT90), .Z(n333) );
  XNOR2_X1 U386 ( .A(G204GAT), .B(KEYINPUT22), .ZN(n332) );
  XNOR2_X1 U387 ( .A(n333), .B(n332), .ZN(n337) );
  XOR2_X1 U388 ( .A(KEYINPUT89), .B(KEYINPUT23), .Z(n335) );
  XOR2_X1 U389 ( .A(G50GAT), .B(G162GAT), .Z(n401) );
  XOR2_X1 U390 ( .A(G22GAT), .B(G155GAT), .Z(n378) );
  XNOR2_X1 U391 ( .A(n401), .B(n378), .ZN(n334) );
  XNOR2_X1 U392 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U393 ( .A(n337), .B(n336), .Z(n339) );
  NAND2_X1 U394 ( .A1(G228GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U395 ( .A(n339), .B(n338), .ZN(n341) );
  XNOR2_X1 U396 ( .A(G106GAT), .B(G78GAT), .ZN(n340) );
  XNOR2_X1 U397 ( .A(n340), .B(G148GAT), .ZN(n359) );
  XOR2_X1 U398 ( .A(n341), .B(n359), .Z(n348) );
  XOR2_X1 U399 ( .A(KEYINPUT91), .B(G218GAT), .Z(n343) );
  XNOR2_X1 U400 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n342) );
  XNOR2_X1 U401 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U402 ( .A(G197GAT), .B(n344), .Z(n350) );
  XOR2_X1 U403 ( .A(KEYINPUT3), .B(KEYINPUT92), .Z(n346) );
  XNOR2_X1 U404 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n345) );
  XNOR2_X1 U405 ( .A(n346), .B(n345), .ZN(n446) );
  XNOR2_X1 U406 ( .A(n350), .B(n446), .ZN(n347) );
  XNOR2_X1 U407 ( .A(n348), .B(n347), .ZN(n483) );
  XOR2_X1 U408 ( .A(G36GAT), .B(KEYINPUT80), .Z(n402) );
  XNOR2_X1 U409 ( .A(G204GAT), .B(G92GAT), .ZN(n349) );
  XNOR2_X1 U410 ( .A(n349), .B(G64GAT), .ZN(n366) );
  XOR2_X1 U411 ( .A(KEYINPUT98), .B(n366), .Z(n352) );
  XNOR2_X1 U412 ( .A(G8GAT), .B(n350), .ZN(n351) );
  XNOR2_X1 U413 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U414 ( .A(n402), .B(n353), .Z(n355) );
  NAND2_X1 U415 ( .A1(G226GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U416 ( .A(n355), .B(n354), .ZN(n357) );
  XOR2_X1 U417 ( .A(n357), .B(n356), .Z(n536) );
  XOR2_X1 U418 ( .A(KEYINPUT122), .B(n536), .Z(n434) );
  XNOR2_X1 U419 ( .A(G176GAT), .B(KEYINPUT13), .ZN(n358) );
  XNOR2_X1 U420 ( .A(G85GAT), .B(G57GAT), .ZN(n451) );
  XNOR2_X1 U421 ( .A(n358), .B(n451), .ZN(n374) );
  NAND2_X1 U422 ( .A1(n359), .A2(KEYINPUT75), .ZN(n363) );
  INV_X1 U423 ( .A(n359), .ZN(n361) );
  INV_X1 U424 ( .A(KEYINPUT75), .ZN(n360) );
  NAND2_X1 U425 ( .A1(n361), .A2(n360), .ZN(n362) );
  NAND2_X1 U426 ( .A1(n363), .A2(n362), .ZN(n365) );
  AND2_X1 U427 ( .A1(G230GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U428 ( .A(n365), .B(n364), .ZN(n372) );
  XNOR2_X1 U429 ( .A(n367), .B(n366), .ZN(n370) );
  XOR2_X1 U430 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n369) );
  XNOR2_X1 U431 ( .A(KEYINPUT33), .B(KEYINPUT76), .ZN(n368) );
  XNOR2_X1 U432 ( .A(n374), .B(n373), .ZN(n585) );
  XOR2_X1 U433 ( .A(KEYINPUT115), .B(KEYINPUT45), .Z(n375) );
  XNOR2_X1 U434 ( .A(KEYINPUT67), .B(n375), .ZN(n421) );
  XNOR2_X1 U435 ( .A(n376), .B(G211GAT), .ZN(n377) );
  XNOR2_X1 U436 ( .A(n377), .B(G78GAT), .ZN(n392) );
  XOR2_X1 U437 ( .A(n378), .B(KEYINPUT82), .Z(n380) );
  NAND2_X1 U438 ( .A1(G231GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U439 ( .A(n380), .B(n379), .ZN(n384) );
  XOR2_X1 U440 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n382) );
  XNOR2_X1 U441 ( .A(KEYINPUT13), .B(G64GAT), .ZN(n381) );
  XNOR2_X1 U442 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U443 ( .A(n384), .B(n383), .Z(n390) );
  XOR2_X1 U444 ( .A(G57GAT), .B(KEYINPUT14), .Z(n386) );
  XNOR2_X1 U445 ( .A(G183GAT), .B(G71GAT), .ZN(n385) );
  XNOR2_X1 U446 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U447 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U448 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U449 ( .A(n392), .B(n391), .Z(n490) );
  INV_X1 U450 ( .A(n490), .ZN(n588) );
  XNOR2_X1 U451 ( .A(KEYINPUT36), .B(KEYINPUT102), .ZN(n415) );
  XOR2_X1 U452 ( .A(KEYINPUT10), .B(KEYINPUT79), .Z(n394) );
  XNOR2_X1 U453 ( .A(KEYINPUT66), .B(KEYINPUT78), .ZN(n393) );
  XNOR2_X1 U454 ( .A(n394), .B(n393), .ZN(n414) );
  XOR2_X1 U455 ( .A(KEYINPUT81), .B(KEYINPUT11), .Z(n396) );
  XNOR2_X1 U456 ( .A(G218GAT), .B(G106GAT), .ZN(n395) );
  XNOR2_X1 U457 ( .A(n396), .B(n395), .ZN(n400) );
  XOR2_X1 U458 ( .A(KEYINPUT9), .B(G85GAT), .Z(n398) );
  XNOR2_X1 U459 ( .A(G99GAT), .B(G92GAT), .ZN(n397) );
  XNOR2_X1 U460 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U461 ( .A(n400), .B(n399), .Z(n408) );
  XOR2_X1 U462 ( .A(n402), .B(n401), .Z(n406) );
  NAND2_X1 U463 ( .A1(G232GAT), .A2(G233GAT), .ZN(n403) );
  XNOR2_X1 U464 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U465 ( .A(n409), .B(KEYINPUT77), .Z(n412) );
  XNOR2_X1 U466 ( .A(n410), .B(G190GAT), .ZN(n411) );
  XNOR2_X1 U467 ( .A(n412), .B(n411), .ZN(n413) );
  NAND2_X1 U468 ( .A1(n415), .A2(n573), .ZN(n419) );
  INV_X1 U469 ( .A(n415), .ZN(n417) );
  INV_X1 U470 ( .A(n573), .ZN(n416) );
  NAND2_X1 U471 ( .A1(n417), .A2(n416), .ZN(n418) );
  NAND2_X1 U472 ( .A1(n419), .A2(n418), .ZN(n591) );
  NAND2_X1 U473 ( .A1(n588), .A2(n591), .ZN(n420) );
  XOR2_X1 U474 ( .A(n421), .B(n420), .Z(n422) );
  NOR2_X1 U475 ( .A1(n585), .A2(n422), .ZN(n423) );
  NAND2_X1 U476 ( .A1(n423), .A2(n580), .ZN(n431) );
  XNOR2_X1 U477 ( .A(KEYINPUT47), .B(KEYINPUT114), .ZN(n429) );
  XNOR2_X1 U478 ( .A(n424), .B(KEYINPUT46), .ZN(n425) );
  NOR2_X1 U479 ( .A1(n588), .A2(n425), .ZN(n426) );
  XNOR2_X1 U480 ( .A(n426), .B(KEYINPUT113), .ZN(n427) );
  NOR2_X1 U481 ( .A1(n427), .A2(n573), .ZN(n428) );
  XNOR2_X1 U482 ( .A(n429), .B(n428), .ZN(n430) );
  NAND2_X1 U483 ( .A1(n431), .A2(n430), .ZN(n433) );
  XNOR2_X1 U484 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n432) );
  XNOR2_X1 U485 ( .A(n433), .B(n432), .ZN(n546) );
  NAND2_X1 U486 ( .A1(n434), .A2(n546), .ZN(n435) );
  XNOR2_X1 U487 ( .A(n435), .B(KEYINPUT123), .ZN(n436) );
  XNOR2_X1 U488 ( .A(n436), .B(KEYINPUT54), .ZN(n461) );
  XOR2_X1 U489 ( .A(KEYINPUT1), .B(KEYINPUT96), .Z(n438) );
  XNOR2_X1 U490 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n437) );
  XNOR2_X1 U491 ( .A(n438), .B(n437), .ZN(n460) );
  XOR2_X1 U492 ( .A(KEYINPUT95), .B(G120GAT), .Z(n440) );
  XNOR2_X1 U493 ( .A(G1GAT), .B(G127GAT), .ZN(n439) );
  XNOR2_X1 U494 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U495 ( .A(KEYINPUT93), .B(KEYINPUT97), .Z(n442) );
  XNOR2_X1 U496 ( .A(KEYINPUT94), .B(KEYINPUT6), .ZN(n441) );
  XNOR2_X1 U497 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U498 ( .A(n444), .B(n443), .Z(n458) );
  XOR2_X1 U499 ( .A(n446), .B(n445), .Z(n448) );
  NAND2_X1 U500 ( .A1(G225GAT), .A2(G233GAT), .ZN(n447) );
  XNOR2_X1 U501 ( .A(n448), .B(n447), .ZN(n456) );
  XOR2_X1 U502 ( .A(G155GAT), .B(G162GAT), .Z(n450) );
  XNOR2_X1 U503 ( .A(G134GAT), .B(G148GAT), .ZN(n449) );
  XNOR2_X1 U504 ( .A(n450), .B(n449), .ZN(n452) );
  XNOR2_X1 U505 ( .A(n452), .B(n451), .ZN(n454) );
  XNOR2_X1 U506 ( .A(G29GAT), .B(KEYINPUT79), .ZN(n453) );
  XNOR2_X1 U507 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U508 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U509 ( .A(n458), .B(n457), .ZN(n459) );
  XOR2_X1 U510 ( .A(n460), .B(n459), .Z(n534) );
  INV_X1 U511 ( .A(n534), .ZN(n481) );
  XNOR2_X1 U512 ( .A(KEYINPUT55), .B(n462), .ZN(n575) );
  OR2_X1 U513 ( .A1(n463), .A2(n575), .ZN(n466) );
  XOR2_X1 U514 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n464) );
  XNOR2_X1 U515 ( .A(n464), .B(G169GAT), .ZN(n465) );
  XNOR2_X1 U516 ( .A(n466), .B(n465), .ZN(G1348GAT) );
  NAND2_X1 U517 ( .A1(n477), .A2(n565), .ZN(n467) );
  OR2_X1 U518 ( .A1(n467), .A2(n575), .ZN(n471) );
  XOR2_X1 U519 ( .A(G176GAT), .B(KEYINPUT126), .Z(n469) );
  XNOR2_X1 U520 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n468) );
  XNOR2_X1 U521 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U522 ( .A(n471), .B(n470), .ZN(G1349GAT) );
  OR2_X1 U523 ( .A1(n293), .A2(n575), .ZN(n474) );
  XOR2_X1 U524 ( .A(KEYINPUT58), .B(KEYINPUT127), .Z(n472) );
  NOR2_X1 U525 ( .A1(n580), .A2(n585), .ZN(n508) );
  INV_X1 U526 ( .A(n477), .ZN(n576) );
  OR2_X1 U527 ( .A1(n536), .A2(n576), .ZN(n475) );
  NAND2_X1 U528 ( .A1(n483), .A2(n475), .ZN(n476) );
  XNOR2_X1 U529 ( .A(n476), .B(KEYINPUT25), .ZN(n480) );
  NOR2_X1 U530 ( .A1(n483), .A2(n477), .ZN(n478) );
  XOR2_X1 U531 ( .A(KEYINPUT26), .B(n478), .Z(n560) );
  XNOR2_X1 U532 ( .A(n536), .B(KEYINPUT27), .ZN(n485) );
  NOR2_X1 U533 ( .A1(n560), .A2(n485), .ZN(n479) );
  NOR2_X1 U534 ( .A1(n480), .A2(n479), .ZN(n482) );
  NOR2_X1 U535 ( .A1(n482), .A2(n481), .ZN(n489) );
  XOR2_X1 U536 ( .A(KEYINPUT88), .B(n576), .Z(n487) );
  XNOR2_X1 U537 ( .A(n483), .B(KEYINPUT68), .ZN(n484) );
  XNOR2_X1 U538 ( .A(n484), .B(KEYINPUT28), .ZN(n548) );
  NOR2_X1 U539 ( .A1(n534), .A2(n485), .ZN(n545) );
  NAND2_X1 U540 ( .A1(n548), .A2(n545), .ZN(n486) );
  NOR2_X1 U541 ( .A1(n487), .A2(n486), .ZN(n488) );
  NOR2_X1 U542 ( .A1(n489), .A2(n488), .ZN(n504) );
  NOR2_X1 U543 ( .A1(n490), .A2(n573), .ZN(n492) );
  XNOR2_X1 U544 ( .A(KEYINPUT16), .B(KEYINPUT83), .ZN(n491) );
  XNOR2_X1 U545 ( .A(n492), .B(n491), .ZN(n493) );
  NOR2_X1 U546 ( .A1(n504), .A2(n493), .ZN(n522) );
  NAND2_X1 U547 ( .A1(n508), .A2(n522), .ZN(n502) );
  NOR2_X1 U548 ( .A1(n534), .A2(n502), .ZN(n495) );
  XNOR2_X1 U549 ( .A(KEYINPUT34), .B(KEYINPUT99), .ZN(n494) );
  XNOR2_X1 U550 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U551 ( .A(G1GAT), .B(n496), .ZN(G1324GAT) );
  NOR2_X1 U552 ( .A1(n536), .A2(n502), .ZN(n497) );
  XOR2_X1 U553 ( .A(KEYINPUT100), .B(n497), .Z(n498) );
  XNOR2_X1 U554 ( .A(G8GAT), .B(n498), .ZN(G1325GAT) );
  NOR2_X1 U555 ( .A1(n576), .A2(n502), .ZN(n500) );
  XNOR2_X1 U556 ( .A(KEYINPUT101), .B(KEYINPUT35), .ZN(n499) );
  XNOR2_X1 U557 ( .A(n500), .B(n499), .ZN(n501) );
  XOR2_X1 U558 ( .A(G15GAT), .B(n501), .Z(G1326GAT) );
  NOR2_X1 U559 ( .A1(n548), .A2(n502), .ZN(n503) );
  XOR2_X1 U560 ( .A(G22GAT), .B(n503), .Z(G1327GAT) );
  XOR2_X1 U561 ( .A(KEYINPUT103), .B(KEYINPUT37), .Z(n507) );
  NOR2_X1 U562 ( .A1(n504), .A2(n588), .ZN(n505) );
  NAND2_X1 U563 ( .A1(n505), .A2(n591), .ZN(n506) );
  XNOR2_X1 U564 ( .A(n507), .B(n506), .ZN(n533) );
  NAND2_X1 U565 ( .A1(n533), .A2(n508), .ZN(n510) );
  XNOR2_X1 U566 ( .A(KEYINPUT38), .B(KEYINPUT104), .ZN(n509) );
  XNOR2_X1 U567 ( .A(n510), .B(n509), .ZN(n519) );
  NOR2_X1 U568 ( .A1(n534), .A2(n519), .ZN(n512) );
  XNOR2_X1 U569 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n511) );
  XNOR2_X1 U570 ( .A(n512), .B(n511), .ZN(G1328GAT) );
  NOR2_X1 U571 ( .A1(n536), .A2(n519), .ZN(n514) );
  XNOR2_X1 U572 ( .A(G36GAT), .B(KEYINPUT105), .ZN(n513) );
  XNOR2_X1 U573 ( .A(n514), .B(n513), .ZN(G1329GAT) );
  XOR2_X1 U574 ( .A(KEYINPUT40), .B(KEYINPUT106), .Z(n516) );
  XNOR2_X1 U575 ( .A(G43GAT), .B(KEYINPUT107), .ZN(n515) );
  XNOR2_X1 U576 ( .A(n516), .B(n515), .ZN(n518) );
  NOR2_X1 U577 ( .A1(n576), .A2(n519), .ZN(n517) );
  XOR2_X1 U578 ( .A(n518), .B(n517), .Z(G1330GAT) );
  NOR2_X1 U579 ( .A1(n548), .A2(n519), .ZN(n520) );
  XOR2_X1 U580 ( .A(G50GAT), .B(n520), .Z(G1331GAT) );
  INV_X1 U581 ( .A(n565), .ZN(n521) );
  NOR2_X1 U582 ( .A1(n563), .A2(n521), .ZN(n532) );
  NAND2_X1 U583 ( .A1(n532), .A2(n522), .ZN(n528) );
  NOR2_X1 U584 ( .A1(n534), .A2(n528), .ZN(n524) );
  XNOR2_X1 U585 ( .A(KEYINPUT108), .B(KEYINPUT42), .ZN(n523) );
  XNOR2_X1 U586 ( .A(n524), .B(n523), .ZN(n525) );
  XOR2_X1 U587 ( .A(G57GAT), .B(n525), .Z(G1332GAT) );
  NOR2_X1 U588 ( .A1(n536), .A2(n528), .ZN(n526) );
  XOR2_X1 U589 ( .A(G64GAT), .B(n526), .Z(G1333GAT) );
  NOR2_X1 U590 ( .A1(n576), .A2(n528), .ZN(n527) );
  XOR2_X1 U591 ( .A(G71GAT), .B(n527), .Z(G1334GAT) );
  NOR2_X1 U592 ( .A1(n548), .A2(n528), .ZN(n530) );
  XNOR2_X1 U593 ( .A(KEYINPUT109), .B(KEYINPUT43), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n530), .B(n529), .ZN(n531) );
  XOR2_X1 U595 ( .A(G78GAT), .B(n531), .Z(G1335GAT) );
  NAND2_X1 U596 ( .A1(n533), .A2(n532), .ZN(n541) );
  NOR2_X1 U597 ( .A1(n534), .A2(n541), .ZN(n535) );
  XOR2_X1 U598 ( .A(G85GAT), .B(n535), .Z(G1336GAT) );
  NOR2_X1 U599 ( .A1(n536), .A2(n541), .ZN(n537) );
  XOR2_X1 U600 ( .A(KEYINPUT110), .B(n537), .Z(n538) );
  XNOR2_X1 U601 ( .A(G92GAT), .B(n538), .ZN(G1337GAT) );
  NOR2_X1 U602 ( .A1(n576), .A2(n541), .ZN(n540) );
  XNOR2_X1 U603 ( .A(G99GAT), .B(KEYINPUT111), .ZN(n539) );
  XNOR2_X1 U604 ( .A(n540), .B(n539), .ZN(G1338GAT) );
  NOR2_X1 U605 ( .A1(n548), .A2(n541), .ZN(n543) );
  XNOR2_X1 U606 ( .A(KEYINPUT44), .B(KEYINPUT112), .ZN(n542) );
  XNOR2_X1 U607 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U608 ( .A(G106GAT), .B(n544), .Z(G1339GAT) );
  NAND2_X1 U609 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U610 ( .A(KEYINPUT116), .B(n547), .Z(n561) );
  NAND2_X1 U611 ( .A1(n548), .A2(n561), .ZN(n549) );
  NOR2_X1 U612 ( .A1(n576), .A2(n549), .ZN(n557) );
  NAND2_X1 U613 ( .A1(n557), .A2(n563), .ZN(n550) );
  XNOR2_X1 U614 ( .A(G113GAT), .B(n550), .ZN(G1340GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT117), .B(KEYINPUT49), .Z(n552) );
  NAND2_X1 U616 ( .A1(n557), .A2(n565), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n552), .B(n551), .ZN(n553) );
  XOR2_X1 U618 ( .A(G120GAT), .B(n553), .Z(G1341GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n555) );
  NAND2_X1 U620 ( .A1(n557), .A2(n588), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U622 ( .A(G127GAT), .B(n556), .Z(G1342GAT) );
  XOR2_X1 U623 ( .A(G134GAT), .B(KEYINPUT51), .Z(n559) );
  NAND2_X1 U624 ( .A1(n557), .A2(n573), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(G1343GAT) );
  INV_X1 U626 ( .A(n560), .ZN(n579) );
  NAND2_X1 U627 ( .A1(n561), .A2(n579), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(KEYINPUT119), .ZN(n572) );
  NAND2_X1 U629 ( .A1(n572), .A2(n563), .ZN(n564) );
  XNOR2_X1 U630 ( .A(G141GAT), .B(n564), .ZN(G1344GAT) );
  XNOR2_X1 U631 ( .A(G148GAT), .B(KEYINPUT120), .ZN(n569) );
  XOR2_X1 U632 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n567) );
  NAND2_X1 U633 ( .A1(n572), .A2(n565), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(G1345GAT) );
  XOR2_X1 U636 ( .A(G155GAT), .B(KEYINPUT121), .Z(n571) );
  NAND2_X1 U637 ( .A1(n572), .A2(n588), .ZN(n570) );
  XNOR2_X1 U638 ( .A(n571), .B(n570), .ZN(G1346GAT) );
  NAND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n574), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U642 ( .A1(n588), .A2(n577), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n578), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U644 ( .A1(n294), .A2(n579), .ZN(n584) );
  NOR2_X1 U645 ( .A1(n580), .A2(n584), .ZN(n582) );
  XNOR2_X1 U646 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(G197GAT), .B(n583), .ZN(G1352GAT) );
  XOR2_X1 U649 ( .A(G204GAT), .B(KEYINPUT61), .Z(n587) );
  INV_X1 U650 ( .A(n584), .ZN(n590) );
  NAND2_X1 U651 ( .A1(n590), .A2(n585), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(G1353GAT) );
  NAND2_X1 U653 ( .A1(n588), .A2(n590), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n589), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U656 ( .A(n592), .B(KEYINPUT62), .ZN(n593) );
  XNOR2_X1 U657 ( .A(G218GAT), .B(n593), .ZN(G1355GAT) );
endmodule

