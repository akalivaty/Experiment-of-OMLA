

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593;

  XNOR2_X1 U326 ( .A(n340), .B(n295), .ZN(n524) );
  AND2_X1 U327 ( .A1(G226GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U328 ( .A(G218GAT), .B(n325), .ZN(n295) );
  INV_X1 U329 ( .A(KEYINPUT27), .ZN(n341) );
  XNOR2_X1 U330 ( .A(n524), .B(n341), .ZN(n384) );
  INV_X1 U331 ( .A(G169GAT), .ZN(n299) );
  XNOR2_X1 U332 ( .A(n300), .B(n299), .ZN(n302) );
  XNOR2_X1 U333 ( .A(n467), .B(KEYINPUT48), .ZN(n533) );
  XNOR2_X1 U334 ( .A(n302), .B(n301), .ZN(n334) );
  INV_X1 U335 ( .A(KEYINPUT55), .ZN(n472) );
  XNOR2_X1 U336 ( .A(n393), .B(n294), .ZN(n337) );
  XNOR2_X1 U337 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U338 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U339 ( .A(n475), .B(n474), .ZN(n476) );
  INV_X1 U340 ( .A(n524), .ZN(n499) );
  XNOR2_X1 U341 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U342 ( .A(n452), .B(KEYINPUT40), .ZN(n453) );
  XNOR2_X1 U343 ( .A(n480), .B(n479), .ZN(G1349GAT) );
  XNOR2_X1 U344 ( .A(n454), .B(n453), .ZN(G1330GAT) );
  XOR2_X1 U345 ( .A(G176GAT), .B(KEYINPUT20), .Z(n297) );
  NAND2_X1 U346 ( .A1(G227GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U347 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U348 ( .A(n298), .B(KEYINPUT64), .Z(n307) );
  XNOR2_X1 U349 ( .A(KEYINPUT19), .B(G183GAT), .ZN(n300) );
  XOR2_X1 U350 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n301) );
  XOR2_X1 U351 ( .A(KEYINPUT86), .B(G99GAT), .Z(n304) );
  XNOR2_X1 U352 ( .A(G43GAT), .B(G190GAT), .ZN(n303) );
  XNOR2_X1 U353 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U354 ( .A(n334), .B(n305), .ZN(n306) );
  XNOR2_X1 U355 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U356 ( .A(G120GAT), .B(G71GAT), .Z(n438) );
  XOR2_X1 U357 ( .A(n308), .B(n438), .Z(n311) );
  XNOR2_X1 U358 ( .A(G113GAT), .B(G134GAT), .ZN(n309) );
  XNOR2_X1 U359 ( .A(n309), .B(KEYINPUT0), .ZN(n345) );
  XOR2_X1 U360 ( .A(G15GAT), .B(G127GAT), .Z(n405) );
  XNOR2_X1 U361 ( .A(n345), .B(n405), .ZN(n310) );
  XOR2_X1 U362 ( .A(n311), .B(n310), .Z(n526) );
  INV_X1 U363 ( .A(n526), .ZN(n536) );
  INV_X1 U364 ( .A(KEYINPUT38), .ZN(n451) );
  XNOR2_X1 U365 ( .A(G43GAT), .B(KEYINPUT73), .ZN(n312) );
  XNOR2_X1 U366 ( .A(n312), .B(G29GAT), .ZN(n313) );
  XOR2_X1 U367 ( .A(n313), .B(KEYINPUT72), .Z(n315) );
  XNOR2_X1 U368 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n314) );
  XNOR2_X1 U369 ( .A(n315), .B(n314), .ZN(n430) );
  XNOR2_X1 U370 ( .A(KEYINPUT66), .B(KEYINPUT10), .ZN(n317) );
  XNOR2_X1 U371 ( .A(G134GAT), .B(KEYINPUT9), .ZN(n316) );
  XNOR2_X1 U372 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U373 ( .A(G50GAT), .B(G162GAT), .Z(n366) );
  XNOR2_X1 U374 ( .A(n318), .B(n366), .ZN(n320) );
  NAND2_X1 U375 ( .A1(G232GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U376 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U377 ( .A(KEYINPUT11), .B(KEYINPUT65), .Z(n322) );
  XNOR2_X1 U378 ( .A(KEYINPUT79), .B(KEYINPUT80), .ZN(n321) );
  XOR2_X1 U379 ( .A(n322), .B(n321), .Z(n323) );
  XNOR2_X1 U380 ( .A(n324), .B(n323), .ZN(n329) );
  XOR2_X1 U381 ( .A(G36GAT), .B(G190GAT), .Z(n325) );
  XOR2_X1 U382 ( .A(G92GAT), .B(G85GAT), .Z(n327) );
  XNOR2_X1 U383 ( .A(G99GAT), .B(G106GAT), .ZN(n326) );
  XNOR2_X1 U384 ( .A(n327), .B(n326), .ZN(n435) );
  XOR2_X1 U385 ( .A(n295), .B(n435), .Z(n328) );
  XNOR2_X1 U386 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U387 ( .A(n430), .B(n330), .Z(n461) );
  INV_X1 U388 ( .A(n461), .ZN(n560) );
  XOR2_X1 U389 ( .A(n560), .B(KEYINPUT81), .Z(n567) );
  INV_X1 U390 ( .A(KEYINPUT36), .ZN(n331) );
  XNOR2_X1 U391 ( .A(n567), .B(n331), .ZN(n591) );
  XOR2_X1 U392 ( .A(G204GAT), .B(G211GAT), .Z(n333) );
  XNOR2_X1 U393 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n332) );
  XNOR2_X1 U394 ( .A(n333), .B(n332), .ZN(n375) );
  XOR2_X1 U395 ( .A(G176GAT), .B(G64GAT), .Z(n445) );
  XOR2_X1 U396 ( .A(n445), .B(KEYINPUT92), .Z(n336) );
  XNOR2_X1 U397 ( .A(n334), .B(G92GAT), .ZN(n335) );
  XNOR2_X1 U398 ( .A(n336), .B(n335), .ZN(n338) );
  XOR2_X1 U399 ( .A(G8GAT), .B(KEYINPUT82), .Z(n393) );
  XNOR2_X1 U400 ( .A(n375), .B(n339), .ZN(n340) );
  XOR2_X1 U401 ( .A(KEYINPUT2), .B(KEYINPUT88), .Z(n343) );
  XNOR2_X1 U402 ( .A(KEYINPUT3), .B(KEYINPUT87), .ZN(n342) );
  XNOR2_X1 U403 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U404 ( .A(G141GAT), .B(n344), .Z(n371) );
  XOR2_X1 U405 ( .A(G85GAT), .B(G155GAT), .Z(n347) );
  XNOR2_X1 U406 ( .A(n345), .B(G162GAT), .ZN(n346) );
  XNOR2_X1 U407 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U408 ( .A(G29GAT), .B(n348), .ZN(n361) );
  XOR2_X1 U409 ( .A(G148GAT), .B(G120GAT), .Z(n350) );
  XNOR2_X1 U410 ( .A(G1GAT), .B(G127GAT), .ZN(n349) );
  XNOR2_X1 U411 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U412 ( .A(KEYINPUT5), .B(KEYINPUT1), .Z(n352) );
  XNOR2_X1 U413 ( .A(KEYINPUT91), .B(KEYINPUT6), .ZN(n351) );
  XNOR2_X1 U414 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U415 ( .A(n354), .B(n353), .Z(n359) );
  XOR2_X1 U416 ( .A(KEYINPUT4), .B(G57GAT), .Z(n356) );
  NAND2_X1 U417 ( .A1(G225GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U418 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U419 ( .A(KEYINPUT90), .B(n357), .ZN(n358) );
  XNOR2_X1 U420 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U421 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U422 ( .A(n371), .B(n362), .Z(n520) );
  INV_X1 U423 ( .A(n520), .ZN(n575) );
  NOR2_X1 U424 ( .A1(n384), .A2(n575), .ZN(n363) );
  XOR2_X1 U425 ( .A(n363), .B(KEYINPUT93), .Z(n534) );
  XOR2_X1 U426 ( .A(G22GAT), .B(G155GAT), .Z(n402) );
  XOR2_X1 U427 ( .A(G148GAT), .B(G78GAT), .Z(n437) );
  XOR2_X1 U428 ( .A(n402), .B(n437), .Z(n365) );
  NAND2_X1 U429 ( .A1(G228GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U430 ( .A(n365), .B(n364), .ZN(n367) );
  XOR2_X1 U431 ( .A(n367), .B(n366), .Z(n373) );
  XOR2_X1 U432 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n369) );
  XNOR2_X1 U433 ( .A(G218GAT), .B(G106GAT), .ZN(n368) );
  XNOR2_X1 U434 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U435 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U436 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U437 ( .A(n374), .B(KEYINPUT23), .Z(n377) );
  XNOR2_X1 U438 ( .A(n375), .B(KEYINPUT89), .ZN(n376) );
  XNOR2_X1 U439 ( .A(n377), .B(n376), .ZN(n470) );
  XNOR2_X1 U440 ( .A(n470), .B(KEYINPUT67), .ZN(n378) );
  XOR2_X1 U441 ( .A(n378), .B(KEYINPUT28), .Z(n529) );
  NOR2_X1 U442 ( .A1(n529), .A2(n526), .ZN(n379) );
  AND2_X1 U443 ( .A1(n534), .A2(n379), .ZN(n389) );
  AND2_X1 U444 ( .A1(n526), .A2(n524), .ZN(n380) );
  OR2_X1 U445 ( .A1(n470), .A2(n380), .ZN(n381) );
  XNOR2_X1 U446 ( .A(n381), .B(KEYINPUT25), .ZN(n382) );
  XNOR2_X1 U447 ( .A(n382), .B(KEYINPUT94), .ZN(n386) );
  NAND2_X1 U448 ( .A1(n470), .A2(n536), .ZN(n383) );
  XNOR2_X1 U449 ( .A(n383), .B(KEYINPUT26), .ZN(n578) );
  NOR2_X1 U450 ( .A1(n578), .A2(n384), .ZN(n385) );
  NOR2_X1 U451 ( .A1(n386), .A2(n385), .ZN(n387) );
  NOR2_X1 U452 ( .A1(n387), .A2(n520), .ZN(n388) );
  NOR2_X1 U453 ( .A1(n389), .A2(n388), .ZN(n483) );
  XOR2_X1 U454 ( .A(KEYINPUT85), .B(KEYINPUT83), .Z(n391) );
  NAND2_X1 U455 ( .A1(G231GAT), .A2(G233GAT), .ZN(n390) );
  XNOR2_X1 U456 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U457 ( .A(KEYINPUT84), .B(n392), .Z(n409) );
  XOR2_X1 U458 ( .A(G57GAT), .B(KEYINPUT13), .Z(n444) );
  XOR2_X1 U459 ( .A(n444), .B(n393), .Z(n395) );
  XNOR2_X1 U460 ( .A(G211GAT), .B(G78GAT), .ZN(n394) );
  XNOR2_X1 U461 ( .A(n395), .B(n394), .ZN(n399) );
  XOR2_X1 U462 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n397) );
  XNOR2_X1 U463 ( .A(G64GAT), .B(KEYINPUT15), .ZN(n396) );
  XNOR2_X1 U464 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U465 ( .A(n399), .B(n398), .Z(n401) );
  XNOR2_X1 U466 ( .A(G183GAT), .B(G71GAT), .ZN(n400) );
  XNOR2_X1 U467 ( .A(n401), .B(n400), .ZN(n403) );
  XOR2_X1 U468 ( .A(n403), .B(n402), .Z(n407) );
  XNOR2_X1 U469 ( .A(G1GAT), .B(KEYINPUT74), .ZN(n404) );
  XNOR2_X1 U470 ( .A(n404), .B(KEYINPUT75), .ZN(n425) );
  XNOR2_X1 U471 ( .A(n425), .B(n405), .ZN(n406) );
  XNOR2_X1 U472 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U473 ( .A(n409), .B(n408), .Z(n481) );
  INV_X1 U474 ( .A(n481), .ZN(n586) );
  NOR2_X1 U475 ( .A1(n483), .A2(n586), .ZN(n411) );
  INV_X1 U476 ( .A(KEYINPUT98), .ZN(n410) );
  XNOR2_X1 U477 ( .A(n411), .B(n410), .ZN(n412) );
  NOR2_X1 U478 ( .A1(n591), .A2(n412), .ZN(n413) );
  XNOR2_X1 U479 ( .A(n413), .B(KEYINPUT37), .ZN(n519) );
  XOR2_X1 U480 ( .A(G15GAT), .B(G113GAT), .Z(n415) );
  XNOR2_X1 U481 ( .A(G169GAT), .B(G141GAT), .ZN(n414) );
  XNOR2_X1 U482 ( .A(n415), .B(n414), .ZN(n419) );
  XOR2_X1 U483 ( .A(KEYINPUT69), .B(KEYINPUT70), .Z(n417) );
  XNOR2_X1 U484 ( .A(G8GAT), .B(KEYINPUT71), .ZN(n416) );
  XNOR2_X1 U485 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U486 ( .A(n419), .B(n418), .Z(n424) );
  XOR2_X1 U487 ( .A(KEYINPUT30), .B(KEYINPUT68), .Z(n421) );
  NAND2_X1 U488 ( .A1(G229GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U489 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U490 ( .A(KEYINPUT29), .B(n422), .ZN(n423) );
  XNOR2_X1 U491 ( .A(n424), .B(n423), .ZN(n429) );
  XOR2_X1 U492 ( .A(G36GAT), .B(G50GAT), .Z(n427) );
  XNOR2_X1 U493 ( .A(G22GAT), .B(n425), .ZN(n426) );
  XNOR2_X1 U494 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U495 ( .A(n429), .B(n428), .Z(n432) );
  XNOR2_X1 U496 ( .A(n430), .B(G197GAT), .ZN(n431) );
  XOR2_X1 U497 ( .A(n432), .B(n431), .Z(n504) );
  INV_X1 U498 ( .A(n504), .ZN(n579) );
  XOR2_X1 U499 ( .A(KEYINPUT77), .B(KEYINPUT76), .Z(n434) );
  XNOR2_X1 U500 ( .A(G204GAT), .B(KEYINPUT32), .ZN(n433) );
  XNOR2_X1 U501 ( .A(n434), .B(n433), .ZN(n436) );
  XOR2_X1 U502 ( .A(n436), .B(n435), .Z(n440) );
  XNOR2_X1 U503 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U504 ( .A(n440), .B(n439), .ZN(n449) );
  XOR2_X1 U505 ( .A(KEYINPUT78), .B(KEYINPUT31), .Z(n442) );
  NAND2_X1 U506 ( .A1(G230GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U507 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U508 ( .A(n443), .B(KEYINPUT33), .Z(n447) );
  XNOR2_X1 U509 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U510 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U511 ( .A(n449), .B(n448), .Z(n582) );
  NAND2_X1 U512 ( .A1(n579), .A2(n582), .ZN(n486) );
  NOR2_X1 U513 ( .A1(n519), .A2(n486), .ZN(n450) );
  XNOR2_X1 U514 ( .A(n451), .B(n450), .ZN(n501) );
  NOR2_X1 U515 ( .A1(n536), .A2(n501), .ZN(n454) );
  INV_X1 U516 ( .A(G43GAT), .ZN(n452) );
  XOR2_X1 U517 ( .A(KEYINPUT118), .B(KEYINPUT54), .Z(n469) );
  NOR2_X1 U518 ( .A1(n481), .A2(n591), .ZN(n455) );
  XNOR2_X1 U519 ( .A(KEYINPUT45), .B(n455), .ZN(n456) );
  NAND2_X1 U520 ( .A1(n456), .A2(n582), .ZN(n457) );
  NOR2_X1 U521 ( .A1(n579), .A2(n457), .ZN(n458) );
  XNOR2_X1 U522 ( .A(n458), .B(KEYINPUT109), .ZN(n466) );
  XOR2_X1 U523 ( .A(KEYINPUT108), .B(KEYINPUT47), .Z(n464) );
  XNOR2_X1 U524 ( .A(n582), .B(KEYINPUT41), .ZN(n555) );
  NAND2_X1 U525 ( .A1(n579), .A2(n555), .ZN(n459) );
  XOR2_X1 U526 ( .A(KEYINPUT46), .B(n459), .Z(n460) );
  NOR2_X1 U527 ( .A1(n586), .A2(n460), .ZN(n462) );
  NAND2_X1 U528 ( .A1(n462), .A2(n461), .ZN(n463) );
  XNOR2_X1 U529 ( .A(n464), .B(n463), .ZN(n465) );
  NAND2_X1 U530 ( .A1(n466), .A2(n465), .ZN(n467) );
  NAND2_X1 U531 ( .A1(n533), .A2(n524), .ZN(n468) );
  XNOR2_X1 U532 ( .A(n469), .B(n468), .ZN(n576) );
  NOR2_X1 U533 ( .A1(n470), .A2(n520), .ZN(n471) );
  AND2_X1 U534 ( .A1(n576), .A2(n471), .ZN(n475) );
  XNOR2_X1 U535 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n473) );
  NOR2_X1 U536 ( .A1(n536), .A2(n476), .ZN(n566) );
  NAND2_X1 U537 ( .A1(n566), .A2(n555), .ZN(n480) );
  XOR2_X1 U538 ( .A(KEYINPUT121), .B(KEYINPUT57), .Z(n478) );
  XOR2_X1 U539 ( .A(G176GAT), .B(KEYINPUT56), .Z(n477) );
  XNOR2_X1 U540 ( .A(KEYINPUT34), .B(KEYINPUT97), .ZN(n491) );
  XOR2_X1 U541 ( .A(G1GAT), .B(KEYINPUT96), .Z(n489) );
  NOR2_X1 U542 ( .A1(n481), .A2(n567), .ZN(n482) );
  XNOR2_X1 U543 ( .A(n482), .B(KEYINPUT16), .ZN(n485) );
  INV_X1 U544 ( .A(n483), .ZN(n484) );
  NAND2_X1 U545 ( .A1(n485), .A2(n484), .ZN(n505) );
  NOR2_X1 U546 ( .A1(n486), .A2(n505), .ZN(n487) );
  XOR2_X1 U547 ( .A(KEYINPUT95), .B(n487), .Z(n495) );
  NAND2_X1 U548 ( .A1(n495), .A2(n520), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U550 ( .A(n491), .B(n490), .ZN(G1324GAT) );
  NAND2_X1 U551 ( .A1(n524), .A2(n495), .ZN(n492) );
  XNOR2_X1 U552 ( .A(n492), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U553 ( .A(G15GAT), .B(KEYINPUT35), .Z(n494) );
  NAND2_X1 U554 ( .A1(n495), .A2(n526), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n494), .B(n493), .ZN(G1326GAT) );
  NAND2_X1 U556 ( .A1(n529), .A2(n495), .ZN(n496) );
  XNOR2_X1 U557 ( .A(n496), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U558 ( .A1(n501), .A2(n575), .ZN(n498) );
  XNOR2_X1 U559 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n498), .B(n497), .ZN(G1328GAT) );
  NOR2_X1 U561 ( .A1(n499), .A2(n501), .ZN(n500) );
  XOR2_X1 U562 ( .A(G36GAT), .B(n500), .Z(G1329GAT) );
  XNOR2_X1 U563 ( .A(G50GAT), .B(KEYINPUT99), .ZN(n503) );
  INV_X1 U564 ( .A(n529), .ZN(n538) );
  NOR2_X1 U565 ( .A1(n538), .A2(n501), .ZN(n502) );
  XNOR2_X1 U566 ( .A(n503), .B(n502), .ZN(G1331GAT) );
  XOR2_X1 U567 ( .A(KEYINPUT100), .B(KEYINPUT42), .Z(n507) );
  NAND2_X1 U568 ( .A1(n504), .A2(n555), .ZN(n518) );
  NOR2_X1 U569 ( .A1(n518), .A2(n505), .ZN(n514) );
  NAND2_X1 U570 ( .A1(n514), .A2(n520), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n507), .B(n506), .ZN(n508) );
  XOR2_X1 U572 ( .A(G57GAT), .B(n508), .Z(G1332GAT) );
  XOR2_X1 U573 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n510) );
  NAND2_X1 U574 ( .A1(n514), .A2(n524), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U576 ( .A(G64GAT), .B(n511), .ZN(G1333GAT) );
  XOR2_X1 U577 ( .A(G71GAT), .B(KEYINPUT103), .Z(n513) );
  NAND2_X1 U578 ( .A1(n514), .A2(n526), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n513), .B(n512), .ZN(G1334GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT104), .B(KEYINPUT43), .Z(n516) );
  NAND2_X1 U581 ( .A1(n514), .A2(n529), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U583 ( .A(G78GAT), .B(n517), .ZN(G1335GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n522) );
  NOR2_X1 U585 ( .A1(n519), .A2(n518), .ZN(n530) );
  NAND2_X1 U586 ( .A1(n530), .A2(n520), .ZN(n521) );
  XNOR2_X1 U587 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U588 ( .A(G85GAT), .B(n523), .ZN(G1336GAT) );
  NAND2_X1 U589 ( .A1(n524), .A2(n530), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n525), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U591 ( .A(G99GAT), .B(KEYINPUT107), .Z(n528) );
  NAND2_X1 U592 ( .A1(n530), .A2(n526), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n528), .B(n527), .ZN(G1338GAT) );
  XNOR2_X1 U594 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n532) );
  NAND2_X1 U595 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n532), .B(n531), .ZN(G1339GAT) );
  NAND2_X1 U597 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U598 ( .A(n535), .B(KEYINPUT110), .ZN(n551) );
  NOR2_X1 U599 ( .A1(n536), .A2(n551), .ZN(n537) );
  NAND2_X1 U600 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U601 ( .A(KEYINPUT111), .B(n539), .ZN(n547) );
  NAND2_X1 U602 ( .A1(n579), .A2(n547), .ZN(n540) );
  XNOR2_X1 U603 ( .A(G113GAT), .B(n540), .ZN(G1340GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT49), .B(KEYINPUT112), .Z(n542) );
  NAND2_X1 U605 ( .A1(n547), .A2(n555), .ZN(n541) );
  XNOR2_X1 U606 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U607 ( .A(G120GAT), .B(n543), .ZN(G1341GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT50), .B(KEYINPUT113), .Z(n545) );
  NAND2_X1 U609 ( .A1(n547), .A2(n586), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(n546), .ZN(G1342GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT51), .B(KEYINPUT114), .Z(n549) );
  NAND2_X1 U613 ( .A1(n547), .A2(n567), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U615 ( .A(G134GAT), .B(n550), .ZN(G1343GAT) );
  NOR2_X1 U616 ( .A1(n551), .A2(n578), .ZN(n552) );
  XOR2_X1 U617 ( .A(KEYINPUT115), .B(n552), .Z(n561) );
  NAND2_X1 U618 ( .A1(n561), .A2(n579), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n553), .B(KEYINPUT116), .ZN(n554) );
  XNOR2_X1 U620 ( .A(G141GAT), .B(n554), .ZN(G1344GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n557) );
  NAND2_X1 U622 ( .A1(n561), .A2(n555), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U624 ( .A(G148GAT), .B(n558), .ZN(G1345GAT) );
  NAND2_X1 U625 ( .A1(n586), .A2(n561), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U627 ( .A(G162GAT), .B(KEYINPUT117), .Z(n563) );
  NAND2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(G1347GAT) );
  NAND2_X1 U630 ( .A1(n579), .A2(n566), .ZN(n564) );
  XNOR2_X1 U631 ( .A(G169GAT), .B(n564), .ZN(G1348GAT) );
  NAND2_X1 U632 ( .A1(n586), .A2(n566), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n565), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n568), .B(KEYINPUT58), .ZN(n569) );
  XNOR2_X1 U636 ( .A(G190GAT), .B(n569), .ZN(G1351GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT122), .B(KEYINPUT124), .Z(n571) );
  XNOR2_X1 U638 ( .A(KEYINPUT59), .B(KEYINPUT60), .ZN(n570) );
  XNOR2_X1 U639 ( .A(n571), .B(n570), .ZN(n572) );
  XOR2_X1 U640 ( .A(n572), .B(KEYINPUT125), .Z(n574) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT123), .ZN(n573) );
  XNOR2_X1 U642 ( .A(n574), .B(n573), .ZN(n581) );
  NAND2_X1 U643 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U644 ( .A1(n578), .A2(n577), .ZN(n587) );
  NAND2_X1 U645 ( .A1(n587), .A2(n579), .ZN(n580) );
  XOR2_X1 U646 ( .A(n581), .B(n580), .Z(G1352GAT) );
  XOR2_X1 U647 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n584) );
  INV_X1 U648 ( .A(n587), .ZN(n590) );
  OR2_X1 U649 ( .A1(n590), .A2(n582), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U651 ( .A(G204GAT), .B(n585), .ZN(G1353GAT) );
  XOR2_X1 U652 ( .A(G211GAT), .B(KEYINPUT127), .Z(n589) );
  NAND2_X1 U653 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n589), .B(n588), .ZN(G1354GAT) );
  NOR2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U656 ( .A(KEYINPUT62), .B(n592), .Z(n593) );
  XNOR2_X1 U657 ( .A(G218GAT), .B(n593), .ZN(G1355GAT) );
endmodule

