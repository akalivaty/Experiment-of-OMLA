//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 1 0 1 1 1 1 1 1 1 0 1 1 1 0 0 0 0 0 0 0 1 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 1 1 0 1 1 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:38 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n554, new_n555, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n604, new_n605, new_n608, new_n610, new_n611, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT65), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT66), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  XOR2_X1   g028(.A(KEYINPUT67), .B(KEYINPUT68), .Z(new_n454));
  XNOR2_X1  g029(.A(new_n453), .B(new_n454), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n452), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n456), .A2(G567), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n459), .A2(KEYINPUT69), .ZN(new_n460));
  AND2_X1   g035(.A1(new_n459), .A2(KEYINPUT69), .ZN(new_n461));
  AOI211_X1 g036(.A(new_n460), .B(new_n461), .C1(G2106), .C2(new_n452), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(G125), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI211_X1 g043(.A(G137), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n463), .A2(G101), .A3(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n468), .A2(new_n471), .ZN(G160));
  NOR2_X1   g047(.A1(new_n464), .A2(new_n465), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G136), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n473), .A2(new_n463), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n475), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  INV_X1    g056(.A(KEYINPUT70), .ZN(new_n482));
  NAND2_X1  g057(.A1(KEYINPUT4), .A2(G138), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n484), .B1(new_n464), .B2(new_n465), .ZN(new_n485));
  NAND2_X1  g060(.A1(G102), .A2(G2104), .ZN(new_n486));
  AOI21_X1  g061(.A(G2105), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g062(.A(G126), .B1(new_n464), .B2(new_n465), .ZN(new_n488));
  NAND2_X1  g063(.A1(G114), .A2(G2104), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n463), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  OAI211_X1 g066(.A(G138), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n482), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT3), .ZN(new_n496));
  INV_X1    g071(.A(G2104), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n483), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n486), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n463), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(G126), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n503), .B1(new_n498), .B2(new_n499), .ZN(new_n504));
  INV_X1    g079(.A(new_n489), .ZN(new_n505));
  OAI21_X1  g080(.A(G2105), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n502), .A2(new_n506), .A3(new_n482), .A4(new_n494), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n495), .A2(new_n508), .ZN(G164));
  OR2_X1    g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT72), .A2(G651), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT71), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT71), .A2(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(KEYINPUT6), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n516), .A2(new_n517), .A3(KEYINPUT6), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n521), .A2(G543), .A3(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G50), .ZN(new_n525));
  AND3_X1   g100(.A1(new_n521), .A2(new_n522), .A3(new_n512), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G88), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n515), .A2(new_n525), .A3(new_n527), .ZN(G303));
  INV_X1    g103(.A(G303), .ZN(G166));
  NAND2_X1  g104(.A1(new_n524), .A2(G51), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n526), .A2(G89), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n532), .A2(KEYINPUT7), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(KEYINPUT7), .ZN(new_n534));
  AND2_X1   g109(.A1(G63), .A2(G651), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n533), .A2(new_n534), .B1(new_n512), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n530), .A2(new_n531), .A3(new_n536), .ZN(G286));
  INV_X1    g112(.A(G286), .ZN(G168));
  AOI22_X1  g113(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n514), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT73), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n540), .B(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(G52), .A2(new_n524), .B1(new_n526), .B2(G90), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(G301));
  INV_X1    g119(.A(G301), .ZN(G171));
  AOI22_X1  g120(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(new_n514), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n524), .A2(G43), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n526), .A2(G81), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  AND2_X1   g131(.A1(KEYINPUT74), .A2(G53), .ZN(new_n557));
  NAND4_X1  g132(.A1(new_n521), .A2(G543), .A3(new_n522), .A4(new_n557), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT9), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n526), .A2(G91), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n512), .A2(KEYINPUT75), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT75), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n510), .A2(new_n562), .A3(new_n511), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n564), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n565));
  OAI211_X1 g140(.A(new_n559), .B(new_n560), .C1(new_n514), .C2(new_n565), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT76), .ZN(G299));
  NAND4_X1  g142(.A1(new_n521), .A2(G49), .A3(G543), .A4(new_n522), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n521), .A2(G87), .A3(new_n512), .A4(new_n522), .ZN(new_n569));
  OAI21_X1  g144(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(G288));
  INV_X1    g146(.A(G61), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n572), .B1(new_n510), .B2(new_n511), .ZN(new_n573));
  AND2_X1   g148(.A1(G73), .A2(G543), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n521), .A2(G48), .A3(G543), .A4(new_n522), .ZN(new_n576));
  AND2_X1   g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n521), .A2(G86), .A3(new_n512), .A4(new_n522), .ZN(new_n578));
  AND2_X1   g153(.A1(new_n578), .A2(KEYINPUT77), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n578), .A2(KEYINPUT77), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n577), .B1(new_n579), .B2(new_n580), .ZN(G305));
  XOR2_X1   g156(.A(KEYINPUT79), .B(G85), .Z(new_n582));
  AOI22_X1  g157(.A1(G47), .A2(new_n524), .B1(new_n526), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT80), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n583), .A2(new_n584), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n587), .A2(new_n514), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT78), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n588), .B(new_n589), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n585), .A2(new_n586), .A3(new_n590), .ZN(G290));
  NAND2_X1  g166(.A1(G301), .A2(G868), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n526), .A2(G92), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n593), .B(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n524), .A2(G54), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n564), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n597), .A2(new_n514), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n595), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n592), .B1(new_n600), .B2(G868), .ZN(G284));
  OAI21_X1  g176(.A(new_n592), .B1(new_n600), .B2(G868), .ZN(G321));
  NAND2_X1  g177(.A1(G286), .A2(G868), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT76), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n566), .B(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n603), .B1(new_n605), .B2(G868), .ZN(G297));
  OAI21_X1  g181(.A(new_n603), .B1(new_n605), .B2(G868), .ZN(G280));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n600), .B1(new_n608), .B2(G860), .ZN(G148));
  NAND2_X1  g184(.A1(new_n600), .A2(new_n608), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(G868), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(G868), .B2(new_n551), .ZN(G323));
  XNOR2_X1  g187(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AOI22_X1  g188(.A1(G123), .A2(new_n476), .B1(new_n474), .B2(G135), .ZN(new_n614));
  OAI21_X1  g189(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n615));
  INV_X1    g190(.A(G111), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n615), .A2(KEYINPUT81), .B1(new_n616), .B2(G2105), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(KEYINPUT81), .B2(new_n615), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n614), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(G2096), .Z(new_n620));
  NAND3_X1  g195(.A1(new_n463), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT12), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT13), .ZN(new_n623));
  INV_X1    g198(.A(G2100), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n620), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT82), .ZN(G156));
  XNOR2_X1  g203(.A(G2427), .B(G2438), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2430), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT15), .B(G2435), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n632), .A2(KEYINPUT14), .A3(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(KEYINPUT83), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G1341), .ZN(new_n637));
  INV_X1    g212(.A(G1348), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g214(.A(G1341), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n636), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(G1348), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G2451), .B(G2454), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n645), .B(new_n646), .Z(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n643), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n639), .A2(new_n642), .A3(new_n647), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n649), .A2(G14), .A3(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(G401));
  XNOR2_X1  g227(.A(G2072), .B(G2078), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2067), .B(G2678), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT84), .ZN(new_n655));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT85), .B(KEYINPUT18), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n653), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(new_n658), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n655), .A2(new_n657), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n661), .A2(KEYINPUT17), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n663), .A2(new_n659), .ZN(new_n664));
  MUX2_X1   g239(.A(new_n653), .B(new_n660), .S(new_n664), .Z(new_n665));
  XNOR2_X1  g240(.A(G2096), .B(G2100), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(G227));
  XNOR2_X1  g243(.A(G1971), .B(G1976), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT86), .B(KEYINPUT19), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1956), .B(G2474), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1961), .B(G1966), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n672), .B(new_n673), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n672), .A2(new_n673), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n671), .A2(new_n676), .ZN(new_n677));
  AND2_X1   g252(.A1(new_n677), .A2(KEYINPUT20), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n677), .A2(KEYINPUT20), .ZN(new_n679));
  OAI221_X1 g254(.A(new_n674), .B1(new_n671), .B2(new_n675), .C1(new_n678), .C2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(G1991), .B(G1996), .Z(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n684), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1981), .B(G1986), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n685), .A2(new_n688), .A3(new_n686), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(G229));
  INV_X1    g267(.A(KEYINPUT34), .ZN(new_n693));
  INV_X1    g268(.A(G16), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G23), .ZN(new_n695));
  INV_X1    g270(.A(G288), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(new_n694), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT87), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT33), .B(G1976), .Z(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n697), .A2(KEYINPUT87), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n697), .A2(KEYINPUT87), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n702), .A2(new_n699), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  AND2_X1   g281(.A1(new_n694), .A2(G6), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G305), .B2(G16), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT32), .B(G1981), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(G303), .A2(G16), .ZN(new_n712));
  INV_X1    g287(.A(G22), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n712), .B1(G16), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G1971), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n708), .A2(new_n710), .ZN(new_n716));
  INV_X1    g291(.A(G1971), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n712), .B(new_n717), .C1(G16), .C2(new_n713), .ZN(new_n718));
  NAND4_X1  g293(.A1(new_n711), .A2(new_n715), .A3(new_n716), .A4(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n693), .B1(new_n706), .B2(new_n720), .ZN(new_n721));
  NOR3_X1   g296(.A1(new_n705), .A2(new_n719), .A3(KEYINPUT34), .ZN(new_n722));
  INV_X1    g297(.A(G29), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G25), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n474), .A2(G131), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n476), .A2(G119), .ZN(new_n726));
  OR2_X1    g301(.A1(G95), .A2(G2105), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n727), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n725), .A2(new_n726), .A3(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n724), .B1(new_n730), .B2(new_n723), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT35), .B(G1991), .Z(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n731), .B(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(G290), .A2(G16), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n694), .A2(G24), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n736), .A2(G1986), .A3(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(G1986), .B1(new_n736), .B2(new_n737), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n735), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(KEYINPUT88), .B1(new_n722), .B2(new_n741), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n706), .A2(new_n720), .A3(new_n693), .ZN(new_n743));
  INV_X1    g318(.A(new_n740), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n734), .B1(new_n744), .B2(new_n738), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT88), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n743), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n721), .B1(new_n742), .B2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT36), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n749), .A2(KEYINPUT89), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n748), .B(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(G286), .A2(G16), .ZN(new_n753));
  INV_X1    g328(.A(G1966), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n694), .A2(G21), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n753), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n694), .A2(G5), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G301), .B2(G16), .ZN(new_n758));
  INV_X1    g333(.A(G1961), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n756), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n753), .A2(new_n755), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n761), .A2(G1966), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT96), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(new_n619), .B2(new_n723), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT31), .B(G11), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT30), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n766), .A2(G28), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT97), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n768), .B(new_n723), .C1(new_n766), .C2(G28), .ZN(new_n769));
  AND3_X1   g344(.A1(new_n764), .A2(new_n765), .A3(new_n769), .ZN(new_n770));
  NAND4_X1  g345(.A1(new_n614), .A2(KEYINPUT96), .A3(G29), .A4(new_n618), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n762), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  OR3_X1    g347(.A1(new_n760), .A2(KEYINPUT98), .A3(new_n772), .ZN(new_n773));
  OR2_X1    g348(.A1(G4), .A2(G16), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n599), .B2(new_n694), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G1348), .ZN(new_n776));
  OAI21_X1  g351(.A(KEYINPUT98), .B1(new_n760), .B2(new_n772), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n723), .A2(G27), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G164), .B2(new_n723), .ZN(new_n779));
  INV_X1    g354(.A(G2078), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NAND4_X1  g356(.A1(new_n773), .A2(new_n776), .A3(new_n777), .A4(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n694), .A2(G20), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT23), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(new_n605), .B2(new_n694), .ZN(new_n786));
  INV_X1    g361(.A(G1956), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  AND2_X1   g363(.A1(KEYINPUT24), .A2(G34), .ZN(new_n789));
  NOR2_X1   g364(.A1(KEYINPUT24), .A2(G34), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n723), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT93), .Z(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G29), .B2(G160), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G2084), .ZN(new_n794));
  NOR2_X1   g369(.A1(G29), .A2(G33), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT91), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT92), .B(KEYINPUT25), .ZN(new_n797));
  AND3_X1   g372(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n474), .A2(G139), .ZN(new_n800));
  INV_X1    g375(.A(new_n473), .ZN(new_n801));
  AOI22_X1  g376(.A1(new_n801), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n799), .B(new_n800), .C1(new_n802), .C2(new_n463), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n796), .B1(new_n803), .B2(new_n723), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n804), .A2(G2072), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n804), .A2(G2072), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n794), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n480), .A2(G29), .ZN(new_n808));
  INV_X1    g383(.A(G35), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n808), .B1(G29), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n810), .A2(KEYINPUT29), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT29), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n808), .B(new_n812), .C1(G29), .C2(new_n809), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(G2090), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n723), .A2(G26), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT90), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT28), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n474), .A2(G140), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n476), .A2(G128), .ZN(new_n820));
  OR2_X1    g395(.A1(G104), .A2(G2105), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n821), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n819), .A2(new_n820), .A3(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n818), .B1(new_n824), .B2(new_n723), .ZN(new_n825));
  INV_X1    g400(.A(G2067), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  OR2_X1    g402(.A1(G16), .A2(G19), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(new_n550), .B2(new_n694), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(new_n640), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n807), .A2(new_n815), .A3(new_n827), .A4(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(G2090), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n811), .A2(new_n832), .A3(new_n813), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT99), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n758), .A2(new_n759), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n829), .A2(new_n640), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n723), .A2(G32), .ZN(new_n838));
  NAND3_X1  g413(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT94), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT26), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n474), .A2(G141), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n476), .A2(G129), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n463), .A2(G105), .A3(G2104), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n842), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n838), .B1(new_n847), .B2(new_n723), .ZN(new_n848));
  XNOR2_X1  g423(.A(KEYINPUT27), .B(G1996), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT95), .ZN(new_n850));
  AND2_X1   g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n848), .A2(new_n850), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n836), .B(new_n837), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  NOR3_X1   g428(.A1(new_n831), .A2(new_n835), .A3(new_n853), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n783), .A2(KEYINPUT100), .A3(new_n788), .A4(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT100), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n788), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n856), .B1(new_n857), .B2(new_n782), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  AND2_X1   g434(.A1(new_n752), .A2(new_n859), .ZN(G311));
  AOI21_X1  g435(.A(KEYINPUT101), .B1(new_n752), .B2(new_n859), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n742), .A2(new_n747), .ZN(new_n862));
  INV_X1    g437(.A(new_n721), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n751), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI211_X1 g439(.A(new_n721), .B(new_n750), .C1(new_n742), .C2(new_n747), .ZN(new_n865));
  OAI211_X1 g440(.A(new_n859), .B(KEYINPUT101), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n861), .A2(new_n867), .ZN(G150));
  NAND2_X1  g443(.A1(new_n600), .A2(G559), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT38), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n524), .A2(G55), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n526), .A2(G93), .ZN(new_n872));
  AOI22_X1  g447(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n873));
  OAI211_X1 g448(.A(new_n871), .B(new_n872), .C1(new_n514), .C2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n551), .B(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n870), .B(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT39), .ZN(new_n878));
  AOI21_X1  g453(.A(G860), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n879), .B1(new_n878), .B2(new_n877), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n874), .A2(G860), .ZN(new_n881));
  XOR2_X1   g456(.A(new_n881), .B(KEYINPUT37), .Z(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(new_n882), .ZN(G145));
  NAND2_X1  g458(.A1(new_n476), .A2(G130), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n463), .A2(G118), .ZN(new_n885));
  OAI21_X1  g460(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n884), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n887), .B1(G142), .B2(new_n474), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(new_n622), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(new_n730), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n803), .A2(KEYINPUT102), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(new_n847), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n892), .A2(new_n494), .A3(new_n491), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n892), .B1(new_n494), .B2(new_n491), .ZN(new_n894));
  OR3_X1    g469(.A1(new_n893), .A2(new_n894), .A3(new_n823), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n823), .B1(new_n893), .B2(new_n894), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n890), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n619), .B(G160), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(G162), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n895), .A2(KEYINPUT103), .A3(new_n890), .A4(new_n896), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT103), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n895), .A2(new_n896), .ZN(new_n903));
  INV_X1    g478(.A(new_n890), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n902), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n900), .A2(new_n901), .A3(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(G37), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n903), .A2(new_n904), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n899), .B1(new_n908), .B2(new_n897), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n906), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n910), .B(new_n911), .ZN(G395));
  INV_X1    g487(.A(G868), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n874), .A2(new_n913), .ZN(new_n914));
  XOR2_X1   g489(.A(G290), .B(G305), .Z(new_n915));
  XNOR2_X1  g490(.A(G303), .B(G288), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n915), .B(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(KEYINPUT42), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n610), .B(new_n875), .ZN(new_n919));
  NOR2_X1   g494(.A1(G299), .A2(new_n600), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n605), .A2(new_n599), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n919), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT41), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n924), .B1(new_n920), .B2(new_n921), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n605), .A2(new_n599), .ZN(new_n926));
  NAND2_X1  g501(.A1(G299), .A2(new_n600), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n926), .A2(new_n927), .A3(KEYINPUT41), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n923), .B1(new_n919), .B2(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n918), .B(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n914), .B1(new_n931), .B2(new_n913), .ZN(G295));
  OAI21_X1  g507(.A(new_n914), .B1(new_n931), .B2(new_n913), .ZN(G331));
  NAND2_X1  g508(.A1(G171), .A2(G168), .ZN(new_n934));
  NAND2_X1  g509(.A1(G301), .A2(G286), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n934), .A2(new_n875), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n935), .ZN(new_n937));
  AND3_X1   g512(.A1(new_n937), .A2(KEYINPUT105), .A3(new_n876), .ZN(new_n938));
  AOI21_X1  g513(.A(KEYINPUT105), .B1(new_n937), .B2(new_n876), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n936), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n936), .B1(new_n920), .B2(new_n921), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n937), .A2(new_n876), .ZN(new_n943));
  AOI22_X1  g518(.A1(new_n929), .A2(new_n940), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n917), .ZN(new_n945));
  AOI21_X1  g520(.A(G37), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n929), .A2(new_n940), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n942), .A2(new_n943), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(new_n917), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT43), .B1(new_n946), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n945), .A2(new_n947), .A3(new_n948), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n938), .A2(new_n939), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n953), .A2(new_n941), .ZN(new_n954));
  AOI22_X1  g529(.A1(new_n925), .A2(new_n928), .B1(new_n936), .B2(new_n943), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n917), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AND4_X1   g531(.A1(KEYINPUT43), .A2(new_n952), .A3(new_n956), .A4(new_n907), .ZN(new_n957));
  OAI21_X1  g532(.A(KEYINPUT44), .B1(new_n951), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT44), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT43), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n960), .B1(new_n946), .B2(new_n950), .ZN(new_n961));
  AND4_X1   g536(.A1(new_n960), .A2(new_n952), .A3(new_n956), .A4(new_n907), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n959), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n958), .A2(new_n963), .ZN(G397));
  NAND3_X1  g539(.A1(new_n502), .A2(new_n506), .A3(new_n494), .ZN(new_n965));
  XOR2_X1   g540(.A(KEYINPUT106), .B(G1384), .Z(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT45), .ZN(new_n968));
  INV_X1    g543(.A(G40), .ZN(new_n969));
  NOR3_X1   g544(.A1(new_n468), .A2(new_n471), .A3(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n967), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  XOR2_X1   g546(.A(new_n971), .B(KEYINPUT107), .Z(new_n972));
  XNOR2_X1  g547(.A(new_n823), .B(new_n826), .ZN(new_n973));
  INV_X1    g548(.A(G1996), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n973), .B1(new_n974), .B2(new_n847), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n971), .A2(G1996), .ZN(new_n976));
  AOI22_X1  g551(.A1(new_n972), .A2(new_n975), .B1(new_n847), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n729), .A2(new_n733), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n730), .A2(new_n732), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n972), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  OR2_X1    g556(.A1(G290), .A2(G1986), .ZN(new_n982));
  NAND2_X1  g557(.A1(G290), .A2(G1986), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n971), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  XOR2_X1   g560(.A(new_n985), .B(KEYINPUT108), .Z(new_n986));
  NAND2_X1  g561(.A1(G303), .A2(G8), .ZN(new_n987));
  XNOR2_X1  g562(.A(KEYINPUT110), .B(KEYINPUT55), .ZN(new_n988));
  XOR2_X1   g563(.A(new_n987), .B(new_n988), .Z(new_n989));
  AOI21_X1  g564(.A(G1384), .B1(new_n491), .B2(new_n494), .ZN(new_n990));
  XOR2_X1   g565(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n965), .A2(KEYINPUT70), .ZN(new_n993));
  AOI21_X1  g568(.A(G1384), .B1(new_n993), .B2(new_n507), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT50), .ZN(new_n995));
  OAI211_X1 g570(.A(new_n970), .B(new_n992), .C1(new_n994), .C2(new_n995), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n996), .A2(G2090), .ZN(new_n997));
  INV_X1    g572(.A(G1384), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n998), .B1(new_n495), .B2(new_n508), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(new_n968), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n965), .A2(KEYINPUT45), .A3(new_n966), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n1001), .A2(new_n970), .ZN(new_n1002));
  AOI21_X1  g577(.A(G1971), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  OAI211_X1 g578(.A(G8), .B(new_n989), .C1(new_n997), .C2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G1981), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n577), .B(new_n1005), .C1(new_n579), .C2(new_n580), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT113), .ZN(new_n1007));
  OR2_X1    g582(.A1(new_n578), .A2(KEYINPUT77), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n578), .A2(KEYINPUT77), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT113), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1010), .A2(new_n1011), .A3(new_n1005), .A4(new_n577), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1007), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1005), .B1(new_n577), .B2(new_n578), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT49), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1014), .B1(new_n1007), .B2(new_n1012), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT49), .ZN(new_n1020));
  INV_X1    g595(.A(G8), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1021), .B1(new_n990), .B2(new_n970), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1018), .A2(new_n1020), .A3(new_n1022), .ZN(new_n1023));
  AND2_X1   g598(.A1(new_n569), .A2(new_n570), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1024), .A2(KEYINPUT111), .A3(G1976), .A4(new_n568), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n970), .A2(new_n965), .A3(new_n998), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT111), .ZN(new_n1027));
  INV_X1    g602(.A(G1976), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1027), .B1(G288), .B2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1025), .A2(new_n1026), .A3(new_n1029), .A4(G8), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT52), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT112), .ZN(new_n1032));
  AND4_X1   g607(.A1(G8), .A2(new_n1025), .A3(new_n1026), .A4(new_n1029), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n696), .A2(G1976), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1034), .A2(KEYINPUT52), .ZN(new_n1035));
  AOI22_X1  g610(.A1(new_n1031), .A2(new_n1032), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  NOR4_X1   g611(.A1(new_n1030), .A2(KEYINPUT112), .A3(KEYINPUT52), .A4(new_n1034), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1004), .A2(new_n1023), .A3(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n970), .B1(new_n990), .B2(new_n991), .ZN(new_n1040));
  NOR2_X1   g615(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1042), .B1(new_n993), .B2(new_n507), .ZN(new_n1043));
  OAI21_X1  g618(.A(KEYINPUT115), .B1(new_n1040), .B2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1041), .B1(new_n495), .B2(new_n508), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT115), .ZN(new_n1046));
  NAND2_X1  g621(.A1(G160), .A2(G40), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n965), .A2(new_n998), .ZN(new_n1048));
  INV_X1    g623(.A(new_n991), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1047), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1045), .A2(new_n1046), .A3(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1044), .A2(new_n832), .A3(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1002), .B1(new_n994), .B2(KEYINPUT45), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(new_n717), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n989), .B1(new_n1055), .B2(G8), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1057), .B1(new_n1053), .B2(G2078), .ZN(new_n1058));
  AOI211_X1 g633(.A(new_n968), .B(G1384), .C1(new_n993), .C2(new_n507), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n970), .B1(new_n990), .B2(KEYINPUT45), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n780), .A2(KEYINPUT53), .ZN(new_n1061));
  OR3_X1    g636(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n996), .A2(new_n759), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1058), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(G171), .ZN(new_n1065));
  NOR3_X1   g640(.A1(new_n1039), .A2(new_n1056), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT51), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n754), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1047), .A2(G2084), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n992), .B(new_n1069), .C1(new_n994), .C2(new_n995), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1067), .B1(new_n1071), .B2(G286), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1068), .A2(G168), .A3(new_n1070), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(G8), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1067), .B1(new_n1073), .B2(G8), .ZN(new_n1076));
  OAI21_X1  g651(.A(KEYINPUT62), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1074), .A2(KEYINPUT51), .ZN(new_n1078));
  AOI21_X1  g653(.A(G168), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1079));
  OAI211_X1 g654(.A(G8), .B(new_n1073), .C1(new_n1079), .C2(new_n1067), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT62), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1078), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1066), .A2(new_n1077), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT124), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT124), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1066), .A2(new_n1077), .A3(new_n1085), .A4(new_n1082), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1088));
  INV_X1    g663(.A(new_n471), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1089), .A2(KEYINPUT123), .ZN(new_n1090));
  NOR4_X1   g665(.A1(new_n1090), .A2(new_n969), .A3(new_n468), .A4(new_n1061), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n967), .A2(new_n968), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1089), .A2(KEYINPUT123), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1091), .A2(new_n1092), .A3(new_n1001), .A4(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1058), .A2(new_n1063), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(G171), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1058), .A2(new_n1062), .A3(G301), .A4(new_n1063), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1096), .A2(KEYINPUT54), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1088), .A2(new_n1098), .ZN(new_n1099));
  AND2_X1   g674(.A1(new_n1023), .A2(new_n1038), .ZN(new_n1100));
  INV_X1    g675(.A(new_n989), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1045), .A2(new_n1050), .ZN(new_n1102));
  AOI21_X1  g677(.A(G2090), .B1(new_n1102), .B2(KEYINPUT115), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n1103), .A2(new_n1051), .B1(new_n717), .B2(new_n1053), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1101), .B1(new_n1104), .B2(new_n1021), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1100), .A2(new_n1004), .A3(new_n1105), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1058), .A2(G301), .A3(new_n1063), .A4(new_n1094), .ZN(new_n1107));
  AOI21_X1  g682(.A(KEYINPUT54), .B1(new_n1065), .B2(new_n1107), .ZN(new_n1108));
  NOR3_X1   g683(.A1(new_n1099), .A2(new_n1106), .A3(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1026), .A2(G2067), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1110), .B1(new_n996), .B2(new_n638), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1111), .A2(KEYINPUT60), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT60), .ZN(new_n1113));
  AOI211_X1 g688(.A(new_n1113), .B(new_n1110), .C1(new_n996), .C2(new_n638), .ZN(new_n1114));
  NOR3_X1   g689(.A1(new_n1112), .A2(new_n1114), .A3(new_n599), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1111), .A2(KEYINPUT60), .A3(new_n599), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT59), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1002), .B(new_n974), .C1(new_n994), .C2(KEYINPUT45), .ZN(new_n1118));
  XOR2_X1   g693(.A(KEYINPUT58), .B(G1341), .Z(new_n1119));
  NAND2_X1  g694(.A1(new_n1026), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1117), .B1(new_n1121), .B2(new_n551), .ZN(new_n1122));
  AOI211_X1 g697(.A(KEYINPUT59), .B(new_n550), .C1(new_n1118), .C2(new_n1120), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1116), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1115), .A2(new_n1124), .ZN(new_n1125));
  XNOR2_X1  g700(.A(KEYINPUT56), .B(G2072), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1002), .B(new_n1126), .C1(new_n994), .C2(KEYINPUT45), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(KEYINPUT121), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT121), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1000), .A2(new_n1129), .A3(new_n1002), .A4(new_n1126), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g706(.A(KEYINPUT118), .B(G1956), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1102), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT119), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n566), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1136), .A2(KEYINPUT120), .A3(KEYINPUT57), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT120), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1138), .B1(new_n566), .B2(new_n1135), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT57), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1140), .B1(new_n566), .B2(new_n1138), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1137), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1134), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1131), .A2(new_n1142), .A3(new_n1133), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1144), .A2(KEYINPUT61), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT61), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1131), .A2(new_n1133), .A3(new_n1142), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1142), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1147), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  AND3_X1   g725(.A1(new_n1125), .A2(new_n1146), .A3(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1111), .A2(new_n599), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1145), .B1(new_n1149), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(KEYINPUT122), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT122), .ZN(new_n1155));
  OAI211_X1 g730(.A(new_n1155), .B(new_n1145), .C1(new_n1149), .C2(new_n1152), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1109), .B1(new_n1151), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1087), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n999), .A2(KEYINPUT50), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1160), .A2(new_n832), .A3(new_n970), .A4(new_n992), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1021), .B1(new_n1161), .B2(new_n1054), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1101), .B1(new_n1162), .B2(KEYINPUT116), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT116), .ZN(new_n1164));
  AOI211_X1 g739(.A(new_n1164), .B(new_n1021), .C1(new_n1161), .C2(new_n1054), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g741(.A1(G286), .A2(new_n1021), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1023), .A2(new_n1038), .A3(new_n1071), .A4(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(KEYINPUT63), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n1022), .B(KEYINPUT114), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1022), .B1(new_n1019), .B2(KEYINPUT49), .ZN(new_n1171));
  AOI211_X1 g746(.A(new_n1017), .B(new_n1014), .C1(new_n1007), .C2(new_n1012), .ZN(new_n1172));
  OAI211_X1 g747(.A(new_n1028), .B(new_n696), .C1(new_n1171), .C2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1170), .B1(new_n1173), .B2(new_n1013), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT63), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1071), .A2(new_n1175), .A3(new_n1167), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1004), .B1(new_n1056), .B2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1174), .B1(new_n1177), .B2(new_n1100), .ZN(new_n1178));
  AND3_X1   g753(.A1(new_n1169), .A2(new_n1178), .A3(KEYINPUT117), .ZN(new_n1179));
  AOI21_X1  g754(.A(KEYINPUT117), .B1(new_n1169), .B2(new_n1178), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n986), .B1(new_n1159), .B2(new_n1181), .ZN(new_n1182));
  XOR2_X1   g757(.A(new_n976), .B(KEYINPUT46), .Z(new_n1183));
  INV_X1    g758(.A(new_n972), .ZN(new_n1184));
  AND2_X1   g759(.A1(new_n973), .A2(new_n847), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1183), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n1186), .B(KEYINPUT47), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n982), .A2(new_n971), .ZN(new_n1188));
  XNOR2_X1  g763(.A(new_n1188), .B(KEYINPUT48), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1187), .B1(new_n981), .B2(new_n1189), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n978), .B(KEYINPUT125), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n977), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n824), .A2(new_n826), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1184), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT126), .ZN(new_n1195));
  AND2_X1   g770(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1197));
  NOR3_X1   g772(.A1(new_n1190), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1182), .A2(new_n1198), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g774(.A1(new_n961), .A2(new_n962), .ZN(new_n1201));
  NAND2_X1  g775(.A1(new_n667), .A2(G319), .ZN(new_n1202));
  AOI21_X1  g776(.A(new_n1202), .B1(new_n690), .B2(new_n691), .ZN(new_n1203));
  AND3_X1   g777(.A1(new_n1203), .A2(KEYINPUT127), .A3(new_n651), .ZN(new_n1204));
  AOI21_X1  g778(.A(KEYINPUT127), .B1(new_n1203), .B2(new_n651), .ZN(new_n1205));
  OAI21_X1  g779(.A(new_n910), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  NOR2_X1   g780(.A1(new_n1201), .A2(new_n1206), .ZN(G308));
  OAI221_X1 g781(.A(new_n910), .B1(new_n1204), .B2(new_n1205), .C1(new_n961), .C2(new_n962), .ZN(G225));
endmodule


