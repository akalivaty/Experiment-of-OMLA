//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 0 0 0 0 1 1 1 1 1 1 1 0 0 1 1 1 0 1 0 0 1 0 1 0 0 1 1 0 1 0 0 1 0 0 1 0 0 0 0 1 1 0 1 1 0 0 0 1 1 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:26 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XOR2_X1   g002(.A(KEYINPUT2), .B(G113), .Z(new_n189));
  XOR2_X1   g003(.A(G116), .B(G119), .Z(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G107), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(G104), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT3), .ZN(new_n195));
  INV_X1    g009(.A(G104), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(G107), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n194), .B1(new_n195), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT77), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n199), .B1(new_n197), .B2(new_n195), .ZN(new_n200));
  OAI211_X1 g014(.A(KEYINPUT77), .B(KEYINPUT3), .C1(new_n196), .C2(G107), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n198), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT78), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n198), .A2(new_n200), .A3(KEYINPUT78), .A4(new_n201), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(G101), .A3(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT4), .ZN(new_n207));
  AND2_X1   g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G101), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n198), .A2(new_n200), .A3(new_n209), .A4(new_n201), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n207), .B1(new_n206), .B2(new_n210), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n192), .B1(new_n208), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT5), .ZN(new_n213));
  INV_X1    g027(.A(G119), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(new_n214), .A3(G116), .ZN(new_n215));
  OAI211_X1 g029(.A(G113), .B(new_n215), .C1(new_n190), .C2(new_n213), .ZN(new_n216));
  INV_X1    g030(.A(new_n189), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n216), .B1(new_n217), .B2(new_n190), .ZN(new_n218));
  OAI21_X1  g032(.A(G101), .B1(new_n194), .B2(new_n197), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n210), .A2(new_n219), .ZN(new_n220));
  OR2_X1    g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n212), .A2(new_n221), .ZN(new_n222));
  XOR2_X1   g036(.A(G110), .B(G122), .Z(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n223), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n212), .A2(new_n221), .A3(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n224), .A2(KEYINPUT6), .A3(new_n226), .ZN(new_n227));
  XNOR2_X1  g041(.A(G143), .B(G146), .ZN(new_n228));
  NAND2_X1  g042(.A1(KEYINPUT0), .A2(G128), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  XOR2_X1   g044(.A(KEYINPUT0), .B(G128), .Z(new_n231));
  OAI21_X1  g045(.A(new_n230), .B1(new_n228), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G125), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(KEYINPUT82), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT1), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n228), .A2(new_n236), .A3(G128), .ZN(new_n237));
  INV_X1    g051(.A(G146), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n236), .B1(G143), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G128), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n237), .B1(new_n241), .B2(new_n228), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G125), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  OR3_X1    g059(.A1(new_n232), .A2(KEYINPUT82), .A3(new_n244), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n235), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  XOR2_X1   g061(.A(KEYINPUT83), .B(G224), .Z(new_n248));
  INV_X1    g062(.A(G953), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(new_n250), .B(KEYINPUT84), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n247), .A2(new_n252), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n235), .A2(new_n251), .A3(new_n245), .A4(new_n246), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n255), .B(KEYINPUT85), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT6), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n222), .A2(new_n257), .A3(new_n223), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n227), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  AOI22_X1  g073(.A1(new_n245), .A2(new_n234), .B1(new_n251), .B2(KEYINPUT7), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n218), .B(new_n220), .ZN(new_n261));
  XOR2_X1   g075(.A(new_n223), .B(KEYINPUT8), .Z(new_n262));
  AOI21_X1  g076(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT7), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n226), .B(new_n263), .C1(new_n264), .C2(new_n254), .ZN(new_n265));
  INV_X1    g079(.A(G902), .ZN(new_n266));
  AND2_X1   g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n259), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(G210), .B1(G237), .B2(G902), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n259), .A2(new_n267), .A3(new_n269), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n188), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(G475), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT17), .ZN(new_n275));
  INV_X1    g089(.A(G237), .ZN(new_n276));
  AND4_X1   g090(.A1(G143), .A2(new_n276), .A3(new_n249), .A4(G214), .ZN(new_n277));
  NOR2_X1   g091(.A1(G237), .A2(G953), .ZN(new_n278));
  AOI21_X1  g092(.A(G143), .B1(new_n278), .B2(G214), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G131), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT88), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n276), .A2(new_n249), .A3(G214), .ZN(new_n284));
  INV_X1    g098(.A(G143), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n278), .A2(G143), .A3(G214), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n283), .B1(new_n288), .B2(G131), .ZN(new_n289));
  AOI211_X1 g103(.A(KEYINPUT88), .B(new_n281), .C1(new_n286), .C2(new_n287), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n275), .B(new_n282), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G140), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G125), .ZN(new_n293));
  OAI21_X1  g107(.A(KEYINPUT72), .B1(new_n293), .B2(KEYINPUT16), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n244), .A2(G140), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT72), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT16), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n244), .A2(G140), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n293), .A2(new_n299), .A3(KEYINPUT16), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n294), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n238), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n294), .A2(new_n298), .A3(new_n300), .A4(G146), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(G131), .B1(new_n277), .B2(new_n279), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT88), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n288), .A2(new_n283), .A3(G131), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n307), .A2(KEYINPUT17), .A3(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n291), .A2(new_n305), .A3(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(G113), .B(G122), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n311), .B(new_n196), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT87), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n286), .A2(new_n313), .A3(new_n287), .ZN(new_n314));
  NAND2_X1  g128(.A1(KEYINPUT18), .A2(G131), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n314), .B(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n293), .A2(new_n299), .A3(new_n238), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n292), .A2(G125), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT86), .B1(new_n295), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT86), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n293), .A2(new_n299), .A3(new_n320), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n317), .B1(new_n322), .B2(new_n238), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n316), .A2(new_n323), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n310), .A2(new_n312), .A3(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n282), .B1(new_n289), .B2(new_n290), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT19), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n327), .B1(new_n319), .B2(new_n321), .ZN(new_n328));
  NOR3_X1   g142(.A1(new_n295), .A2(new_n318), .A3(KEYINPUT19), .ZN(new_n329));
  OR2_X1    g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n326), .B(new_n303), .C1(new_n330), .C2(G146), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n312), .B1(new_n331), .B2(new_n324), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n274), .B(new_n266), .C1(new_n325), .C2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT89), .ZN(new_n334));
  INV_X1    g148(.A(new_n312), .ZN(new_n335));
  AOI22_X1  g149(.A1(new_n307), .A2(new_n308), .B1(new_n281), .B2(new_n280), .ZN(new_n336));
  NOR3_X1   g150(.A1(new_n328), .A2(G146), .A3(new_n329), .ZN(new_n337));
  INV_X1    g151(.A(new_n303), .ZN(new_n338));
  NOR3_X1   g152(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n324), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n335), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n310), .A2(new_n312), .A3(new_n324), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n334), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n333), .B1(KEYINPUT20), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(KEYINPUT89), .B1(new_n325), .B2(new_n332), .ZN(new_n345));
  AOI21_X1  g159(.A(G475), .B1(new_n341), .B2(new_n342), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT20), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n345), .A2(new_n346), .A3(new_n347), .A4(new_n266), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n310), .A2(new_n324), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n335), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n342), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n274), .B1(new_n352), .B2(new_n266), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(KEYINPUT90), .B1(new_n349), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT90), .ZN(new_n356));
  AOI211_X1 g170(.A(new_n356), .B(new_n353), .C1(new_n344), .C2(new_n348), .ZN(new_n357));
  XNOR2_X1  g171(.A(G116), .B(G122), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n193), .ZN(new_n359));
  INV_X1    g173(.A(G116), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n360), .A2(KEYINPUT14), .A3(G122), .ZN(new_n361));
  INV_X1    g175(.A(new_n358), .ZN(new_n362));
  OAI211_X1 g176(.A(G107), .B(new_n361), .C1(new_n362), .C2(KEYINPUT14), .ZN(new_n363));
  XNOR2_X1  g177(.A(G128), .B(G143), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT92), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n364), .B(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(G134), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n366), .A2(new_n367), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n359), .B(new_n363), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n366), .A2(new_n367), .ZN(new_n371));
  XOR2_X1   g185(.A(KEYINPUT91), .B(KEYINPUT13), .Z(new_n372));
  NAND3_X1  g186(.A1(new_n372), .A2(G128), .A3(new_n285), .ZN(new_n373));
  INV_X1    g187(.A(new_n364), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n373), .B(G134), .C1(new_n372), .C2(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n358), .B(new_n193), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n371), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  XOR2_X1   g191(.A(KEYINPUT9), .B(G234), .Z(new_n378));
  XOR2_X1   g192(.A(KEYINPUT71), .B(G217), .Z(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(new_n379), .A3(new_n249), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n370), .A2(new_n377), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n381), .B1(new_n370), .B2(new_n377), .ZN(new_n383));
  OR2_X1    g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n266), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT15), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(new_n386), .A3(G478), .ZN(new_n387));
  INV_X1    g201(.A(G478), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n384), .B(new_n266), .C1(KEYINPUT15), .C2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G952), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n390), .A2(G953), .ZN(new_n391));
  NAND2_X1  g205(.A1(G234), .A2(G237), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n393), .B(KEYINPUT93), .ZN(new_n394));
  XNOR2_X1  g208(.A(KEYINPUT21), .B(G898), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n395), .A2(G902), .A3(G953), .A4(new_n392), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  XOR2_X1   g211(.A(new_n397), .B(KEYINPUT94), .Z(new_n398));
  NAND3_X1  g212(.A1(new_n387), .A2(new_n389), .A3(new_n398), .ZN(new_n399));
  NOR3_X1   g213(.A1(new_n355), .A2(new_n357), .A3(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(G221), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n401), .B1(new_n378), .B2(new_n266), .ZN(new_n402));
  INV_X1    g216(.A(G469), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n403), .A2(new_n266), .ZN(new_n404));
  XOR2_X1   g218(.A(new_n232), .B(KEYINPUT68), .Z(new_n405));
  OAI21_X1  g219(.A(new_n405), .B1(new_n208), .B2(new_n211), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT11), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n407), .B1(new_n367), .B2(G137), .ZN(new_n408));
  INV_X1    g222(.A(G137), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n409), .A2(KEYINPUT11), .A3(G134), .ZN(new_n410));
  AND2_X1   g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(KEYINPUT64), .B1(new_n409), .B2(G134), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT64), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n413), .A2(new_n367), .A3(G137), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n281), .B1(new_n411), .B2(new_n415), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n415), .A2(new_n281), .A3(new_n408), .A4(new_n410), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT65), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n411), .A2(KEYINPUT65), .A3(new_n281), .A4(new_n415), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n416), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n228), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n239), .A2(KEYINPUT80), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(G128), .B1(new_n239), .B2(KEYINPUT80), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n422), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT79), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n237), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n228), .A2(KEYINPUT79), .A3(new_n236), .A4(G128), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n426), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n220), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT10), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n431), .A2(KEYINPUT10), .A3(new_n242), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n406), .A2(new_n421), .A3(new_n434), .A4(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n249), .A2(G227), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n437), .B(KEYINPUT76), .ZN(new_n438));
  XNOR2_X1  g252(.A(G110), .B(G140), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n438), .B(new_n439), .ZN(new_n440));
  AND2_X1   g254(.A1(new_n436), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n406), .A2(new_n434), .A3(new_n435), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n419), .A2(new_n420), .ZN(new_n443));
  INV_X1    g257(.A(new_n416), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT12), .ZN(new_n447));
  OR2_X1    g261(.A1(new_n447), .A2(KEYINPUT81), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(KEYINPUT81), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n242), .B1(new_n210), .B2(new_n219), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n450), .B1(new_n431), .B2(new_n430), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n448), .B(new_n449), .C1(new_n451), .C2(new_n421), .ZN(new_n452));
  INV_X1    g266(.A(new_n450), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n432), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n454), .A2(KEYINPUT81), .A3(new_n447), .A4(new_n445), .ZN(new_n455));
  AND2_X1   g269(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n436), .ZN(new_n457));
  INV_X1    g271(.A(new_n440), .ZN(new_n458));
  AOI22_X1  g272(.A1(new_n441), .A2(new_n446), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n404), .B1(new_n459), .B2(G469), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n440), .B1(new_n446), .B2(new_n436), .ZN(new_n461));
  AND3_X1   g275(.A1(new_n456), .A2(new_n436), .A3(new_n440), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n403), .B(new_n266), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n402), .B1(new_n460), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n273), .A2(new_n400), .A3(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT95), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n273), .A2(new_n400), .A3(new_n464), .A4(KEYINPUT95), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n278), .A2(G210), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n469), .B(new_n209), .ZN(new_n470));
  XNOR2_X1  g284(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n471));
  XOR2_X1   g285(.A(new_n470), .B(new_n471), .Z(new_n472));
  NAND3_X1  g286(.A1(new_n445), .A2(KEYINPUT66), .A3(new_n232), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT66), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n474), .B1(new_n421), .B2(new_n233), .ZN(new_n475));
  AND2_X1   g289(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n409), .A2(G134), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n367), .A2(G137), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n281), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(KEYINPUT67), .B1(new_n443), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT67), .ZN(new_n483));
  AOI211_X1 g297(.A(new_n483), .B(new_n479), .C1(new_n419), .C2(new_n420), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n482), .A2(new_n485), .A3(new_n242), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n191), .B1(new_n476), .B2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(KEYINPUT69), .B1(new_n443), .B2(new_n480), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT69), .ZN(new_n489));
  AOI211_X1 g303(.A(new_n489), .B(new_n479), .C1(new_n419), .C2(new_n420), .ZN(new_n490));
  NOR3_X1   g304(.A1(new_n488), .A2(new_n490), .A3(new_n243), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n405), .A2(new_n445), .ZN(new_n492));
  NOR3_X1   g306(.A1(new_n491), .A2(new_n492), .A3(new_n192), .ZN(new_n493));
  OAI21_X1  g307(.A(KEYINPUT28), .B1(new_n487), .B2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT70), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n495), .B1(new_n493), .B2(KEYINPUT28), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT29), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n443), .A2(new_n480), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n489), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n443), .A2(KEYINPUT69), .A3(new_n480), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n499), .A2(new_n242), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n405), .A2(new_n445), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n501), .A2(new_n191), .A3(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT28), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n503), .A2(KEYINPUT70), .A3(new_n504), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n494), .A2(new_n496), .A3(new_n497), .A4(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n192), .B1(new_n491), .B2(new_n492), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n504), .B1(new_n507), .B2(new_n503), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n503), .A2(KEYINPUT70), .A3(new_n504), .ZN(new_n509));
  AOI21_X1  g323(.A(KEYINPUT70), .B1(new_n503), .B2(new_n504), .ZN(new_n510));
  NOR3_X1   g324(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n472), .B(new_n506), .C1(new_n511), .C2(new_n497), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT30), .ZN(new_n513));
  NOR3_X1   g327(.A1(new_n481), .A2(new_n484), .A3(new_n243), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n473), .A2(new_n475), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n501), .A2(KEYINPUT30), .A3(new_n502), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(new_n192), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n503), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n519), .A2(new_n472), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n497), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n512), .A2(new_n266), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(G472), .ZN(new_n523));
  NOR2_X1   g337(.A1(G472), .A2(G902), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n518), .A2(new_n503), .A3(new_n472), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT31), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT31), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n518), .A2(new_n527), .A3(new_n503), .A4(new_n472), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n509), .A2(new_n510), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n472), .B1(new_n530), .B2(new_n494), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n524), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT32), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n192), .B1(new_n514), .B2(new_n515), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n504), .B1(new_n535), .B2(new_n503), .ZN(new_n536));
  NOR3_X1   g350(.A1(new_n536), .A2(new_n509), .A3(new_n510), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n526), .B(new_n528), .C1(new_n537), .C2(new_n472), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n538), .A2(KEYINPUT32), .A3(new_n524), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n523), .A2(new_n534), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n240), .A2(G119), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n214), .A2(G128), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT24), .B(G110), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(G110), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n542), .A2(KEYINPUT23), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n541), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n240), .A2(KEYINPUT23), .A3(G119), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n546), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AOI211_X1 g364(.A(new_n545), .B(new_n550), .C1(new_n302), .C2(new_n303), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n548), .A2(new_n549), .ZN(new_n553));
  XNOR2_X1  g367(.A(KEYINPUT73), .B(G110), .ZN(new_n554));
  AOI22_X1  g368(.A1(new_n553), .A2(new_n554), .B1(new_n543), .B2(new_n544), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n303), .A2(new_n317), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(KEYINPUT22), .B(G137), .ZN(new_n559));
  INV_X1    g373(.A(G234), .ZN(new_n560));
  NOR3_X1   g374(.A1(new_n401), .A2(new_n560), .A3(G953), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n559), .B(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n552), .A2(new_n558), .A3(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n562), .B1(new_n551), .B2(new_n557), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n564), .A2(new_n565), .A3(new_n266), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(KEYINPUT74), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT25), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT74), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n564), .A2(new_n565), .A3(new_n569), .A4(new_n266), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n567), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT75), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n564), .A2(new_n565), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n574), .A2(KEYINPUT25), .A3(new_n266), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n567), .A2(KEYINPUT75), .A3(new_n568), .A4(new_n570), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n573), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n379), .B1(new_n560), .B2(G902), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n579), .A2(G902), .ZN(new_n580));
  AOI22_X1  g394(.A1(new_n577), .A2(new_n579), .B1(new_n574), .B2(new_n580), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n467), .A2(new_n468), .A3(new_n540), .A4(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(G101), .ZN(G3));
  NAND2_X1  g397(.A1(new_n460), .A2(new_n463), .ZN(new_n584));
  INV_X1    g398(.A(new_n402), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n532), .ZN(new_n587));
  INV_X1    g401(.A(G472), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n588), .B1(new_n538), .B2(new_n266), .ZN(new_n589));
  NOR3_X1   g403(.A1(new_n586), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n382), .A2(new_n383), .ZN(new_n591));
  AND2_X1   g405(.A1(KEYINPUT96), .A2(KEYINPUT33), .ZN(new_n592));
  NOR2_X1   g406(.A1(KEYINPUT96), .A2(KEYINPUT33), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n592), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n595), .B1(new_n382), .B2(new_n383), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n594), .A2(G478), .A3(new_n266), .A4(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n385), .A2(new_n388), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n349), .A2(new_n354), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n356), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n349), .A2(KEYINPUT90), .A3(new_n354), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n600), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n398), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n590), .A2(new_n273), .A3(new_n581), .A4(new_n606), .ZN(new_n607));
  XOR2_X1   g421(.A(new_n607), .B(KEYINPUT97), .Z(new_n608));
  XNOR2_X1  g422(.A(KEYINPUT34), .B(G104), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(G6));
  XNOR2_X1  g424(.A(new_n333), .B(new_n347), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n611), .A2(new_n353), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n387), .A2(new_n389), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g428(.A(new_n398), .B(KEYINPUT98), .Z(new_n615));
  AND3_X1   g429(.A1(new_n273), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n590), .A2(new_n616), .A3(new_n581), .ZN(new_n617));
  XOR2_X1   g431(.A(KEYINPUT35), .B(G107), .Z(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G9));
  NOR2_X1   g433(.A1(new_n587), .A2(new_n589), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n577), .A2(new_n579), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n552), .A2(new_n558), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n562), .A2(KEYINPUT36), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n580), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n467), .A2(new_n468), .A3(new_n620), .A4(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT37), .B(G110), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G12));
  AND2_X1   g443(.A1(new_n464), .A2(new_n626), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n534), .A2(new_n539), .ZN(new_n631));
  INV_X1    g445(.A(new_n472), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n191), .B1(new_n501), .B2(new_n502), .ZN(new_n633));
  OAI21_X1  g447(.A(KEYINPUT28), .B1(new_n493), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n634), .A2(new_n496), .A3(new_n505), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n632), .B1(new_n635), .B2(KEYINPUT29), .ZN(new_n636));
  AOI22_X1  g450(.A1(new_n636), .A2(new_n506), .B1(new_n497), .B2(new_n520), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n588), .B1(new_n637), .B2(new_n266), .ZN(new_n638));
  OAI211_X1 g452(.A(new_n630), .B(new_n273), .C1(new_n631), .C2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(G900), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n392), .A2(new_n640), .A3(G902), .A4(G953), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(KEYINPUT99), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n394), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(new_n643), .B(KEYINPUT100), .Z(new_n644));
  NAND2_X1  g458(.A1(new_n614), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n639), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(new_n240), .ZN(G30));
  XOR2_X1   g461(.A(new_n644), .B(KEYINPUT39), .Z(new_n648));
  NOR2_X1   g462(.A1(new_n586), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(new_n649), .B(KEYINPUT101), .Z(new_n650));
  INV_X1    g464(.A(KEYINPUT40), .ZN(new_n651));
  OR2_X1    g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n519), .A2(new_n472), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n493), .A2(new_n633), .ZN(new_n654));
  AOI21_X1  g468(.A(G902), .B1(new_n654), .B2(new_n632), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n588), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n631), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n657), .A2(new_n626), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n271), .A2(new_n272), .ZN(new_n659));
  XOR2_X1   g473(.A(new_n659), .B(KEYINPUT38), .Z(new_n660));
  NAND2_X1  g474(.A1(new_n602), .A2(new_n603), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n613), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n660), .A2(new_n188), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n650), .A2(new_n651), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n652), .A2(new_n658), .A3(new_n663), .A4(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G143), .ZN(G45));
  INV_X1    g480(.A(KEYINPUT103), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT102), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n661), .A2(new_n668), .A3(new_n599), .A4(new_n644), .ZN(new_n669));
  OAI211_X1 g483(.A(new_n599), .B(new_n644), .C1(new_n355), .C2(new_n357), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(KEYINPUT102), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n667), .B1(new_n639), .B2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n273), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n538), .A2(KEYINPUT32), .A3(new_n524), .ZN(new_n675));
  AOI21_X1  g489(.A(KEYINPUT32), .B1(new_n538), .B2(new_n524), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n674), .B1(new_n677), .B2(new_n523), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n669), .A2(new_n671), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n678), .A2(KEYINPUT103), .A3(new_n630), .A4(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n673), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G146), .ZN(G48));
  NOR2_X1   g496(.A1(new_n461), .A2(new_n462), .ZN(new_n683));
  OAI21_X1  g497(.A(G469), .B1(new_n683), .B2(G902), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n463), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n402), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n686), .A2(new_n273), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n687), .A2(new_n540), .A3(new_n581), .A4(new_n606), .ZN(new_n688));
  XNOR2_X1  g502(.A(KEYINPUT41), .B(G113), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G15));
  NAND4_X1  g504(.A1(new_n616), .A2(new_n540), .A3(new_n581), .A4(new_n686), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G116), .ZN(G18));
  NAND4_X1  g506(.A1(new_n687), .A2(new_n540), .A3(new_n400), .A4(new_n626), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G119), .ZN(G21));
  XNOR2_X1  g508(.A(new_n589), .B(KEYINPUT104), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n511), .A2(new_n472), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n524), .B1(new_n696), .B2(new_n529), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n695), .A2(new_n581), .A3(new_n615), .A4(new_n697), .ZN(new_n698));
  AOI21_X1  g512(.A(KEYINPUT105), .B1(new_n661), .B2(new_n613), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n661), .A2(KEYINPUT105), .A3(new_n613), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n687), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  OR2_X1    g516(.A1(new_n698), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G122), .ZN(G24));
  OAI21_X1  g518(.A(new_n266), .B1(new_n529), .B2(new_n531), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(G472), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(KEYINPUT104), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT104), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n589), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n707), .A2(new_n626), .A3(new_n709), .A4(new_n697), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n686), .A2(new_n273), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n669), .A2(new_n671), .A3(KEYINPUT106), .ZN(new_n713));
  AOI21_X1  g527(.A(KEYINPUT106), .B1(new_n669), .B2(new_n671), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT107), .B(G125), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G27));
  INV_X1    g532(.A(KEYINPUT108), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n719), .A2(KEYINPUT42), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n713), .A2(new_n714), .A3(new_n720), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n659), .A2(new_n188), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n540), .A2(new_n464), .A3(new_n722), .A4(new_n581), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n719), .A2(KEYINPUT42), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n721), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(new_n725), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT106), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n672), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n669), .A2(new_n671), .A3(KEYINPUT106), .ZN(new_n730));
  INV_X1    g544(.A(new_n720), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n729), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n727), .B1(new_n732), .B2(new_n723), .ZN(new_n733));
  AND2_X1   g547(.A1(new_n726), .A2(new_n733), .ZN(new_n734));
  XOR2_X1   g548(.A(KEYINPUT109), .B(G131), .Z(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(G33));
  AND3_X1   g550(.A1(new_n540), .A2(new_n581), .A3(new_n722), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT110), .ZN(new_n738));
  INV_X1    g552(.A(new_n645), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n737), .A2(new_n738), .A3(new_n464), .A4(new_n739), .ZN(new_n740));
  OAI21_X1  g554(.A(KEYINPUT110), .B1(new_n723), .B2(new_n645), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G134), .ZN(G36));
  INV_X1    g557(.A(new_n661), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n599), .ZN(new_n745));
  OR2_X1    g559(.A1(new_n745), .A2(KEYINPUT43), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(KEYINPUT43), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AOI22_X1  g562(.A1(new_n748), .A2(KEYINPUT111), .B1(new_n621), .B2(new_n625), .ZN(new_n749));
  OAI221_X1 g563(.A(new_n749), .B1(KEYINPUT111), .B2(new_n748), .C1(new_n587), .C2(new_n589), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT44), .ZN(new_n751));
  OR2_X1    g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n722), .B(KEYINPUT112), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT45), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n459), .B(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(G469), .ZN(new_n757));
  INV_X1    g571(.A(new_n404), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n757), .A2(KEYINPUT46), .A3(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT46), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n760), .B(G469), .C1(new_n756), .C2(G902), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n759), .A2(new_n463), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n585), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n763), .A2(new_n648), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n750), .A2(new_n751), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n752), .A2(new_n754), .A3(new_n765), .A4(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G137), .ZN(G39));
  NAND2_X1  g582(.A1(new_n763), .A2(KEYINPUT47), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT47), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n762), .A2(new_n770), .A3(new_n585), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n769), .A2(new_n679), .A3(new_n722), .A4(new_n771), .ZN(new_n772));
  OR3_X1    g586(.A1(new_n772), .A2(new_n540), .A3(new_n581), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G140), .ZN(G42));
  AND2_X1   g588(.A1(new_n685), .A2(KEYINPUT49), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n685), .A2(KEYINPUT49), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n775), .A2(new_n745), .A3(new_n776), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n581), .A2(new_n187), .A3(new_n585), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n777), .A2(new_n660), .A3(new_n657), .A4(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT51), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT50), .ZN(new_n781));
  INV_X1    g595(.A(new_n394), .ZN(new_n782));
  AND3_X1   g596(.A1(new_n746), .A2(new_n782), .A3(new_n747), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n707), .A2(new_n697), .A3(new_n709), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n783), .A2(new_n581), .A3(new_n686), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n660), .A2(new_n188), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n781), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n785), .A2(new_n581), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n789), .A2(new_n748), .A3(new_n394), .ZN(new_n790));
  INV_X1    g604(.A(new_n787), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n790), .A2(KEYINPUT50), .A3(new_n686), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n788), .A2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n581), .A2(new_n782), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n722), .A2(new_n686), .ZN(new_n796));
  NOR4_X1   g610(.A1(new_n795), .A2(new_n796), .A3(new_n631), .A4(new_n656), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n797), .A2(new_n744), .A3(new_n600), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n748), .A2(new_n394), .A3(new_n796), .ZN(new_n799));
  INV_X1    g613(.A(new_n710), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR4_X1   g615(.A1(new_n789), .A2(new_n748), .A3(new_n753), .A4(new_n394), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n685), .A2(new_n585), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n804), .B1(new_n769), .B2(new_n771), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n798), .B(new_n801), .C1(new_n803), .C2(new_n805), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n780), .B1(new_n794), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n790), .A2(new_n687), .ZN(new_n808));
  INV_X1    g622(.A(new_n805), .ZN(new_n809));
  AOI22_X1  g623(.A1(new_n809), .A2(new_n802), .B1(new_n800), .B2(new_n799), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n810), .A2(new_n793), .A3(KEYINPUT51), .A4(new_n798), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n807), .A2(new_n391), .A3(new_n808), .A4(new_n811), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n540), .A2(new_n581), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n799), .A2(new_n813), .ZN(new_n814));
  XOR2_X1   g628(.A(new_n814), .B(KEYINPUT48), .Z(new_n815));
  AND2_X1   g629(.A1(new_n797), .A2(new_n604), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n812), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n713), .A2(new_n784), .A3(new_n714), .ZN(new_n818));
  INV_X1    g632(.A(new_n613), .ZN(new_n819));
  AND4_X1   g633(.A1(new_n819), .A2(new_n540), .A3(new_n612), .A4(new_n644), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n630), .B(new_n722), .C1(new_n818), .C2(new_n820), .ZN(new_n821));
  AND4_X1   g635(.A1(new_n733), .A2(new_n821), .A3(new_n742), .A4(new_n726), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n688), .B(new_n691), .C1(new_n698), .C2(new_n702), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT113), .ZN(new_n824));
  OAI22_X1  g638(.A1(new_n604), .A2(new_n824), .B1(new_n661), .B2(new_n819), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n744), .A2(KEYINPUT113), .A3(new_n613), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n273), .A2(new_n615), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n827), .A2(new_n581), .A3(new_n590), .A4(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n830), .A2(new_n582), .A3(new_n627), .A4(new_n693), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n823), .A2(new_n831), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n540), .A2(new_n273), .A3(new_n630), .ZN(new_n833));
  AOI22_X1  g647(.A1(new_n712), .A2(new_n715), .B1(new_n833), .B2(new_n739), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT52), .ZN(new_n835));
  INV_X1    g649(.A(new_n699), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n674), .B1(new_n836), .B2(new_n700), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n658), .A2(new_n464), .A3(new_n644), .A4(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n834), .A2(new_n681), .A3(new_n835), .A4(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n834), .A2(new_n681), .A3(new_n838), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(KEYINPUT52), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n822), .A2(new_n832), .A3(new_n839), .A4(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT53), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n841), .A2(new_n839), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(KEYINPUT114), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n734), .A2(new_n832), .A3(new_n742), .A4(new_n821), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT114), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n841), .A2(new_n849), .A3(new_n839), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n846), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n844), .B1(new_n851), .B2(new_n843), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(KEYINPUT54), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n851), .A2(new_n843), .ZN(new_n854));
  XOR2_X1   g668(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT115), .B1(new_n842), .B2(new_n843), .ZN(new_n857));
  INV_X1    g671(.A(new_n845), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT115), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n858), .A2(new_n848), .A3(new_n859), .A4(KEYINPUT53), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n854), .A2(new_n856), .A3(new_n857), .A4(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n817), .A2(new_n853), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(KEYINPUT117), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT117), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n817), .A2(new_n853), .A3(new_n861), .A4(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n390), .A2(new_n249), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(KEYINPUT118), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n779), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(KEYINPUT119), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT119), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n872), .B(new_n779), .C1(new_n866), .C2(new_n869), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n871), .A2(new_n873), .ZN(G75));
  NOR2_X1   g688(.A1(new_n845), .A2(new_n847), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n859), .B1(new_n875), .B2(KEYINPUT53), .ZN(new_n876));
  NOR4_X1   g690(.A1(new_n845), .A2(new_n847), .A3(KEYINPUT115), .A4(new_n843), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n266), .B1(new_n878), .B2(new_n854), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(G210), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT56), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n227), .A2(new_n258), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(new_n256), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT55), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n880), .A2(new_n881), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n884), .B1(new_n880), .B2(new_n881), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n390), .A2(G953), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n887), .B(KEYINPUT120), .Z(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n885), .A2(new_n886), .A3(new_n889), .ZN(G51));
  INV_X1    g704(.A(KEYINPUT121), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n758), .A2(KEYINPUT57), .ZN(new_n892));
  INV_X1    g706(.A(new_n850), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n849), .B1(new_n841), .B2(new_n839), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(KEYINPUT53), .B1(new_n895), .B2(new_n848), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n857), .A2(new_n860), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n855), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n892), .B1(new_n898), .B2(new_n861), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n758), .A2(KEYINPUT57), .ZN(new_n900));
  AOI211_X1 g714(.A(new_n891), .B(new_n683), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(new_n892), .ZN(new_n902));
  INV_X1    g716(.A(new_n861), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n856), .B1(new_n878), .B2(new_n854), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n900), .B(new_n902), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n683), .ZN(new_n906));
  AOI21_X1  g720(.A(KEYINPUT121), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n901), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n879), .A2(G469), .A3(new_n756), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n889), .B1(new_n908), .B2(new_n909), .ZN(G54));
  NAND3_X1  g724(.A1(new_n879), .A2(KEYINPUT58), .A3(G475), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n341), .A2(new_n342), .ZN(new_n912));
  OR2_X1    g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n911), .A2(new_n912), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n889), .B1(new_n913), .B2(new_n914), .ZN(G60));
  NAND2_X1  g729(.A1(new_n594), .A2(new_n596), .ZN(new_n916));
  XNOR2_X1  g730(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n388), .A2(new_n266), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n917), .B(new_n918), .Z(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  AOI211_X1 g734(.A(new_n916), .B(new_n920), .C1(new_n898), .C2(new_n861), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n853), .A2(new_n861), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(new_n919), .ZN(new_n923));
  AOI211_X1 g737(.A(new_n889), .B(new_n921), .C1(new_n916), .C2(new_n923), .ZN(G63));
  NAND2_X1  g738(.A1(new_n878), .A2(new_n854), .ZN(new_n925));
  NAND2_X1  g739(.A1(G217), .A2(G902), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT60), .Z(new_n927));
  AOI21_X1  g741(.A(new_n574), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n925), .A2(new_n624), .A3(new_n927), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n888), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT61), .ZN(new_n931));
  OAI22_X1  g745(.A1(new_n928), .A2(new_n930), .B1(KEYINPUT123), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(KEYINPUT123), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n932), .B(new_n933), .ZN(G66));
  INV_X1    g748(.A(new_n248), .ZN(new_n935));
  OAI21_X1  g749(.A(G953), .B1(new_n935), .B2(new_n395), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n936), .B1(new_n832), .B2(G953), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n882), .B1(G898), .B2(new_n249), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n937), .B(new_n938), .ZN(G69));
  INV_X1    g753(.A(new_n766), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n765), .B1(new_n750), .B2(new_n751), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n940), .A2(new_n941), .A3(new_n753), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n765), .A2(new_n813), .A3(new_n837), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n834), .A2(new_n681), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n773), .A2(new_n734), .A3(new_n742), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n942), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n249), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n516), .A2(new_n517), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(new_n330), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n948), .B(new_n950), .C1(new_n640), .C2(new_n249), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n737), .A2(new_n649), .ZN(new_n952));
  INV_X1    g766(.A(new_n827), .ZN(new_n953));
  OR3_X1    g767(.A1(new_n952), .A2(KEYINPUT124), .A3(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(KEYINPUT124), .B1(new_n952), .B2(new_n953), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(KEYINPUT125), .B1(new_n942), .B2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT125), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n767), .A2(new_n958), .A3(new_n955), .A4(new_n954), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n665), .A2(new_n944), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT62), .Z(new_n962));
  AND2_X1   g776(.A1(new_n962), .A2(new_n773), .ZN(new_n963));
  AOI21_X1  g777(.A(G953), .B1(new_n960), .B2(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n951), .B1(new_n964), .B2(new_n950), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(KEYINPUT126), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n249), .B1(G227), .B2(G900), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT126), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n951), .B(new_n968), .C1(new_n964), .C2(new_n950), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n966), .A2(new_n967), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n967), .B1(new_n966), .B2(new_n969), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n970), .A2(new_n971), .ZN(G72));
  INV_X1    g786(.A(new_n520), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n947), .A2(new_n832), .ZN(new_n974));
  NAND2_X1  g788(.A1(G472), .A2(G902), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT63), .Z(new_n976));
  AOI21_X1  g790(.A(new_n973), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n960), .A2(new_n963), .A3(new_n832), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n979), .A2(new_n976), .ZN(new_n980));
  OAI211_X1 g794(.A(new_n888), .B(new_n978), .C1(new_n980), .C2(new_n653), .ZN(new_n981));
  AND4_X1   g795(.A1(new_n973), .A2(new_n852), .A3(new_n653), .A4(new_n976), .ZN(new_n982));
  OAI21_X1  g796(.A(KEYINPUT127), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n653), .B1(new_n979), .B2(new_n976), .ZN(new_n984));
  NOR4_X1   g798(.A1(new_n984), .A2(new_n889), .A3(new_n977), .A4(new_n982), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT127), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n983), .A2(new_n987), .ZN(G57));
endmodule


