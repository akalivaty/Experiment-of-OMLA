//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 1 0 1 0 0 1 0 1 0 1 0 0 1 0 1 0 0 1 1 1 0 1 0 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:52 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n560, new_n562, new_n563, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n596, new_n597, new_n600, new_n602, new_n603, new_n604, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1113, new_n1114, new_n1115, new_n1117, new_n1118, new_n1119;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  AND3_X1   g037(.A1(new_n462), .A2(KEYINPUT67), .A3(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(KEYINPUT67), .B1(new_n462), .B2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n466), .B1(new_n462), .B2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n468), .A2(KEYINPUT66), .A3(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n471), .A2(G137), .B1(G101), .B2(G2104), .ZN(new_n472));
  OR2_X1    g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n462), .A2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n475));
  OR2_X1    g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  AOI22_X1  g052(.A1(new_n477), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n478));
  INV_X1    g053(.A(G2105), .ZN(new_n479));
  OR2_X1    g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n473), .A2(new_n480), .ZN(G160));
  NAND2_X1  g056(.A1(new_n465), .A2(new_n470), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(new_n479), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n482), .A2(G2105), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n479), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n484), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  NAND4_X1  g065(.A1(new_n465), .A2(G138), .A3(new_n479), .A4(new_n470), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT69), .ZN(new_n493));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  NOR4_X1   g069(.A1(new_n476), .A2(KEYINPUT4), .A3(new_n494), .A4(G2105), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT69), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n491), .A2(new_n497), .A3(KEYINPUT4), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n493), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n471), .A2(G126), .A3(G2105), .ZN(new_n500));
  OR2_X1    g075(.A1(new_n479), .A2(G114), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT68), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n468), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI221_X1 g078(.A(new_n503), .B1(new_n502), .B2(new_n501), .C1(G102), .C2(G2105), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n499), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n499), .A2(new_n506), .A3(KEYINPUT70), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(G164));
  NAND2_X1  g086(.A1(G50), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT71), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  OR3_X1    g089(.A1(new_n513), .A2(new_n514), .A3(KEYINPUT5), .ZN(new_n515));
  OAI21_X1  g090(.A(KEYINPUT5), .B1(new_n513), .B2(new_n514), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n512), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT6), .B(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  XOR2_X1   g096(.A(new_n521), .B(KEYINPUT72), .Z(new_n522));
  NAND2_X1  g097(.A1(G75), .A2(G543), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT73), .ZN(new_n524));
  INV_X1    g099(.A(G62), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n524), .B1(new_n517), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n522), .A2(new_n527), .ZN(G303));
  INV_X1    g103(.A(G303), .ZN(G166));
  XOR2_X1   g104(.A(KEYINPUT6), .B(G651), .Z(new_n530));
  INV_X1    g105(.A(KEYINPUT74), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n520), .A2(KEYINPUT74), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n532), .A2(G543), .A3(new_n533), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT75), .ZN(new_n535));
  XNOR2_X1  g110(.A(KEYINPUT76), .B(G51), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n520), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n538), .A2(new_n517), .ZN(new_n539));
  XOR2_X1   g114(.A(KEYINPUT77), .B(KEYINPUT7), .Z(new_n540));
  NAND3_X1  g115(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n540), .B(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n537), .A2(new_n539), .A3(new_n542), .ZN(G286));
  INV_X1    g118(.A(G286), .ZN(G168));
  NAND2_X1  g119(.A1(new_n535), .A2(G52), .ZN(new_n545));
  NAND2_X1  g120(.A1(G77), .A2(G543), .ZN(new_n546));
  INV_X1    g121(.A(G64), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n517), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n517), .A2(new_n530), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n548), .A2(G651), .B1(new_n549), .B2(G90), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n545), .A2(new_n550), .ZN(G301));
  INV_X1    g126(.A(G301), .ZN(G171));
  NAND2_X1  g127(.A1(new_n535), .A2(G43), .ZN(new_n553));
  NAND2_X1  g128(.A1(G68), .A2(G543), .ZN(new_n554));
  INV_X1    g129(.A(G56), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n517), .B2(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n556), .A2(G651), .B1(new_n549), .B2(G81), .ZN(new_n557));
  AND2_X1   g132(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  AND3_X1   g134(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G36), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n560), .A2(new_n563), .ZN(G188));
  AND3_X1   g139(.A1(new_n532), .A2(G543), .A3(new_n533), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n565), .A2(KEYINPUT78), .A3(G53), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT9), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n549), .A2(G91), .ZN(new_n568));
  INV_X1    g143(.A(G651), .ZN(new_n569));
  INV_X1    g144(.A(new_n517), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n570), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n571));
  OAI211_X1 g146(.A(new_n567), .B(new_n568), .C1(new_n569), .C2(new_n571), .ZN(G299));
  NAND2_X1  g147(.A1(new_n565), .A2(G49), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT79), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n573), .B(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n549), .A2(G87), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n570), .B2(G74), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(G288));
  AOI22_X1  g153(.A1(new_n570), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n570), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n580));
  OAI22_X1  g155(.A1(new_n569), .A2(new_n579), .B1(new_n580), .B2(new_n530), .ZN(G305));
  NAND2_X1  g156(.A1(new_n535), .A2(G47), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n549), .A2(G85), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n570), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  OAI211_X1 g159(.A(new_n582), .B(new_n583), .C1(new_n569), .C2(new_n584), .ZN(G290));
  NAND2_X1  g160(.A1(G301), .A2(G868), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n549), .A2(G92), .ZN(new_n587));
  XOR2_X1   g162(.A(new_n587), .B(KEYINPUT10), .Z(new_n588));
  NAND2_X1  g163(.A1(new_n535), .A2(G54), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n570), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n590));
  OR2_X1    g165(.A1(new_n590), .A2(new_n569), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n588), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n586), .B1(new_n593), .B2(G868), .ZN(G284));
  XNOR2_X1  g169(.A(G284), .B(KEYINPUT80), .ZN(G321));
  INV_X1    g170(.A(G868), .ZN(new_n596));
  NAND2_X1  g171(.A1(G299), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(new_n596), .B2(G168), .ZN(G297));
  OAI21_X1  g173(.A(new_n597), .B1(new_n596), .B2(G168), .ZN(G280));
  INV_X1    g174(.A(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n593), .B1(new_n600), .B2(G860), .ZN(G148));
  INV_X1    g176(.A(new_n558), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(new_n596), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n592), .A2(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(new_n596), .ZN(G323));
  XNOR2_X1  g180(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g181(.A1(new_n485), .A2(G135), .ZN(new_n607));
  OR2_X1    g182(.A1(new_n607), .A2(KEYINPUT81), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n607), .A2(KEYINPUT81), .B1(G123), .B2(new_n483), .ZN(new_n609));
  OR2_X1    g184(.A1(new_n479), .A2(G111), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n468), .B1(new_n610), .B2(KEYINPUT82), .ZN(new_n611));
  OAI221_X1 g186(.A(new_n611), .B1(KEYINPUT82), .B2(new_n610), .C1(G99), .C2(G2105), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n608), .A2(new_n609), .A3(new_n612), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(G2096), .Z(new_n614));
  NAND3_X1  g189(.A1(new_n479), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(KEYINPUT12), .Z(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT13), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(G2100), .Z(new_n618));
  NAND2_X1  g193(.A1(new_n614), .A2(new_n618), .ZN(G156));
  XNOR2_X1  g194(.A(G2451), .B(G2454), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT16), .ZN(new_n621));
  XOR2_X1   g196(.A(G2443), .B(G2446), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(G1341), .B(G1348), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT15), .B(G2435), .ZN(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT83), .B(G2438), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(G2427), .B(G2430), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(KEYINPUT14), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n625), .B(new_n631), .ZN(new_n632));
  AND2_X1   g207(.A1(new_n632), .A2(G14), .ZN(G401));
  XOR2_X1   g208(.A(G2072), .B(G2078), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT84), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n635), .A2(KEYINPUT17), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(KEYINPUT17), .ZN(new_n637));
  XOR2_X1   g212(.A(G2067), .B(G2678), .Z(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G2084), .B(G2090), .Z(new_n640));
  NOR2_X1   g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n639), .A2(new_n640), .ZN(new_n643));
  NAND4_X1  g218(.A1(new_n636), .A2(new_n637), .A3(new_n642), .A4(new_n643), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n643), .A2(new_n634), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT18), .ZN(new_n646));
  OAI211_X1 g221(.A(new_n644), .B(new_n646), .C1(new_n634), .C2(new_n642), .ZN(new_n647));
  XOR2_X1   g222(.A(G2096), .B(G2100), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT85), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n647), .B(new_n649), .ZN(G227));
  INV_X1    g225(.A(KEYINPUT20), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1956), .B(G2474), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT86), .ZN(new_n653));
  XOR2_X1   g228(.A(G1961), .B(G1966), .Z(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1971), .B(G1976), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT19), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n651), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n653), .A2(new_n654), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n660), .A2(new_n657), .A3(new_n655), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n655), .A2(new_n651), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n662), .A2(new_n659), .ZN(new_n663));
  OAI211_X1 g238(.A(new_n658), .B(new_n661), .C1(new_n663), .C2(new_n657), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G1991), .ZN(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G1981), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1986), .B(G1996), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n665), .B(new_n669), .ZN(G229));
  INV_X1    g245(.A(G29), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(G25), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n485), .A2(G131), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT87), .Z(new_n674));
  OR2_X1    g249(.A1(G95), .A2(G2105), .ZN(new_n675));
  OAI211_X1 g250(.A(new_n675), .B(G2104), .C1(G107), .C2(new_n479), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n483), .A2(G119), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n674), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n672), .B1(new_n679), .B2(new_n671), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT35), .B(G1991), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT88), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n680), .B(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(G1986), .ZN(new_n685));
  INV_X1    g260(.A(G16), .ZN(new_n686));
  AND2_X1   g261(.A1(new_n686), .A2(G24), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(G290), .B2(G16), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n684), .B1(new_n685), .B2(new_n688), .ZN(new_n689));
  AND2_X1   g264(.A1(new_n686), .A2(G22), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n690), .B1(G303), .B2(G16), .ZN(new_n691));
  INV_X1    g266(.A(G1971), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n686), .A2(G23), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(G288), .B2(G16), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT33), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n693), .B1(new_n696), .B2(G1976), .ZN(new_n697));
  MUX2_X1   g272(.A(G6), .B(G305), .S(G16), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT89), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT32), .B(G1981), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n697), .B(new_n701), .C1(G1976), .C2(new_n696), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n689), .B1(new_n702), .B2(KEYINPUT34), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n688), .A2(new_n685), .ZN(new_n704));
  OAI211_X1 g279(.A(new_n703), .B(new_n704), .C1(KEYINPUT34), .C2(new_n702), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT90), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n705), .A2(new_n706), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n707), .A2(KEYINPUT36), .A3(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT91), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n709), .B(new_n710), .C1(KEYINPUT36), .C2(new_n705), .ZN(new_n711));
  NAND2_X1  g286(.A1(G299), .A2(G16), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(KEYINPUT23), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n686), .A2(G20), .ZN(new_n714));
  MUX2_X1   g289(.A(KEYINPUT23), .B(new_n713), .S(new_n714), .Z(new_n715));
  INV_X1    g290(.A(G1956), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NAND4_X1  g292(.A1(new_n707), .A2(KEYINPUT91), .A3(KEYINPUT36), .A4(new_n708), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n671), .A2(G35), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G162), .B2(new_n671), .ZN(new_n720));
  MUX2_X1   g295(.A(new_n719), .B(new_n720), .S(KEYINPUT98), .Z(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT99), .B(KEYINPUT29), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n721), .B(new_n722), .Z(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G2090), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT100), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G2090), .B2(new_n723), .ZN(new_n726));
  NOR2_X1   g301(.A1(G29), .A2(G33), .ZN(new_n727));
  AOI22_X1  g302(.A1(new_n477), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n728), .A2(new_n479), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n485), .A2(G139), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n479), .A2(G103), .A3(G2104), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT25), .Z(new_n732));
  NAND3_X1  g307(.A1(new_n729), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT93), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n727), .B1(new_n734), .B2(G29), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(G2072), .Z(new_n736));
  OR2_X1    g311(.A1(KEYINPUT24), .A2(G34), .ZN(new_n737));
  NAND2_X1  g312(.A1(KEYINPUT24), .A2(G34), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n737), .A2(new_n671), .A3(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G160), .B2(new_n671), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(G2084), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT27), .B(G1996), .Z(new_n742));
  NAND2_X1  g317(.A1(new_n671), .A2(G32), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n485), .A2(G141), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n483), .A2(G129), .ZN(new_n745));
  NAND3_X1  g320(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT26), .Z(new_n747));
  NAND3_X1  g322(.A1(new_n479), .A2(G105), .A3(G2104), .ZN(new_n748));
  NAND4_X1  g323(.A1(new_n744), .A2(new_n745), .A3(new_n747), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT94), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n743), .B1(new_n750), .B2(new_n671), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n736), .B(new_n741), .C1(new_n742), .C2(new_n751), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT95), .ZN(new_n753));
  NOR2_X1   g328(.A1(G168), .A2(new_n686), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(new_n686), .B2(G21), .ZN(new_n755));
  INV_X1    g330(.A(G1966), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n558), .A2(new_n686), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n686), .B2(G19), .ZN(new_n758));
  INV_X1    g333(.A(G1341), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n755), .A2(new_n756), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(G5), .A2(G16), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G171), .B2(G16), .ZN(new_n762));
  INV_X1    g337(.A(G1961), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  OAI211_X1 g339(.A(new_n760), .B(new_n764), .C1(new_n759), .C2(new_n758), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n740), .A2(G2084), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT31), .B(G11), .ZN(new_n767));
  INV_X1    g342(.A(G28), .ZN(new_n768));
  AOI21_X1  g343(.A(G29), .B1(new_n768), .B2(KEYINPUT30), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n769), .A2(KEYINPUT96), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n769), .A2(KEYINPUT96), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n770), .B(new_n771), .C1(KEYINPUT30), .C2(new_n768), .ZN(new_n772));
  OAI211_X1 g347(.A(new_n767), .B(new_n772), .C1(new_n613), .C2(new_n671), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT97), .Z(new_n774));
  NAND2_X1  g349(.A1(new_n751), .A2(new_n742), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n774), .B(new_n775), .C1(new_n756), .C2(new_n755), .ZN(new_n776));
  NOR3_X1   g351(.A1(new_n765), .A2(new_n766), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n686), .A2(G4), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n593), .B2(new_n686), .ZN(new_n779));
  INV_X1    g354(.A(G1348), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n483), .A2(G128), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n485), .A2(G140), .ZN(new_n783));
  OR2_X1    g358(.A1(G104), .A2(G2105), .ZN(new_n784));
  OAI211_X1 g359(.A(new_n784), .B(G2104), .C1(G116), .C2(new_n479), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n782), .A2(new_n783), .A3(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT92), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n788), .A2(new_n671), .ZN(new_n789));
  AND2_X1   g364(.A1(new_n671), .A2(G26), .ZN(new_n790));
  OAI21_X1  g365(.A(KEYINPUT28), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(KEYINPUT28), .B2(new_n790), .ZN(new_n792));
  INV_X1    g367(.A(G2067), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n777), .A2(new_n781), .A3(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(G27), .A2(G29), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G164), .B2(G29), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G2078), .ZN(new_n798));
  NOR4_X1   g373(.A1(new_n726), .A2(new_n753), .A3(new_n795), .A4(new_n798), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n711), .A2(new_n717), .A3(new_n718), .A4(new_n799), .ZN(G150));
  INV_X1    g375(.A(G150), .ZN(G311));
  NOR2_X1   g376(.A1(new_n592), .A2(new_n600), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT39), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n535), .A2(G55), .ZN(new_n806));
  NAND2_X1  g381(.A1(G80), .A2(G543), .ZN(new_n807));
  INV_X1    g382(.A(G67), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n807), .B1(new_n517), .B2(new_n808), .ZN(new_n809));
  AOI22_X1  g384(.A1(new_n809), .A2(G651), .B1(new_n549), .B2(G93), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n806), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n558), .B(new_n811), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n805), .B(new_n812), .Z(new_n813));
  NOR2_X1   g388(.A1(new_n813), .A2(G860), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT102), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n811), .A2(G860), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT37), .Z(new_n817));
  NAND2_X1  g392(.A1(new_n815), .A2(new_n817), .ZN(G145));
  NAND2_X1  g393(.A1(new_n473), .A2(new_n480), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(new_n489), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n678), .B(new_n616), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n483), .A2(G130), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n485), .A2(G142), .ZN(new_n823));
  OR2_X1    g398(.A1(G106), .A2(G2105), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n824), .B(G2104), .C1(G118), .C2(new_n479), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n822), .A2(new_n823), .A3(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(new_n507), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n788), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n786), .B(KEYINPUT92), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(new_n507), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n828), .A2(new_n830), .A3(new_n750), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n750), .B1(new_n828), .B2(new_n830), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT103), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n834), .A2(new_n835), .A3(new_n734), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n828), .A2(new_n830), .ZN(new_n837));
  INV_X1    g412(.A(new_n750), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n839), .A2(new_n734), .A3(new_n831), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(KEYINPUT103), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n836), .A2(new_n841), .ZN(new_n842));
  AND3_X1   g417(.A1(new_n828), .A2(new_n830), .A3(new_n749), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n749), .B1(new_n828), .B2(new_n830), .ZN(new_n844));
  INV_X1    g419(.A(new_n733), .ZN(new_n845));
  NOR3_X1   g420(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n826), .B1(new_n842), .B2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n826), .ZN(new_n849));
  AOI211_X1 g424(.A(new_n849), .B(new_n846), .C1(new_n836), .C2(new_n841), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n821), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n835), .B1(new_n834), .B2(new_n734), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n840), .A2(KEYINPUT103), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n847), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(new_n849), .ZN(new_n855));
  INV_X1    g430(.A(new_n821), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n842), .A2(new_n826), .A3(new_n847), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n613), .ZN(new_n859));
  AND3_X1   g434(.A1(new_n851), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n859), .B1(new_n851), .B2(new_n858), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n820), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NOR3_X1   g437(.A1(new_n848), .A2(new_n850), .A3(new_n821), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n856), .B1(new_n855), .B2(new_n857), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n613), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n820), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n851), .A2(new_n858), .A3(new_n859), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(G37), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n862), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g446(.A1(new_n811), .A2(G868), .ZN(new_n872));
  XNOR2_X1  g447(.A(G290), .B(G305), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(G303), .ZN(new_n874));
  INV_X1    g449(.A(G288), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n874), .B(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT104), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n877), .B1(new_n878), .B2(KEYINPUT42), .ZN(new_n879));
  XNOR2_X1  g454(.A(KEYINPUT104), .B(KEYINPUT42), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n879), .B1(new_n877), .B2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT105), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n812), .B(new_n604), .Z(new_n883));
  XNOR2_X1  g458(.A(G299), .B(new_n592), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n884), .A2(KEYINPUT41), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(KEYINPUT41), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n883), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n884), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n887), .B1(new_n888), .B2(new_n883), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n881), .B1(new_n882), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n882), .ZN(new_n891));
  XOR2_X1   g466(.A(new_n890), .B(new_n891), .Z(new_n892));
  AOI21_X1  g467(.A(new_n872), .B1(new_n892), .B2(G868), .ZN(G295));
  AOI21_X1  g468(.A(new_n872), .B1(new_n892), .B2(G868), .ZN(G331));
  INV_X1    g469(.A(KEYINPUT43), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n812), .B(G301), .ZN(new_n896));
  OR2_X1    g471(.A1(new_n896), .A2(G168), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(G168), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n885), .A2(new_n886), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n897), .A2(new_n888), .A3(new_n898), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n901), .A2(new_n877), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(new_n869), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT106), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n885), .B(new_n905), .ZN(new_n906));
  XOR2_X1   g481(.A(new_n886), .B(KEYINPUT107), .Z(new_n907));
  OAI21_X1  g482(.A(new_n899), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(new_n902), .ZN(new_n909));
  AOI211_X1 g484(.A(new_n895), .B(new_n904), .C1(new_n876), .C2(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n877), .B1(new_n901), .B2(new_n902), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n904), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n912), .A2(KEYINPUT43), .ZN(new_n913));
  OAI21_X1  g488(.A(KEYINPUT44), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n909), .A2(new_n876), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n915), .A2(new_n895), .A3(new_n869), .A4(new_n903), .ZN(new_n916));
  OAI21_X1  g491(.A(KEYINPUT43), .B1(new_n904), .B2(new_n911), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n914), .B1(KEYINPUT44), .B2(new_n918), .ZN(G397));
  XNOR2_X1  g494(.A(KEYINPUT108), .B(G40), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(G160), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(G1384), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n491), .A2(new_n497), .A3(KEYINPUT4), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n497), .B1(new_n491), .B2(KEYINPUT4), .ZN(new_n925));
  NOR3_X1   g500(.A1(new_n924), .A2(new_n925), .A3(new_n495), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n923), .B1(new_n926), .B2(new_n505), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  NOR3_X1   g503(.A1(new_n922), .A2(new_n928), .A3(KEYINPUT45), .ZN(new_n929));
  INV_X1    g504(.A(G1996), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT125), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(KEYINPUT46), .ZN(new_n933));
  XOR2_X1   g508(.A(new_n931), .B(new_n933), .Z(new_n934));
  NAND2_X1  g509(.A1(new_n829), .A2(G2067), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n788), .A2(new_n793), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n929), .B1(new_n938), .B2(new_n749), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n934), .B(new_n939), .C1(new_n932), .C2(KEYINPUT46), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n940), .B(KEYINPUT47), .ZN(new_n941));
  INV_X1    g516(.A(new_n929), .ZN(new_n942));
  NOR3_X1   g517(.A1(new_n942), .A2(G1986), .A3(G290), .ZN(new_n943));
  XOR2_X1   g518(.A(new_n943), .B(KEYINPUT48), .Z(new_n944));
  NAND2_X1  g519(.A1(new_n749), .A2(G1996), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n937), .B(new_n945), .C1(G1996), .C2(new_n838), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n678), .B(new_n682), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n944), .B1(new_n942), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n679), .A2(new_n683), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n936), .B1(new_n946), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n929), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n941), .A2(new_n949), .A3(new_n952), .ZN(new_n953));
  XOR2_X1   g528(.A(new_n953), .B(KEYINPUT126), .Z(new_n954));
  NOR2_X1   g529(.A1(new_n819), .A2(new_n920), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT109), .B1(new_n507), .B2(new_n923), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT109), .ZN(new_n957));
  AOI211_X1 g532(.A(new_n957), .B(G1384), .C1(new_n499), .C2(new_n506), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n955), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(G8), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n960), .B(KEYINPUT110), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n875), .A2(G1976), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(KEYINPUT111), .A2(KEYINPUT52), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OR3_X1    g540(.A1(new_n875), .A2(KEYINPUT52), .A3(G1976), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n961), .A2(KEYINPUT111), .A3(KEYINPUT52), .A4(new_n962), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  XOR2_X1   g543(.A(G305), .B(G1981), .Z(new_n969));
  NOR2_X1   g544(.A1(KEYINPUT112), .A2(KEYINPUT49), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n969), .B(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n961), .A2(new_n971), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n968), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n509), .A2(new_n923), .A3(new_n510), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT45), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n928), .A2(KEYINPUT45), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n976), .A2(new_n955), .A3(new_n977), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n978), .A2(G1971), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n922), .B1(new_n974), .B2(KEYINPUT50), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT50), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n981), .B1(new_n956), .B2(new_n958), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n983), .A2(G2090), .ZN(new_n984));
  OAI21_X1  g559(.A(G8), .B1(new_n979), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(G303), .A2(G8), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n986), .B(KEYINPUT55), .ZN(new_n987));
  OR2_X1    g562(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n927), .A2(new_n957), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n507), .A2(KEYINPUT109), .A3(new_n923), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n989), .A2(new_n975), .A3(new_n990), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n991), .B(new_n955), .C1(new_n975), .C2(new_n974), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n756), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT115), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n992), .A2(KEYINPUT115), .A3(new_n756), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(KEYINPUT116), .B1(new_n983), .B2(G2084), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT116), .ZN(new_n999));
  INV_X1    g574(.A(G2084), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n980), .A2(new_n999), .A3(new_n1000), .A4(new_n982), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n998), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n997), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1003), .A2(G8), .A3(G168), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT63), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1006), .B1(new_n985), .B2(new_n987), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n973), .A2(new_n988), .A3(new_n1005), .A4(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n968), .A2(new_n988), .A3(new_n972), .ZN(new_n1009));
  INV_X1    g584(.A(new_n987), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n989), .A2(KEYINPUT50), .A3(new_n990), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n955), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT114), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n974), .A2(KEYINPUT50), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1011), .A2(KEYINPUT114), .A3(new_n955), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1014), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  OAI22_X1  g593(.A1(new_n1018), .A2(G2090), .B1(G1971), .B2(new_n978), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1010), .B1(new_n1019), .B2(G8), .ZN(new_n1020));
  NOR3_X1   g595(.A1(new_n1009), .A2(new_n1020), .A3(new_n1004), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1008), .B1(new_n1021), .B2(KEYINPUT63), .ZN(new_n1022));
  INV_X1    g597(.A(new_n988), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n973), .A2(new_n1023), .ZN(new_n1024));
  XOR2_X1   g599(.A(new_n961), .B(KEYINPUT113), .Z(new_n1025));
  AOI211_X1 g600(.A(G1976), .B(G288), .C1(new_n961), .C2(new_n971), .ZN(new_n1026));
  NOR2_X1   g601(.A1(G305), .A2(G1981), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1025), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1022), .A2(new_n1024), .A3(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n997), .A2(G168), .A3(new_n1002), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT123), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1030), .A2(new_n1031), .A3(G8), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(KEYINPUT51), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1003), .A2(G8), .A3(G286), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT51), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1030), .A2(new_n1031), .A3(new_n1035), .A4(G8), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1033), .A2(new_n1034), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(KEYINPUT62), .ZN(new_n1038));
  OR2_X1    g613(.A1(new_n992), .A2(G2078), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT124), .ZN(new_n1040));
  OR2_X1    g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1041), .A2(KEYINPUT53), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G2078), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT53), .B1(new_n978), .B2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1045), .B1(new_n763), .B2(new_n983), .ZN(new_n1046));
  AND2_X1   g621(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1047), .A2(G301), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT62), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1033), .A2(new_n1049), .A3(new_n1034), .A4(new_n1036), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1038), .A2(new_n1048), .A3(new_n1050), .ZN(new_n1051));
  XOR2_X1   g626(.A(KEYINPUT58), .B(G1341), .Z(new_n1052));
  AOI22_X1  g627(.A1(new_n978), .A2(new_n930), .B1(new_n959), .B2(new_n1052), .ZN(new_n1053));
  OR2_X1    g628(.A1(new_n1053), .A2(new_n602), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT59), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1054), .A2(KEYINPUT121), .A3(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT61), .ZN(new_n1057));
  XNOR2_X1  g632(.A(KEYINPUT56), .B(G2072), .ZN(new_n1058));
  AND4_X1   g633(.A1(new_n955), .A2(new_n976), .A3(new_n977), .A4(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1059), .B1(new_n1018), .B2(new_n716), .ZN(new_n1060));
  XOR2_X1   g635(.A(G299), .B(KEYINPUT57), .Z(new_n1061));
  OAI21_X1  g636(.A(new_n1057), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  AND2_X1   g637(.A1(new_n1057), .A2(KEYINPUT122), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1063), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1056), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  AND2_X1   g640(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1066));
  XOR2_X1   g641(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n1067));
  NOR2_X1   g642(.A1(new_n1054), .A2(new_n1067), .ZN(new_n1068));
  NOR3_X1   g643(.A1(new_n1065), .A2(new_n1066), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n983), .A2(new_n780), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n922), .B1(new_n989), .B2(new_n990), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(new_n793), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1070), .A2(KEYINPUT117), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT117), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1072), .ZN(new_n1075));
  AOI21_X1  g650(.A(G1348), .B1(new_n980), .B2(new_n982), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1074), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT60), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1073), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(new_n593), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1078), .B1(new_n1073), .B2(new_n1077), .ZN(new_n1081));
  XOR2_X1   g656(.A(new_n1080), .B(new_n1081), .Z(new_n1082));
  INV_X1    g657(.A(new_n1059), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1011), .A2(KEYINPUT114), .A3(new_n955), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT114), .B1(new_n1011), .B2(new_n955), .ZN(new_n1085));
  NOR3_X1   g660(.A1(new_n1084), .A2(new_n1085), .A3(new_n1015), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1083), .B1(new_n1086), .B2(G1956), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT119), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1061), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1060), .A2(KEYINPUT119), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(KEYINPUT120), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT120), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1089), .A2(new_n1091), .A3(new_n1094), .A4(new_n1090), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1073), .A2(new_n1077), .A3(new_n593), .ZN(new_n1096));
  XNOR2_X1  g671(.A(new_n1096), .B(KEYINPUT118), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1093), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1099));
  AOI22_X1  g674(.A1(new_n1069), .A2(new_n1082), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  XOR2_X1   g675(.A(G301), .B(KEYINPUT54), .Z(new_n1101));
  AND4_X1   g676(.A1(KEYINPUT53), .A2(new_n977), .A3(G40), .A4(new_n1044), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1102), .B(G160), .C1(KEYINPUT45), .C2(new_n928), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1046), .A2(new_n1101), .A3(new_n1103), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1037), .B(new_n1104), .C1(new_n1101), .C2(new_n1047), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1051), .B1(new_n1100), .B2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1009), .A2(new_n1020), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1029), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(G290), .B(new_n685), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n942), .B1(new_n948), .B2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n954), .B1(new_n1108), .B2(new_n1110), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g686(.A1(G229), .A2(new_n460), .ZN(new_n1113));
  AOI21_X1  g687(.A(new_n1113), .B1(new_n916), .B2(new_n917), .ZN(new_n1114));
  NOR2_X1   g688(.A1(G401), .A2(G227), .ZN(new_n1115));
  NAND3_X1  g689(.A1(new_n870), .A2(new_n1114), .A3(new_n1115), .ZN(G225));
  NAND2_X1  g690(.A1(G225), .A2(KEYINPUT127), .ZN(new_n1117));
  INV_X1    g691(.A(KEYINPUT127), .ZN(new_n1118));
  NAND4_X1  g692(.A1(new_n870), .A2(new_n1114), .A3(new_n1118), .A4(new_n1115), .ZN(new_n1119));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1119), .ZN(G308));
endmodule


