//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 0 1 0 1 0 0 0 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 1 1 1 0 0 0 1 1 1 1 0 0 1 0 0 0 1 0 1 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n635, new_n636, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n821, new_n823, new_n824, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n870, new_n871, new_n872, new_n873, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n893, new_n894, new_n895, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n947, new_n948;
  XOR2_X1   g000(.A(G211gat), .B(G218gat), .Z(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT77), .ZN(new_n203));
  XNOR2_X1  g002(.A(G197gat), .B(G204gat), .ZN(new_n204));
  INV_X1    g003(.A(G211gat), .ZN(new_n205));
  INV_X1    g004(.A(G218gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n204), .B1(KEYINPUT22), .B2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n203), .B(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G226gat), .A2(G233gat), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  AND3_X1   g010(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT68), .ZN(new_n215));
  NAND2_X1  g014(.A1(G183gat), .A2(G190gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT66), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n216), .B(new_n217), .ZN(new_n218));
  XOR2_X1   g017(.A(KEYINPUT67), .B(KEYINPUT24), .Z(new_n219));
  AOI21_X1  g018(.A(new_n215), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n219), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n221), .A2(KEYINPUT68), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n214), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT25), .ZN(new_n224));
  NOR2_X1   g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n225), .B1(KEYINPUT23), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n225), .B(KEYINPUT65), .ZN(new_n228));
  AOI211_X1 g027(.A(new_n224), .B(new_n227), .C1(new_n228), .C2(KEYINPUT23), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n223), .A2(new_n229), .ZN(new_n230));
  OR2_X1    g029(.A1(new_n212), .A2(KEYINPUT64), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n212), .A2(KEYINPUT64), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT24), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n213), .B1(new_n233), .B2(new_n216), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n231), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n227), .B1(KEYINPUT23), .B2(new_n225), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(new_n224), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n230), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT27), .B(G183gat), .ZN(new_n240));
  INV_X1    g039(.A(G190gat), .ZN(new_n241));
  AND3_X1   g040(.A1(new_n240), .A2(KEYINPUT28), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n241), .ZN(new_n243));
  XNOR2_X1  g042(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT70), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n242), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n245), .A2(KEYINPUT70), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT26), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n228), .A2(new_n251), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n252), .B(new_n226), .C1(new_n251), .C2(new_n225), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n250), .A2(new_n216), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n239), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT29), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n211), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n210), .B1(new_n239), .B2(new_n254), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n209), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n258), .ZN(new_n260));
  INV_X1    g059(.A(new_n209), .ZN(new_n261));
  AOI21_X1  g060(.A(KEYINPUT29), .B1(new_n239), .B2(new_n254), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n260), .B(new_n261), .C1(new_n262), .C2(new_n211), .ZN(new_n263));
  XNOR2_X1  g062(.A(G8gat), .B(G36gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n264), .B(KEYINPUT78), .ZN(new_n265));
  XNOR2_X1  g064(.A(G64gat), .B(G92gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n259), .A2(new_n263), .A3(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT37), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n259), .A2(new_n263), .A3(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n267), .B(KEYINPUT79), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n271), .A2(KEYINPUT38), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n269), .B1(new_n259), .B2(new_n263), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n268), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(G225gat), .A2(G233gat), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(KEYINPUT71), .B(G120gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(G113gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(G127gat), .B(G134gat), .ZN(new_n281));
  INV_X1    g080(.A(G113gat), .ZN(new_n282));
  INV_X1    g081(.A(G120gat), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT1), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n280), .A2(new_n281), .A3(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT72), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n284), .B1(new_n282), .B2(new_n283), .ZN(new_n287));
  INV_X1    g086(.A(new_n281), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n285), .A2(new_n286), .A3(new_n289), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n280), .A2(KEYINPUT72), .A3(new_n281), .A4(new_n284), .ZN(new_n291));
  AND2_X1   g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  XOR2_X1   g091(.A(G141gat), .B(G148gat), .Z(new_n293));
  INV_X1    g092(.A(G155gat), .ZN(new_n294));
  INV_X1    g093(.A(G162gat), .ZN(new_n295));
  OAI21_X1  g094(.A(KEYINPUT2), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  XOR2_X1   g096(.A(G155gat), .B(G162gat), .Z(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n297), .B(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT3), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n297), .B(new_n298), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT3), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n292), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT80), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT80), .ZN(new_n307));
  NAND4_X1  g106(.A1(new_n292), .A2(new_n302), .A3(new_n304), .A4(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n278), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n290), .A2(new_n291), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(new_n300), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n311), .B(KEYINPUT4), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT82), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n292), .A2(new_n303), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n315), .A2(KEYINPUT81), .A3(new_n311), .ZN(new_n316));
  OR3_X1    g115(.A1(new_n310), .A2(new_n300), .A3(KEYINPUT81), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n314), .B1(new_n318), .B2(new_n277), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n316), .A2(KEYINPUT82), .A3(new_n278), .A4(new_n317), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n313), .A2(new_n319), .A3(KEYINPUT5), .A4(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT5), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT4), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n311), .B(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT83), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n312), .A2(KEYINPUT83), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n322), .B(new_n309), .C1(new_n326), .C2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n321), .A2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(G1gat), .B(G29gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n330), .B(KEYINPUT0), .ZN(new_n331));
  XNOR2_X1  g130(.A(G57gat), .B(G85gat), .ZN(new_n332));
  XOR2_X1   g131(.A(new_n331), .B(new_n332), .Z(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n329), .A2(KEYINPUT6), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n329), .A2(new_n334), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT6), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n321), .A2(new_n328), .A3(new_n333), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n267), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n270), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT38), .B1(new_n341), .B2(new_n274), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n276), .A2(new_n335), .A3(new_n339), .A4(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n301), .B1(new_n209), .B2(KEYINPUT29), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(new_n303), .ZN(new_n345));
  INV_X1    g144(.A(G228gat), .ZN(new_n346));
  INV_X1    g145(.A(G233gat), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n261), .B1(new_n302), .B2(new_n256), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT85), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n345), .B(new_n348), .C1(new_n349), .C2(new_n350), .ZN(new_n351));
  AND2_X1   g150(.A1(new_n349), .A2(new_n350), .ZN(new_n352));
  OR2_X1    g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n202), .ZN(new_n354));
  AOI21_X1  g153(.A(KEYINPUT29), .B1(new_n208), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n355), .B1(new_n354), .B2(new_n208), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n300), .B1(new_n356), .B2(new_n301), .ZN(new_n357));
  OAI22_X1  g156(.A1(new_n349), .A2(new_n357), .B1(new_n346), .B2(new_n347), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n353), .A2(KEYINPUT86), .A3(new_n358), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n358), .B1(new_n351), .B2(new_n352), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT86), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(G22gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(KEYINPUT84), .B(KEYINPUT31), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n364), .B(G50gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(G78gat), .B(G106gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n365), .B(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n362), .A2(new_n363), .A3(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n363), .B1(new_n362), .B2(new_n367), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n359), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n370), .ZN(new_n372));
  INV_X1    g171(.A(new_n359), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n372), .A2(new_n373), .A3(new_n368), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n324), .A2(new_n325), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n312), .A2(KEYINPUT83), .ZN(new_n378));
  AOI22_X1  g177(.A1(new_n377), .A2(new_n378), .B1(new_n306), .B2(new_n308), .ZN(new_n379));
  OAI21_X1  g178(.A(KEYINPUT87), .B1(new_n379), .B2(new_n277), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n306), .A2(new_n308), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n381), .B1(new_n326), .B2(new_n327), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT87), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n382), .A2(new_n383), .A3(new_n278), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n380), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT39), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n334), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n386), .B1(new_n318), .B2(new_n277), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n380), .A2(new_n384), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n387), .A2(KEYINPUT40), .A3(new_n389), .ZN(new_n390));
  AND3_X1   g189(.A1(new_n259), .A2(new_n263), .A3(new_n267), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n271), .B1(new_n259), .B2(new_n263), .ZN(new_n392));
  OAI21_X1  g191(.A(KEYINPUT30), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT30), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n268), .A2(new_n394), .ZN(new_n395));
  AOI22_X1  g194(.A1(new_n393), .A2(new_n395), .B1(new_n334), .B2(new_n329), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n390), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT40), .B1(new_n387), .B2(new_n389), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n343), .B(new_n376), .C1(new_n397), .C2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT36), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n253), .A2(new_n216), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n402), .B1(new_n249), .B2(new_n248), .ZN(new_n403));
  AOI22_X1  g202(.A1(new_n223), .A2(new_n229), .B1(new_n224), .B2(new_n237), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n310), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n239), .A2(new_n292), .A3(new_n254), .ZN(new_n406));
  NAND2_X1  g205(.A1(G227gat), .A2(G233gat), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n405), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT32), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT74), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT74), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n409), .A2(new_n412), .A3(KEYINPUT32), .ZN(new_n413));
  XNOR2_X1  g212(.A(G15gat), .B(G43gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(G71gat), .B(G99gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n411), .A2(new_n413), .A3(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT73), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT33), .ZN(new_n420));
  AND3_X1   g219(.A1(new_n409), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n419), .B1(new_n409), .B2(new_n420), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n418), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT34), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n425), .B1(new_n407), .B2(KEYINPUT75), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n405), .A2(new_n406), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n427), .B1(new_n428), .B2(new_n407), .ZN(new_n429));
  AOI211_X1 g228(.A(new_n408), .B(new_n426), .C1(new_n405), .C2(new_n406), .ZN(new_n430));
  OAI21_X1  g229(.A(KEYINPUT76), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n416), .A2(new_n420), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n431), .B1(new_n410), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n428), .A2(new_n407), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(new_n426), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n428), .A2(new_n407), .A3(new_n427), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n437), .A2(KEYINPUT76), .ZN(new_n438));
  NOR3_X1   g237(.A1(new_n424), .A2(new_n433), .A3(new_n438), .ZN(new_n439));
  OR3_X1    g238(.A1(new_n429), .A2(new_n430), .A3(KEYINPUT76), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n410), .A2(new_n432), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n441), .B1(new_n437), .B2(KEYINPUT76), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n416), .B1(new_n410), .B2(KEYINPUT74), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n443), .B(new_n413), .C1(new_n422), .C2(new_n421), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n440), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n401), .B1(new_n439), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n438), .B1(new_n424), .B2(new_n433), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n442), .A2(new_n444), .A3(new_n440), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n447), .A2(KEYINPUT36), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n393), .A2(new_n395), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n450), .B1(new_n335), .B2(new_n339), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n446), .B(new_n449), .C1(new_n451), .C2(new_n376), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n447), .A2(new_n448), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n376), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n339), .A2(new_n335), .ZN(new_n455));
  AND2_X1   g254(.A1(new_n393), .A2(new_n395), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NOR3_X1   g256(.A1(new_n454), .A2(KEYINPUT35), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT35), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n375), .B1(new_n447), .B2(new_n448), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n459), .B1(new_n460), .B2(new_n451), .ZN(new_n461));
  OAI22_X1  g260(.A1(new_n400), .A2(new_n452), .B1(new_n458), .B2(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(G15gat), .B(G22gat), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT16), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n463), .B1(new_n464), .B2(G1gat), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n465), .B1(G1gat), .B2(new_n463), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n466), .B(G8gat), .ZN(new_n467));
  AND2_X1   g266(.A1(G71gat), .A2(G78gat), .ZN(new_n468));
  NOR2_X1   g267(.A1(G71gat), .A2(G78gat), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(G57gat), .B(G64gat), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(G57gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(G64gat), .ZN(new_n475));
  INV_X1    g274(.A(G64gat), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(G57gat), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  XNOR2_X1  g277(.A(G71gat), .B(G78gat), .ZN(new_n479));
  INV_X1    g278(.A(new_n472), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  AND2_X1   g280(.A1(new_n473), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n467), .B1(KEYINPUT21), .B2(new_n482), .ZN(new_n483));
  XOR2_X1   g282(.A(new_n483), .B(KEYINPUT92), .Z(new_n484));
  NOR2_X1   g283(.A1(new_n482), .A2(KEYINPUT21), .ZN(new_n485));
  NAND2_X1  g284(.A1(G231gat), .A2(G233gat), .ZN(new_n486));
  XOR2_X1   g285(.A(new_n485), .B(new_n486), .Z(new_n487));
  XNOR2_X1  g286(.A(new_n487), .B(G127gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n484), .B(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n490), .B(G155gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(G183gat), .B(G211gat), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n491), .B(new_n492), .ZN(new_n493));
  XOR2_X1   g292(.A(new_n489), .B(new_n493), .Z(new_n494));
  XNOR2_X1  g293(.A(G43gat), .B(G50gat), .ZN(new_n495));
  INV_X1    g294(.A(G29gat), .ZN(new_n496));
  INV_X1    g295(.A(G36gat), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n496), .A2(new_n497), .A3(KEYINPUT14), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT14), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n499), .B1(G29gat), .B2(G36gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n496), .A2(new_n497), .ZN(new_n502));
  OAI211_X1 g301(.A(KEYINPUT15), .B(new_n495), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n501), .B(KEYINPUT89), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n502), .B1(new_n495), .B2(KEYINPUT15), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n505), .B1(KEYINPUT15), .B2(new_n495), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n503), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT17), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI211_X1 g308(.A(KEYINPUT17), .B(new_n503), .C1(new_n504), .C2(new_n506), .ZN(new_n510));
  NAND2_X1  g309(.A1(G99gat), .A2(G106gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT8), .ZN(new_n512));
  NAND2_X1  g311(.A1(G85gat), .A2(G92gat), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT7), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(G85gat), .ZN(new_n516));
  INV_X1    g315(.A(G92gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n512), .A2(new_n515), .A3(new_n518), .A4(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(G99gat), .B(G106gat), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  AOI22_X1  g322(.A1(KEYINPUT8), .A2(new_n511), .B1(new_n516), .B2(new_n517), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n524), .A2(new_n521), .A3(new_n515), .A4(new_n519), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n509), .A2(new_n510), .A3(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT94), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(G232gat), .A2(G233gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(KEYINPUT93), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT41), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n526), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n533), .B1(new_n507), .B2(new_n534), .ZN(new_n535));
  OR2_X1    g334(.A1(new_n535), .A2(KEYINPUT95), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n509), .A2(KEYINPUT94), .A3(new_n510), .A4(new_n526), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n535), .A2(KEYINPUT95), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n529), .A2(new_n536), .A3(new_n537), .A4(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G190gat), .B(G218gat), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT96), .ZN(new_n541));
  OR2_X1    g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n531), .A2(new_n532), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n540), .A2(new_n541), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(G134gat), .B(G162gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n539), .A2(new_n542), .A3(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n547), .B1(new_n539), .B2(new_n542), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(G230gat), .A2(G233gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n525), .A2(KEYINPUT97), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n482), .A2(new_n526), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n473), .A2(new_n481), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n525), .B(new_n523), .C1(new_n556), .C2(KEYINPUT97), .ZN(new_n557));
  AOI21_X1  g356(.A(KEYINPUT10), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT10), .ZN(new_n559));
  NOR3_X1   g358(.A1(new_n526), .A2(new_n556), .A3(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n553), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n555), .A2(new_n557), .ZN(new_n562));
  OR2_X1    g361(.A1(new_n562), .A2(new_n553), .ZN(new_n563));
  XNOR2_X1  g362(.A(G120gat), .B(G148gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(G176gat), .B(G204gat), .ZN(new_n565));
  XOR2_X1   g364(.A(new_n564), .B(new_n565), .Z(new_n566));
  NAND3_X1  g365(.A1(new_n561), .A2(new_n563), .A3(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n562), .A2(new_n559), .ZN(new_n569));
  INV_X1    g368(.A(new_n560), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(new_n553), .B(KEYINPUT98), .Z(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(new_n563), .ZN(new_n575));
  INV_X1    g374(.A(new_n566), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n568), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n494), .A2(new_n552), .A3(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(G8gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n466), .B(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n509), .A2(new_n580), .A3(new_n510), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n467), .A2(new_n507), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(G229gat), .A2(G233gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(KEYINPUT90), .ZN(new_n585));
  OAI21_X1  g384(.A(KEYINPUT91), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n467), .B(new_n507), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n585), .B(KEYINPUT13), .ZN(new_n588));
  AOI22_X1  g387(.A1(new_n586), .A2(KEYINPUT18), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT18), .ZN(new_n590));
  OAI211_X1 g389(.A(KEYINPUT91), .B(new_n590), .C1(new_n583), .C2(new_n585), .ZN(new_n591));
  XNOR2_X1  g390(.A(G113gat), .B(G141gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(G169gat), .B(G197gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(KEYINPUT88), .B(KEYINPUT11), .Z(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(KEYINPUT12), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n589), .A2(new_n591), .A3(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n597), .B1(new_n589), .B2(new_n591), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n578), .A2(new_n601), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n462), .A2(new_n602), .ZN(new_n603));
  AND2_X1   g402(.A1(new_n339), .A2(new_n335), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(KEYINPUT99), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT99), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n455), .A2(new_n606), .ZN(new_n607));
  AND2_X1   g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n603), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(G1gat), .ZN(G1324gat));
  INV_X1    g410(.A(KEYINPUT42), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n603), .A2(new_n450), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT100), .ZN(new_n614));
  XOR2_X1   g413(.A(KEYINPUT16), .B(G8gat), .Z(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n612), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n603), .A2(KEYINPUT42), .A3(new_n450), .A4(new_n615), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT100), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n613), .B(new_n619), .ZN(new_n620));
  NOR3_X1   g419(.A1(new_n620), .A2(KEYINPUT101), .A3(new_n579), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT101), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n622), .B1(new_n614), .B2(G8gat), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n617), .B(new_n618), .C1(new_n621), .C2(new_n623), .ZN(G1325gat));
  INV_X1    g423(.A(G15gat), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n603), .A2(new_n625), .A3(new_n453), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT102), .ZN(new_n627));
  INV_X1    g426(.A(new_n449), .ZN(new_n628));
  AOI21_X1  g427(.A(KEYINPUT36), .B1(new_n447), .B2(new_n448), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n446), .A2(KEYINPUT102), .A3(new_n449), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AND2_X1   g431(.A1(new_n603), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n626), .B1(new_n633), .B2(new_n625), .ZN(G1326gat));
  NAND2_X1  g433(.A1(new_n603), .A2(new_n375), .ZN(new_n635));
  XNOR2_X1  g434(.A(KEYINPUT43), .B(G22gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(G1327gat));
  INV_X1    g436(.A(new_n577), .ZN(new_n638));
  NOR3_X1   g437(.A1(new_n494), .A2(new_n601), .A3(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT104), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT103), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n451), .A2(new_n642), .A3(new_n376), .ZN(new_n643));
  AOI21_X1  g442(.A(KEYINPUT103), .B1(new_n457), .B2(new_n375), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n399), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n641), .B1(new_n645), .B2(new_n632), .ZN(new_n646));
  AND3_X1   g445(.A1(new_n446), .A2(KEYINPUT102), .A3(new_n449), .ZN(new_n647));
  AOI21_X1  g446(.A(KEYINPUT102), .B1(new_n446), .B2(new_n449), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n642), .B1(new_n451), .B2(new_n376), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n457), .A2(KEYINPUT103), .A3(new_n375), .ZN(new_n651));
  OR2_X1    g450(.A1(new_n341), .A2(new_n274), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n275), .B1(new_n652), .B2(KEYINPUT38), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n375), .B1(new_n653), .B2(new_n604), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n385), .A2(new_n386), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n655), .A2(new_n333), .A3(new_n389), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT40), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n658), .A2(new_n390), .A3(new_n396), .ZN(new_n659));
  AOI22_X1  g458(.A1(new_n650), .A2(new_n651), .B1(new_n654), .B2(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n649), .A2(new_n660), .A3(KEYINPUT104), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n458), .A2(new_n461), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n646), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n552), .A2(KEYINPUT44), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT44), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n666), .B1(new_n462), .B2(new_n551), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n640), .B1(new_n665), .B2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(G29gat), .B1(new_n670), .B2(new_n608), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n462), .A2(new_n551), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n672), .A2(new_n640), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n673), .A2(new_n496), .A3(new_n609), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT45), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n671), .A2(new_n675), .ZN(G1328gat));
  NAND3_X1  g475(.A1(new_n673), .A2(new_n497), .A3(new_n450), .ZN(new_n677));
  XOR2_X1   g476(.A(new_n677), .B(KEYINPUT46), .Z(new_n678));
  OAI21_X1  g477(.A(G36gat), .B1(new_n670), .B2(new_n456), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(G1329gat));
  AND2_X1   g479(.A1(new_n673), .A2(new_n453), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n681), .A2(G43gat), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n632), .A2(G43gat), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n682), .B1(new_n670), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(KEYINPUT47), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT47), .ZN(new_n686));
  OAI211_X1 g485(.A(new_n682), .B(new_n686), .C1(new_n670), .C2(new_n683), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n685), .A2(new_n687), .ZN(G1330gat));
  INV_X1    g487(.A(KEYINPUT48), .ZN(new_n689));
  INV_X1    g488(.A(G50gat), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n690), .B1(new_n669), .B2(new_n375), .ZN(new_n691));
  NOR4_X1   g490(.A1(new_n672), .A2(G50gat), .A3(new_n376), .A4(new_n640), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n689), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT105), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n694), .B1(new_n669), .B2(new_n375), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n667), .B1(new_n663), .B2(new_n664), .ZN(new_n696));
  NOR4_X1   g495(.A1(new_n696), .A2(KEYINPUT105), .A3(new_n376), .A4(new_n640), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n695), .A2(new_n697), .A3(new_n690), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n692), .A2(new_n689), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n693), .B1(new_n698), .B2(new_n699), .ZN(G1331gat));
  INV_X1    g499(.A(new_n663), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n494), .A2(new_n601), .A3(new_n552), .A4(new_n638), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(new_n609), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(G57gat), .ZN(G1332gat));
  OR2_X1    g504(.A1(new_n701), .A2(new_n702), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT49), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n450), .B1(new_n707), .B2(new_n476), .ZN(new_n708));
  OAI21_X1  g507(.A(KEYINPUT106), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  OR4_X1    g508(.A1(KEYINPUT106), .A2(new_n701), .A3(new_n702), .A4(new_n708), .ZN(new_n710));
  NOR2_X1   g509(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n711));
  AND3_X1   g510(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n711), .B1(new_n709), .B2(new_n710), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n712), .A2(new_n713), .ZN(G1333gat));
  OAI21_X1  g513(.A(G71gat), .B1(new_n706), .B2(new_n649), .ZN(new_n715));
  INV_X1    g514(.A(G71gat), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n703), .A2(new_n716), .A3(new_n453), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT50), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n715), .A2(new_n717), .A3(KEYINPUT50), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(G1334gat));
  NAND2_X1  g521(.A1(new_n703), .A2(new_n375), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(G78gat), .ZN(G1335gat));
  INV_X1    g523(.A(new_n600), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n598), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n494), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(new_n638), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n728), .B1(new_n665), .B2(new_n668), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(G85gat), .B1(new_n730), .B2(new_n608), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT51), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n732), .A2(KEYINPUT107), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n727), .ZN(new_n735));
  AOI211_X1 g534(.A(new_n552), .B(new_n735), .C1(KEYINPUT107), .C2(new_n732), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n734), .B1(new_n663), .B2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n663), .A2(new_n734), .A3(new_n736), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n609), .A2(new_n516), .A3(new_n638), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n731), .B1(new_n740), .B2(new_n741), .ZN(G1336gat));
  AOI21_X1  g541(.A(new_n517), .B1(new_n729), .B2(new_n450), .ZN(new_n743));
  INV_X1    g542(.A(new_n739), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n450), .A2(new_n517), .A3(new_n638), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT108), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n744), .A2(new_n737), .A3(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(KEYINPUT52), .B1(new_n743), .B2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT109), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n749), .B1(new_n729), .B2(new_n450), .ZN(new_n750));
  NOR4_X1   g549(.A1(new_n696), .A2(KEYINPUT109), .A3(new_n456), .A4(new_n728), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n750), .A2(new_n751), .A3(new_n517), .ZN(new_n752));
  OR2_X1    g551(.A1(new_n747), .A2(KEYINPUT52), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n748), .B1(new_n752), .B2(new_n753), .ZN(G1337gat));
  OAI21_X1  g553(.A(G99gat), .B1(new_n730), .B2(new_n649), .ZN(new_n755));
  INV_X1    g554(.A(G99gat), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n453), .A2(new_n756), .A3(new_n638), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n755), .B1(new_n740), .B2(new_n757), .ZN(G1338gat));
  INV_X1    g557(.A(G106gat), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n759), .B1(new_n729), .B2(new_n375), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT53), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n577), .A2(G106gat), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n375), .A2(new_n763), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n744), .A2(new_n737), .A3(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n761), .A2(new_n762), .A3(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(KEYINPUT53), .B1(new_n760), .B2(new_n765), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(G1339gat));
  NAND4_X1  g568(.A1(new_n494), .A2(new_n601), .A3(new_n552), .A4(new_n577), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n583), .A2(new_n585), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n587), .A2(new_n588), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n596), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n598), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n552), .A2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT111), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT54), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n571), .A2(new_n777), .A3(new_n573), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n778), .A2(KEYINPUT55), .A3(new_n576), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT110), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n777), .B1(new_n571), .B2(new_n553), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n558), .A2(new_n573), .A3(new_n560), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n780), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n561), .A2(KEYINPUT54), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n785), .A2(KEYINPUT110), .A3(new_n782), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n779), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(new_n567), .ZN(new_n788));
  OAI21_X1  g587(.A(KEYINPUT110), .B1(new_n785), .B2(new_n782), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n783), .A2(new_n780), .A3(KEYINPUT54), .A4(new_n561), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n778), .A2(new_n576), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT55), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n776), .B1(new_n788), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n568), .B1(new_n791), .B2(new_n779), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n792), .B1(new_n789), .B2(new_n790), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n796), .B(KEYINPUT111), .C1(KEYINPUT55), .C2(new_n797), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n775), .A2(new_n795), .A3(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n795), .A2(new_n726), .A3(new_n798), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n598), .A2(new_n638), .A3(new_n773), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(KEYINPUT112), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT112), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n598), .A2(new_n638), .A3(new_n803), .A4(new_n773), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n800), .A2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT113), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n551), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n800), .A2(new_n805), .A3(KEYINPUT113), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n799), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n770), .B1(new_n810), .B2(new_n494), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n812), .A2(new_n454), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n608), .A2(new_n450), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(G113gat), .B1(new_n815), .B2(new_n601), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n601), .A2(G113gat), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n817), .B(KEYINPUT114), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n816), .B1(new_n815), .B2(new_n818), .ZN(G1340gat));
  NOR2_X1   g618(.A1(new_n815), .A2(new_n577), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n820), .A2(G120gat), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n821), .B1(new_n279), .B2(new_n820), .ZN(G1341gat));
  INV_X1    g621(.A(new_n494), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n815), .A2(new_n823), .ZN(new_n824));
  XOR2_X1   g623(.A(new_n824), .B(G127gat), .Z(G1342gat));
  NAND4_X1  g624(.A1(new_n813), .A2(new_n456), .A3(new_n551), .A4(new_n609), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(G134gat), .ZN(new_n827));
  XNOR2_X1  g626(.A(new_n827), .B(KEYINPUT115), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT116), .ZN(new_n829));
  OAI22_X1  g628(.A1(new_n826), .A2(G134gat), .B1(new_n829), .B2(KEYINPUT56), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(KEYINPUT56), .ZN(new_n831));
  OR2_X1    g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(new_n831), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n828), .A2(new_n832), .A3(new_n833), .ZN(G1343gat));
  NOR3_X1   g633(.A1(new_n632), .A2(new_n450), .A3(new_n608), .ZN(new_n835));
  AOI21_X1  g634(.A(KEYINPUT57), .B1(new_n811), .B2(new_n375), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n375), .A2(KEYINPUT57), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n796), .B1(KEYINPUT55), .B2(new_n797), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n801), .B1(new_n601), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n799), .B1(new_n552), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n841), .A2(new_n494), .ZN(new_n842));
  INV_X1    g641(.A(new_n770), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n838), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n835), .B1(new_n836), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(G141gat), .B1(new_n846), .B2(new_n601), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n812), .A2(new_n376), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n835), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n601), .A2(G141gat), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n850), .B(KEYINPUT117), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n847), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(KEYINPUT58), .ZN(G1344gat));
  OAI211_X1 g652(.A(new_n551), .B(new_n796), .C1(KEYINPUT55), .C2(new_n797), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n854), .A2(KEYINPUT118), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n774), .B1(new_n854), .B2(KEYINPUT118), .ZN(new_n856));
  AOI22_X1  g655(.A1(new_n855), .A2(new_n856), .B1(new_n840), .B2(new_n552), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n770), .B1(new_n857), .B2(new_n494), .ZN(new_n858));
  AOI21_X1  g657(.A(KEYINPUT57), .B1(new_n858), .B2(new_n375), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n859), .B1(new_n811), .B2(new_n838), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  AND3_X1   g660(.A1(new_n861), .A2(new_n638), .A3(new_n835), .ZN(new_n862));
  INV_X1    g661(.A(G148gat), .ZN(new_n863));
  OAI21_X1  g662(.A(KEYINPUT59), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n863), .A2(KEYINPUT59), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n865), .B1(new_n846), .B2(new_n577), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n638), .A2(new_n863), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n867), .B1(new_n849), .B2(new_n868), .ZN(G1345gat));
  NOR3_X1   g668(.A1(new_n846), .A2(new_n294), .A3(new_n823), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n849), .A2(KEYINPUT119), .A3(new_n823), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n871), .A2(G155gat), .ZN(new_n872));
  OAI21_X1  g671(.A(KEYINPUT119), .B1(new_n849), .B2(new_n823), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n870), .B1(new_n872), .B2(new_n873), .ZN(G1346gat));
  NOR4_X1   g673(.A1(new_n608), .A2(G162gat), .A3(new_n450), .A4(new_n552), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n848), .A2(new_n649), .A3(new_n875), .ZN(new_n876));
  XNOR2_X1  g675(.A(new_n876), .B(KEYINPUT120), .ZN(new_n877));
  OAI21_X1  g676(.A(G162gat), .B1(new_n846), .B2(new_n552), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(G1347gat));
  NOR2_X1   g678(.A1(new_n812), .A2(new_n609), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n460), .A2(new_n450), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(G169gat), .B1(new_n884), .B2(new_n726), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n813), .A2(new_n450), .A3(new_n608), .ZN(new_n886));
  INV_X1    g685(.A(G169gat), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n886), .A2(new_n887), .A3(new_n601), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n885), .A2(new_n888), .ZN(G1348gat));
  OAI21_X1  g688(.A(G176gat), .B1(new_n886), .B2(new_n577), .ZN(new_n890));
  OR2_X1    g689(.A1(new_n577), .A2(G176gat), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n890), .B1(new_n883), .B2(new_n891), .ZN(G1349gat));
  OAI21_X1  g691(.A(G183gat), .B1(new_n886), .B2(new_n823), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n494), .A2(new_n240), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n893), .B1(new_n883), .B2(new_n894), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g695(.A(G190gat), .B1(new_n886), .B2(new_n552), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n897), .B(KEYINPUT61), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n884), .A2(new_n241), .A3(new_n551), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(G1351gat));
  NOR3_X1   g699(.A1(new_n632), .A2(new_n456), .A3(new_n376), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n880), .A2(new_n901), .ZN(new_n902));
  OR3_X1    g701(.A1(new_n902), .A2(G197gat), .A3(new_n601), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n904));
  OR2_X1    g703(.A1(new_n860), .A2(KEYINPUT121), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n860), .A2(KEYINPUT121), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n608), .A2(new_n450), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n632), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n905), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n904), .B1(new_n909), .B2(new_n601), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(G197gat), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n909), .A2(new_n904), .A3(new_n601), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n903), .B1(new_n911), .B2(new_n912), .ZN(G1352gat));
  NOR2_X1   g712(.A1(new_n577), .A2(G204gat), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(KEYINPUT123), .B1(new_n902), .B2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT123), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n880), .A2(new_n917), .A3(new_n901), .A4(new_n914), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n919), .A2(KEYINPUT62), .ZN(new_n920));
  OAI21_X1  g719(.A(G204gat), .B1(new_n909), .B2(new_n577), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n916), .A2(KEYINPUT62), .A3(new_n918), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(G1353gat));
  NAND4_X1  g722(.A1(new_n880), .A2(new_n205), .A3(new_n494), .A4(new_n901), .ZN(new_n924));
  NAND2_X1  g723(.A1(KEYINPUT125), .A2(KEYINPUT63), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT124), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n908), .A2(new_n494), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n927), .B1(new_n860), .B2(new_n928), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n632), .A2(new_n907), .A3(new_n823), .ZN(new_n930));
  AND3_X1   g729(.A1(new_n800), .A2(KEYINPUT113), .A3(new_n805), .ZN(new_n931));
  AOI21_X1  g730(.A(KEYINPUT113), .B1(new_n800), .B2(new_n805), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n931), .A2(new_n932), .A3(new_n551), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n823), .B1(new_n933), .B2(new_n799), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n837), .B1(new_n934), .B2(new_n770), .ZN(new_n935));
  OAI211_X1 g734(.A(KEYINPUT124), .B(new_n930), .C1(new_n935), .C2(new_n859), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n929), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g736(.A(G211gat), .B1(KEYINPUT125), .B2(KEYINPUT63), .ZN(new_n938));
  INV_X1    g737(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n926), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  AOI211_X1 g739(.A(new_n925), .B(new_n938), .C1(new_n929), .C2(new_n936), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n924), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT126), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI211_X1 g743(.A(KEYINPUT126), .B(new_n924), .C1(new_n940), .C2(new_n941), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(G1354gat));
  NOR3_X1   g745(.A1(new_n909), .A2(new_n206), .A3(new_n552), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n880), .A2(new_n551), .A3(new_n901), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n947), .B1(new_n206), .B2(new_n948), .ZN(G1355gat));
endmodule


