

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583;

  XNOR2_X1 U322 ( .A(n360), .B(n326), .ZN(n327) );
  XOR2_X1 U323 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n290) );
  AND2_X1 U324 ( .A1(G227GAT), .A2(G233GAT), .ZN(n291) );
  INV_X1 U325 ( .A(KEYINPUT97), .ZN(n370) );
  NOR2_X1 U326 ( .A1(n542), .A2(n541), .ZN(n543) );
  NOR2_X1 U327 ( .A1(n506), .A2(n552), .ZN(n507) );
  XOR2_X1 U328 ( .A(KEYINPUT11), .B(KEYINPUT81), .Z(n293) );
  AND2_X1 U329 ( .A1(n508), .A2(n507), .ZN(n509) );
  XNOR2_X1 U330 ( .A(n362), .B(n294), .ZN(n295) );
  XNOR2_X1 U331 ( .A(n434), .B(n291), .ZN(n326) );
  XNOR2_X1 U332 ( .A(n296), .B(n295), .ZN(n298) );
  XNOR2_X1 U333 ( .A(n546), .B(KEYINPUT65), .ZN(n567) );
  XNOR2_X1 U334 ( .A(n358), .B(n357), .ZN(n566) );
  XNOR2_X1 U335 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U336 ( .A(n304), .B(n303), .ZN(n309) );
  XOR2_X1 U337 ( .A(n339), .B(n338), .Z(n549) );
  XNOR2_X1 U338 ( .A(n447), .B(n446), .ZN(n474) );
  XNOR2_X1 U339 ( .A(n448), .B(KEYINPUT40), .ZN(n449) );
  XNOR2_X1 U340 ( .A(n450), .B(n449), .ZN(G1330GAT) );
  XNOR2_X1 U341 ( .A(G92GAT), .B(KEYINPUT79), .ZN(n292) );
  XOR2_X1 U342 ( .A(n293), .B(n292), .Z(n296) );
  XOR2_X1 U343 ( .A(G36GAT), .B(G190GAT), .Z(n362) );
  XNOR2_X1 U344 ( .A(G218GAT), .B(G106GAT), .ZN(n294) );
  XNOR2_X1 U345 ( .A(G99GAT), .B(G85GAT), .ZN(n297) );
  XNOR2_X1 U346 ( .A(n297), .B(KEYINPUT74), .ZN(n440) );
  XOR2_X1 U347 ( .A(n298), .B(n440), .Z(n304) );
  XOR2_X1 U348 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n300) );
  NAND2_X1 U349 ( .A1(G232GAT), .A2(G233GAT), .ZN(n299) );
  XOR2_X1 U350 ( .A(n300), .B(n299), .Z(n302) );
  XOR2_X1 U351 ( .A(G50GAT), .B(G162GAT), .Z(n341) );
  XOR2_X1 U352 ( .A(G134GAT), .B(KEYINPUT80), .Z(n382) );
  XNOR2_X1 U353 ( .A(n341), .B(n382), .ZN(n301) );
  XOR2_X1 U354 ( .A(KEYINPUT69), .B(KEYINPUT8), .Z(n306) );
  XNOR2_X1 U355 ( .A(G43GAT), .B(G29GAT), .ZN(n305) );
  XNOR2_X1 U356 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U357 ( .A(KEYINPUT7), .B(n307), .Z(n421) );
  XNOR2_X1 U358 ( .A(n421), .B(KEYINPUT66), .ZN(n308) );
  XOR2_X1 U359 ( .A(n309), .B(n308), .Z(n563) );
  XOR2_X1 U360 ( .A(n563), .B(KEYINPUT36), .Z(n580) );
  XOR2_X1 U361 ( .A(G155GAT), .B(G71GAT), .Z(n311) );
  XNOR2_X1 U362 ( .A(G22GAT), .B(G127GAT), .ZN(n310) );
  XNOR2_X1 U363 ( .A(n311), .B(n310), .ZN(n324) );
  XOR2_X1 U364 ( .A(G57GAT), .B(KEYINPUT13), .Z(n431) );
  XOR2_X1 U365 ( .A(G8GAT), .B(G183GAT), .Z(n359) );
  XOR2_X1 U366 ( .A(n431), .B(n359), .Z(n313) );
  NAND2_X1 U367 ( .A1(G231GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U368 ( .A(n313), .B(n312), .ZN(n317) );
  XOR2_X1 U369 ( .A(KEYINPUT83), .B(KEYINPUT14), .Z(n315) );
  XNOR2_X1 U370 ( .A(KEYINPUT82), .B(KEYINPUT15), .ZN(n314) );
  XNOR2_X1 U371 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U372 ( .A(n317), .B(n316), .Z(n322) );
  XOR2_X1 U373 ( .A(G15GAT), .B(G1GAT), .Z(n413) );
  XOR2_X1 U374 ( .A(KEYINPUT12), .B(G64GAT), .Z(n319) );
  XNOR2_X1 U375 ( .A(G211GAT), .B(G78GAT), .ZN(n318) );
  XNOR2_X1 U376 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U377 ( .A(n413), .B(n320), .ZN(n321) );
  XNOR2_X1 U378 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U379 ( .A(n324), .B(n323), .Z(n576) );
  XNOR2_X1 U380 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n325) );
  XNOR2_X1 U381 ( .A(n290), .B(n325), .ZN(n360) );
  XOR2_X1 U382 ( .A(G120GAT), .B(G71GAT), .Z(n434) );
  XOR2_X1 U383 ( .A(n327), .B(G176GAT), .Z(n331) );
  XOR2_X1 U384 ( .A(G127GAT), .B(KEYINPUT0), .Z(n329) );
  XNOR2_X1 U385 ( .A(G113GAT), .B(KEYINPUT85), .ZN(n328) );
  XNOR2_X1 U386 ( .A(n329), .B(n328), .ZN(n381) );
  XNOR2_X1 U387 ( .A(G15GAT), .B(n381), .ZN(n330) );
  XNOR2_X1 U388 ( .A(n331), .B(n330), .ZN(n339) );
  XOR2_X1 U389 ( .A(G190GAT), .B(G134GAT), .Z(n333) );
  XNOR2_X1 U390 ( .A(G43GAT), .B(G99GAT), .ZN(n332) );
  XNOR2_X1 U391 ( .A(n333), .B(n332), .ZN(n337) );
  XOR2_X1 U392 ( .A(KEYINPUT86), .B(KEYINPUT87), .Z(n335) );
  XNOR2_X1 U393 ( .A(KEYINPUT20), .B(G183GAT), .ZN(n334) );
  XNOR2_X1 U394 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U395 ( .A(n337), .B(n336), .Z(n338) );
  XNOR2_X1 U396 ( .A(G106GAT), .B(G78GAT), .ZN(n340) );
  XNOR2_X1 U397 ( .A(n340), .B(G148GAT), .ZN(n441) );
  XOR2_X1 U398 ( .A(n441), .B(n341), .Z(n346) );
  XOR2_X1 U399 ( .A(G141GAT), .B(G22GAT), .Z(n420) );
  XOR2_X1 U400 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n343) );
  XNOR2_X1 U401 ( .A(KEYINPUT89), .B(G155GAT), .ZN(n342) );
  XNOR2_X1 U402 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U403 ( .A(KEYINPUT90), .B(n344), .Z(n386) );
  XNOR2_X1 U404 ( .A(n420), .B(n386), .ZN(n345) );
  XNOR2_X1 U405 ( .A(n346), .B(n345), .ZN(n350) );
  XOR2_X1 U406 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n348) );
  NAND2_X1 U407 ( .A1(G228GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U408 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U409 ( .A(n350), .B(n349), .Z(n356) );
  XNOR2_X1 U410 ( .A(G211GAT), .B(G218GAT), .ZN(n351) );
  XNOR2_X1 U411 ( .A(n351), .B(KEYINPUT21), .ZN(n352) );
  XOR2_X1 U412 ( .A(n352), .B(KEYINPUT88), .Z(n354) );
  XNOR2_X1 U413 ( .A(G197GAT), .B(G204GAT), .ZN(n353) );
  XNOR2_X1 U414 ( .A(n354), .B(n353), .ZN(n368) );
  XNOR2_X1 U415 ( .A(n368), .B(KEYINPUT22), .ZN(n355) );
  XNOR2_X1 U416 ( .A(n356), .B(n355), .ZN(n547) );
  NOR2_X1 U417 ( .A1(n549), .A2(n547), .ZN(n358) );
  XNOR2_X1 U418 ( .A(KEYINPUT96), .B(KEYINPUT26), .ZN(n357) );
  XNOR2_X1 U419 ( .A(KEYINPUT27), .B(KEYINPUT95), .ZN(n369) );
  XNOR2_X1 U420 ( .A(n360), .B(n359), .ZN(n366) );
  XNOR2_X1 U421 ( .A(G176GAT), .B(G92GAT), .ZN(n361) );
  XNOR2_X1 U422 ( .A(n361), .B(G64GAT), .ZN(n435) );
  XOR2_X1 U423 ( .A(n362), .B(n435), .Z(n364) );
  NAND2_X1 U424 ( .A1(G226GAT), .A2(G233GAT), .ZN(n363) );
  XNOR2_X1 U425 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U426 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U427 ( .A(n368), .B(n367), .Z(n490) );
  XOR2_X1 U428 ( .A(n369), .B(n490), .Z(n400) );
  AND2_X1 U429 ( .A1(n566), .A2(n400), .ZN(n526) );
  XNOR2_X1 U430 ( .A(n526), .B(n370), .ZN(n399) );
  XNOR2_X1 U431 ( .A(KEYINPUT99), .B(KEYINPUT25), .ZN(n374) );
  NAND2_X1 U432 ( .A1(n490), .A2(n549), .ZN(n371) );
  NAND2_X1 U433 ( .A1(n371), .A2(n547), .ZN(n372) );
  XNOR2_X1 U434 ( .A(n372), .B(KEYINPUT98), .ZN(n373) );
  XNOR2_X1 U435 ( .A(n374), .B(n373), .ZN(n397) );
  XOR2_X1 U436 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n376) );
  XNOR2_X1 U437 ( .A(G1GAT), .B(KEYINPUT5), .ZN(n375) );
  XNOR2_X1 U438 ( .A(n376), .B(n375), .ZN(n380) );
  XOR2_X1 U439 ( .A(G57GAT), .B(KEYINPUT1), .Z(n378) );
  XNOR2_X1 U440 ( .A(KEYINPUT91), .B(KEYINPUT6), .ZN(n377) );
  XNOR2_X1 U441 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U442 ( .A(n380), .B(n379), .Z(n388) );
  XOR2_X1 U443 ( .A(n382), .B(n381), .Z(n384) );
  NAND2_X1 U444 ( .A1(G225GAT), .A2(G233GAT), .ZN(n383) );
  XNOR2_X1 U445 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U446 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U447 ( .A(n388), .B(n387), .ZN(n396) );
  XOR2_X1 U448 ( .A(KEYINPUT94), .B(KEYINPUT4), .Z(n390) );
  XNOR2_X1 U449 ( .A(G141GAT), .B(G148GAT), .ZN(n389) );
  XNOR2_X1 U450 ( .A(n390), .B(n389), .ZN(n394) );
  XOR2_X1 U451 ( .A(G85GAT), .B(G162GAT), .Z(n392) );
  XNOR2_X1 U452 ( .A(G29GAT), .B(G120GAT), .ZN(n391) );
  XNOR2_X1 U453 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U454 ( .A(n394), .B(n393), .Z(n395) );
  XOR2_X1 U455 ( .A(n396), .B(n395), .Z(n488) );
  INV_X1 U456 ( .A(n488), .ZN(n544) );
  NAND2_X1 U457 ( .A1(n397), .A2(n544), .ZN(n398) );
  NOR2_X1 U458 ( .A1(n399), .A2(n398), .ZN(n403) );
  XOR2_X1 U459 ( .A(n547), .B(KEYINPUT28), .Z(n493) );
  INV_X1 U460 ( .A(n493), .ZN(n473) );
  NAND2_X1 U461 ( .A1(n400), .A2(n473), .ZN(n512) );
  NOR2_X1 U462 ( .A1(n512), .A2(n549), .ZN(n401) );
  NOR2_X1 U463 ( .A1(n544), .A2(n401), .ZN(n402) );
  NOR2_X1 U464 ( .A1(n403), .A2(n402), .ZN(n453) );
  NAND2_X1 U465 ( .A1(n576), .A2(n453), .ZN(n404) );
  XOR2_X1 U466 ( .A(KEYINPUT105), .B(n404), .Z(n405) );
  NOR2_X1 U467 ( .A1(n580), .A2(n405), .ZN(n407) );
  XNOR2_X1 U468 ( .A(KEYINPUT106), .B(KEYINPUT37), .ZN(n406) );
  XNOR2_X1 U469 ( .A(n407), .B(n406), .ZN(n487) );
  XOR2_X1 U470 ( .A(KEYINPUT68), .B(KEYINPUT71), .Z(n409) );
  XNOR2_X1 U471 ( .A(KEYINPUT67), .B(KEYINPUT30), .ZN(n408) );
  XNOR2_X1 U472 ( .A(n409), .B(n408), .ZN(n425) );
  XOR2_X1 U473 ( .A(G8GAT), .B(G197GAT), .Z(n411) );
  XNOR2_X1 U474 ( .A(G50GAT), .B(G36GAT), .ZN(n410) );
  XNOR2_X1 U475 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U476 ( .A(n412), .B(G113GAT), .Z(n415) );
  XNOR2_X1 U477 ( .A(G169GAT), .B(n413), .ZN(n414) );
  XNOR2_X1 U478 ( .A(n415), .B(n414), .ZN(n419) );
  XOR2_X1 U479 ( .A(KEYINPUT70), .B(KEYINPUT29), .Z(n417) );
  NAND2_X1 U480 ( .A1(G229GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U481 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U482 ( .A(n419), .B(n418), .Z(n423) );
  XNOR2_X1 U483 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U484 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U485 ( .A(n425), .B(n424), .ZN(n568) );
  INV_X1 U486 ( .A(n568), .ZN(n552) );
  XOR2_X1 U487 ( .A(KEYINPUT31), .B(KEYINPUT78), .Z(n427) );
  XNOR2_X1 U488 ( .A(KEYINPUT72), .B(KEYINPUT77), .ZN(n426) );
  XNOR2_X1 U489 ( .A(n427), .B(n426), .ZN(n445) );
  XOR2_X1 U490 ( .A(KEYINPUT76), .B(KEYINPUT32), .Z(n429) );
  XNOR2_X1 U491 ( .A(KEYINPUT73), .B(KEYINPUT33), .ZN(n428) );
  XNOR2_X1 U492 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U493 ( .A(n430), .B(KEYINPUT75), .Z(n433) );
  XNOR2_X1 U494 ( .A(G204GAT), .B(n431), .ZN(n432) );
  XNOR2_X1 U495 ( .A(n433), .B(n432), .ZN(n439) );
  XOR2_X1 U496 ( .A(n435), .B(n434), .Z(n437) );
  NAND2_X1 U497 ( .A1(G230GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U498 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U499 ( .A(n439), .B(n438), .Z(n443) );
  XNOR2_X1 U500 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U501 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U502 ( .A(n445), .B(n444), .Z(n572) );
  NAND2_X1 U503 ( .A1(n552), .A2(n572), .ZN(n456) );
  NOR2_X1 U504 ( .A1(n487), .A2(n456), .ZN(n447) );
  XNOR2_X1 U505 ( .A(KEYINPUT38), .B(KEYINPUT107), .ZN(n446) );
  INV_X1 U506 ( .A(n549), .ZN(n513) );
  NOR2_X1 U507 ( .A1(n474), .A2(n513), .ZN(n450) );
  INV_X1 U508 ( .A(G43GAT), .ZN(n448) );
  XOR2_X1 U509 ( .A(KEYINPUT34), .B(KEYINPUT102), .Z(n459) );
  XOR2_X1 U510 ( .A(KEYINPUT84), .B(KEYINPUT16), .Z(n452) );
  INV_X1 U511 ( .A(n563), .ZN(n538) );
  INV_X1 U512 ( .A(n576), .ZN(n560) );
  NAND2_X1 U513 ( .A1(n538), .A2(n560), .ZN(n451) );
  XNOR2_X1 U514 ( .A(n452), .B(n451), .ZN(n454) );
  NAND2_X1 U515 ( .A1(n454), .A2(n453), .ZN(n455) );
  XNOR2_X1 U516 ( .A(n455), .B(KEYINPUT100), .ZN(n477) );
  NOR2_X1 U517 ( .A1(n477), .A2(n456), .ZN(n457) );
  XOR2_X1 U518 ( .A(KEYINPUT101), .B(n457), .Z(n465) );
  NAND2_X1 U519 ( .A1(n465), .A2(n488), .ZN(n458) );
  XNOR2_X1 U520 ( .A(n459), .B(n458), .ZN(n460) );
  XOR2_X1 U521 ( .A(G1GAT), .B(n460), .Z(G1324GAT) );
  NAND2_X1 U522 ( .A1(n465), .A2(n490), .ZN(n461) );
  XNOR2_X1 U523 ( .A(n461), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U524 ( .A(KEYINPUT35), .B(KEYINPUT103), .Z(n463) );
  NAND2_X1 U525 ( .A1(n465), .A2(n549), .ZN(n462) );
  XNOR2_X1 U526 ( .A(n463), .B(n462), .ZN(n464) );
  XOR2_X1 U527 ( .A(G15GAT), .B(n464), .Z(G1326GAT) );
  NAND2_X1 U528 ( .A1(n465), .A2(n493), .ZN(n466) );
  XNOR2_X1 U529 ( .A(n466), .B(KEYINPUT104), .ZN(n467) );
  XNOR2_X1 U530 ( .A(G22GAT), .B(n467), .ZN(G1327GAT) );
  NOR2_X1 U531 ( .A1(n474), .A2(n544), .ZN(n469) );
  XNOR2_X1 U532 ( .A(KEYINPUT108), .B(KEYINPUT39), .ZN(n468) );
  XNOR2_X1 U533 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U534 ( .A(G29GAT), .B(n470), .ZN(G1328GAT) );
  INV_X1 U535 ( .A(n490), .ZN(n542) );
  NOR2_X1 U536 ( .A1(n474), .A2(n542), .ZN(n472) );
  XNOR2_X1 U537 ( .A(G36GAT), .B(KEYINPUT109), .ZN(n471) );
  XNOR2_X1 U538 ( .A(n472), .B(n471), .ZN(G1329GAT) );
  NOR2_X1 U539 ( .A1(n474), .A2(n473), .ZN(n475) );
  XOR2_X1 U540 ( .A(G50GAT), .B(n475), .Z(G1331GAT) );
  XNOR2_X1 U541 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n479) );
  XOR2_X1 U542 ( .A(KEYINPUT41), .B(KEYINPUT64), .Z(n476) );
  XNOR2_X1 U543 ( .A(n572), .B(n476), .ZN(n528) );
  INV_X1 U544 ( .A(n528), .ZN(n557) );
  NAND2_X1 U545 ( .A1(n557), .A2(n568), .ZN(n486) );
  NOR2_X1 U546 ( .A1(n477), .A2(n486), .ZN(n483) );
  NAND2_X1 U547 ( .A1(n488), .A2(n483), .ZN(n478) );
  XNOR2_X1 U548 ( .A(n479), .B(n478), .ZN(G1332GAT) );
  NAND2_X1 U549 ( .A1(n483), .A2(n490), .ZN(n480) );
  XNOR2_X1 U550 ( .A(n480), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U551 ( .A1(n483), .A2(n549), .ZN(n481) );
  XNOR2_X1 U552 ( .A(n481), .B(KEYINPUT110), .ZN(n482) );
  XNOR2_X1 U553 ( .A(G71GAT), .B(n482), .ZN(G1334GAT) );
  XOR2_X1 U554 ( .A(G78GAT), .B(KEYINPUT43), .Z(n485) );
  NAND2_X1 U555 ( .A1(n483), .A2(n493), .ZN(n484) );
  XNOR2_X1 U556 ( .A(n485), .B(n484), .ZN(G1335GAT) );
  NOR2_X1 U557 ( .A1(n487), .A2(n486), .ZN(n494) );
  NAND2_X1 U558 ( .A1(n494), .A2(n488), .ZN(n489) );
  XNOR2_X1 U559 ( .A(n489), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U560 ( .A1(n494), .A2(n490), .ZN(n491) );
  XNOR2_X1 U561 ( .A(n491), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U562 ( .A1(n494), .A2(n549), .ZN(n492) );
  XNOR2_X1 U563 ( .A(n492), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U564 ( .A(KEYINPUT44), .B(KEYINPUT112), .ZN(n498) );
  XOR2_X1 U565 ( .A(G106GAT), .B(KEYINPUT111), .Z(n496) );
  NAND2_X1 U566 ( .A1(n494), .A2(n493), .ZN(n495) );
  XNOR2_X1 U567 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U568 ( .A(n498), .B(n497), .ZN(G1339GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT113), .B(KEYINPUT47), .Z(n503) );
  NOR2_X1 U570 ( .A1(n568), .A2(n528), .ZN(n499) );
  XNOR2_X1 U571 ( .A(n499), .B(KEYINPUT46), .ZN(n500) );
  NOR2_X1 U572 ( .A1(n560), .A2(n500), .ZN(n501) );
  NAND2_X1 U573 ( .A1(n501), .A2(n538), .ZN(n502) );
  XNOR2_X1 U574 ( .A(n503), .B(n502), .ZN(n510) );
  NOR2_X1 U575 ( .A1(n576), .A2(n580), .ZN(n505) );
  XNOR2_X1 U576 ( .A(KEYINPUT45), .B(KEYINPUT114), .ZN(n504) );
  XNOR2_X1 U577 ( .A(n505), .B(n504), .ZN(n508) );
  INV_X1 U578 ( .A(n572), .ZN(n506) );
  NOR2_X1 U579 ( .A1(n510), .A2(n509), .ZN(n511) );
  XNOR2_X1 U580 ( .A(KEYINPUT48), .B(n511), .ZN(n541) );
  NOR2_X1 U581 ( .A1(n544), .A2(n541), .ZN(n525) );
  NOR2_X1 U582 ( .A1(n513), .A2(n512), .ZN(n514) );
  NAND2_X1 U583 ( .A1(n525), .A2(n514), .ZN(n515) );
  XNOR2_X1 U584 ( .A(KEYINPUT115), .B(n515), .ZN(n522) );
  NAND2_X1 U585 ( .A1(n522), .A2(n552), .ZN(n516) );
  XNOR2_X1 U586 ( .A(n516), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U587 ( .A(G120GAT), .B(KEYINPUT49), .Z(n518) );
  NAND2_X1 U588 ( .A1(n522), .A2(n557), .ZN(n517) );
  XNOR2_X1 U589 ( .A(n518), .B(n517), .ZN(G1341GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n520) );
  NAND2_X1 U591 ( .A1(n522), .A2(n560), .ZN(n519) );
  XNOR2_X1 U592 ( .A(n520), .B(n519), .ZN(n521) );
  XOR2_X1 U593 ( .A(G127GAT), .B(n521), .Z(G1342GAT) );
  XOR2_X1 U594 ( .A(G134GAT), .B(KEYINPUT51), .Z(n524) );
  NAND2_X1 U595 ( .A1(n522), .A2(n563), .ZN(n523) );
  XNOR2_X1 U596 ( .A(n524), .B(n523), .ZN(G1343GAT) );
  NAND2_X1 U597 ( .A1(n526), .A2(n525), .ZN(n537) );
  NOR2_X1 U598 ( .A1(n568), .A2(n537), .ZN(n527) );
  XOR2_X1 U599 ( .A(G141GAT), .B(n527), .Z(G1344GAT) );
  NOR2_X1 U600 ( .A1(n528), .A2(n537), .ZN(n533) );
  XOR2_X1 U601 ( .A(KEYINPUT53), .B(KEYINPUT118), .Z(n530) );
  XNOR2_X1 U602 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n529) );
  XNOR2_X1 U603 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U604 ( .A(KEYINPUT117), .B(n531), .ZN(n532) );
  XNOR2_X1 U605 ( .A(n533), .B(n532), .ZN(G1345GAT) );
  NOR2_X1 U606 ( .A1(n576), .A2(n537), .ZN(n535) );
  XNOR2_X1 U607 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n534) );
  XNOR2_X1 U608 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U609 ( .A(G155GAT), .B(n536), .ZN(G1346GAT) );
  NOR2_X1 U610 ( .A1(n538), .A2(n537), .ZN(n540) );
  XNOR2_X1 U611 ( .A(G162GAT), .B(KEYINPUT121), .ZN(n539) );
  XNOR2_X1 U612 ( .A(n540), .B(n539), .ZN(G1347GAT) );
  XNOR2_X1 U613 ( .A(KEYINPUT54), .B(n543), .ZN(n545) );
  NAND2_X1 U614 ( .A1(n545), .A2(n544), .ZN(n546) );
  NAND2_X1 U615 ( .A1(n547), .A2(n567), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n548), .B(KEYINPUT55), .ZN(n550) );
  AND2_X1 U617 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X2 U618 ( .A(KEYINPUT122), .B(n551), .ZN(n562) );
  NAND2_X1 U619 ( .A1(n562), .A2(n552), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n553), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT57), .B(KEYINPUT124), .Z(n555) );
  XNOR2_X1 U622 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U624 ( .A(KEYINPUT123), .B(n556), .Z(n559) );
  NAND2_X1 U625 ( .A1(n557), .A2(n562), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(G1349GAT) );
  NAND2_X1 U627 ( .A1(n562), .A2(n560), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n561), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U629 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n565) );
  NAND2_X1 U630 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(G1351GAT) );
  NAND2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n579) );
  NOR2_X1 U633 ( .A1(n568), .A2(n579), .ZN(n570) );
  XNOR2_X1 U634 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(n571), .ZN(G1352GAT) );
  NOR2_X1 U637 ( .A1(n572), .A2(n579), .ZN(n574) );
  XNOR2_X1 U638 ( .A(KEYINPUT125), .B(KEYINPUT61), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n575) );
  XOR2_X1 U640 ( .A(G204GAT), .B(n575), .Z(G1353GAT) );
  NOR2_X1 U641 ( .A1(n576), .A2(n579), .ZN(n577) );
  XOR2_X1 U642 ( .A(KEYINPUT126), .B(n577), .Z(n578) );
  XNOR2_X1 U643 ( .A(G211GAT), .B(n578), .ZN(G1354GAT) );
  NOR2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n582) );
  XNOR2_X1 U645 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

