//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 1 1 1 0 1 0 0 1 0 0 1 0 1 0 1 0 1 0 1 0 0 1 1 0 1 1 0 0 1 0 1 0 1 1 1 1 1 1 1 1 1 1 0 1 0 0 1 0 1 0 1 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:01 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n444, new_n445, new_n446, new_n451, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n460, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n570, new_n571, new_n572, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n632, new_n633, new_n636, new_n638, new_n639, new_n640,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n824, new_n825, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1184,
    new_n1185, new_n1186, new_n1187;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT66), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  XNOR2_X1  g015(.A(KEYINPUT67), .B(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  INV_X1    g018(.A(G2072), .ZN(new_n444));
  INV_X1    g019(.A(G2078), .ZN(new_n445));
  NOR2_X1   g020(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g021(.A1(new_n446), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g022(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g023(.A(KEYINPUT68), .B(G452), .Z(G391));
  AND2_X1   g024(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g025(.A1(G7), .A2(G661), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g027(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g028(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n455));
  XNOR2_X1  g030(.A(KEYINPUT69), .B(KEYINPUT2), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n455), .B(new_n456), .ZN(new_n457));
  NOR4_X1   g032(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT70), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n457), .A2(new_n460), .ZN(G325));
  INV_X1    g036(.A(G325), .ZN(G261));
  AOI22_X1  g037(.A1(new_n457), .A2(G2106), .B1(G567), .B2(new_n460), .ZN(G319));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT71), .ZN(new_n465));
  XNOR2_X1  g040(.A(new_n464), .B(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OR2_X1    g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g045(.A(G2105), .B1(new_n466), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT72), .ZN(new_n472));
  INV_X1    g047(.A(G2104), .ZN(new_n473));
  NOR3_X1   g048(.A1(new_n472), .A2(new_n473), .A3(G2105), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  AOI21_X1  g050(.A(KEYINPUT72), .B1(new_n475), .B2(G2104), .ZN(new_n476));
  OAI21_X1  g051(.A(G101), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  XNOR2_X1  g052(.A(KEYINPUT3), .B(G2104), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n478), .A2(G137), .A3(new_n475), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n471), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  AOI21_X1  g056(.A(new_n475), .B1(new_n468), .B2(new_n469), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  XOR2_X1   g058(.A(new_n483), .B(KEYINPUT73), .Z(new_n484));
  NAND2_X1  g059(.A1(new_n478), .A2(new_n475), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n475), .A2(G112), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n484), .B(new_n487), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  XOR2_X1   g065(.A(new_n490), .B(KEYINPUT74), .Z(G162));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT75), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n494), .A2(new_n495), .A3(G2105), .ZN(new_n496));
  OAI21_X1  g071(.A(KEYINPUT75), .B1(new_n475), .B2(G114), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n493), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  AND2_X1   g073(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n499));
  NOR2_X1   g074(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n500));
  OAI211_X1 g075(.A(G126), .B(G2105), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  OAI211_X1 g077(.A(G138), .B(new_n475), .C1(new_n499), .C2(new_n500), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT4), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n478), .A2(new_n505), .A3(G138), .A4(new_n475), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n502), .B1(new_n504), .B2(new_n506), .ZN(G164));
  NOR2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT76), .B(G651), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT6), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n512), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT77), .B(G88), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n512), .A2(G50), .A3(G543), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n517), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n522), .A2(new_n510), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n520), .A2(new_n521), .A3(new_n523), .ZN(G303));
  INV_X1    g099(.A(G303), .ZN(G166));
  NAND2_X1  g100(.A1(new_n518), .A2(G89), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n517), .A2(G63), .A3(G651), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT78), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n527), .B(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  AND3_X1   g106(.A1(new_n526), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n512), .A2(G543), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(KEYINPUT79), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT79), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n512), .A2(new_n535), .A3(G543), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G51), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n532), .A2(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  INV_X1    g115(.A(G52), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n541), .B1(new_n534), .B2(new_n536), .ZN(new_n542));
  NAND2_X1  g117(.A1(G77), .A2(G543), .ZN(new_n543));
  AND2_X1   g118(.A1(new_n515), .A2(new_n516), .ZN(new_n544));
  INV_X1    g119(.A(G64), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n510), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(G90), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n512), .A2(new_n517), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n542), .A2(new_n551), .ZN(G171));
  INV_X1    g127(.A(G43), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n553), .B1(new_n534), .B2(new_n536), .ZN(new_n554));
  NAND2_X1  g129(.A1(G68), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G56), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n544), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(new_n547), .ZN(new_n558));
  INV_X1    g133(.A(G81), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n559), .B2(new_n550), .ZN(new_n560));
  OAI21_X1  g135(.A(KEYINPUT80), .B1(new_n554), .B2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n536), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n535), .B1(new_n512), .B2(G543), .ZN(new_n563));
  OAI21_X1  g138(.A(G43), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT80), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n518), .A2(G81), .B1(new_n547), .B2(new_n557), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n561), .A2(new_n567), .A3(G860), .ZN(G153));
  NAND4_X1  g143(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(new_n572));
  XOR2_X1   g147(.A(new_n572), .B(KEYINPUT81), .Z(G188));
  INV_X1    g148(.A(G53), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT82), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n574), .B1(new_n575), .B2(KEYINPUT9), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n512), .A2(G543), .A3(new_n576), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n575), .A2(KEYINPUT9), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n578), .ZN(new_n580));
  NAND4_X1  g155(.A1(new_n512), .A2(G543), .A3(new_n580), .A4(new_n576), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n517), .A2(G65), .ZN(new_n582));
  NAND2_X1  g157(.A1(G78), .A2(G543), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(G651), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n512), .A2(G91), .A3(new_n517), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n579), .A2(new_n581), .A3(new_n585), .A4(new_n586), .ZN(G299));
  INV_X1    g162(.A(G171), .ZN(G301));
  NAND3_X1  g163(.A1(new_n512), .A2(G49), .A3(G543), .ZN(new_n589));
  OAI21_X1  g164(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n590));
  INV_X1    g165(.A(G87), .ZN(new_n591));
  OAI211_X1 g166(.A(new_n589), .B(new_n590), .C1(new_n550), .C2(new_n591), .ZN(G288));
  INV_X1    g167(.A(G651), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(KEYINPUT76), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT76), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(G651), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n511), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  OAI211_X1 g172(.A(G86), .B(new_n517), .C1(new_n597), .C2(new_n508), .ZN(new_n598));
  OAI211_X1 g173(.A(G48), .B(G543), .C1(new_n597), .C2(new_n508), .ZN(new_n599));
  INV_X1    g174(.A(G61), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n600), .B1(new_n515), .B2(new_n516), .ZN(new_n601));
  AND2_X1   g176(.A1(G73), .A2(G543), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n547), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n598), .A2(new_n599), .A3(new_n603), .ZN(G305));
  NAND2_X1  g179(.A1(new_n537), .A2(G47), .ZN(new_n605));
  INV_X1    g180(.A(G60), .ZN(new_n606));
  INV_X1    g181(.A(G72), .ZN(new_n607));
  OAI22_X1  g182(.A1(new_n544), .A2(new_n606), .B1(new_n607), .B2(new_n514), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n510), .B1(new_n608), .B2(KEYINPUT83), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT83), .ZN(new_n610));
  OAI221_X1 g185(.A(new_n610), .B1(new_n607), .B2(new_n514), .C1(new_n544), .C2(new_n606), .ZN(new_n611));
  XNOR2_X1  g186(.A(KEYINPUT84), .B(G85), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n609), .A2(new_n611), .B1(new_n518), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n605), .A2(new_n613), .ZN(G290));
  INV_X1    g189(.A(G868), .ZN(new_n615));
  NOR2_X1   g190(.A1(G301), .A2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT10), .ZN(new_n617));
  INV_X1    g192(.A(G92), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n550), .B2(new_n618), .ZN(new_n619));
  NAND4_X1  g194(.A1(new_n512), .A2(KEYINPUT10), .A3(G92), .A4(new_n517), .ZN(new_n620));
  NAND2_X1  g195(.A1(G79), .A2(G543), .ZN(new_n621));
  INV_X1    g196(.A(G66), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n544), .B2(new_n622), .ZN(new_n623));
  AOI22_X1  g198(.A1(new_n619), .A2(new_n620), .B1(G651), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n537), .A2(G54), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(KEYINPUT85), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n616), .B1(new_n629), .B2(new_n615), .ZN(G284));
  AOI21_X1  g205(.A(new_n616), .B1(new_n629), .B2(new_n615), .ZN(G321));
  NOR2_X1   g206(.A1(G286), .A2(new_n615), .ZN(new_n632));
  XOR2_X1   g207(.A(G299), .B(KEYINPUT86), .Z(new_n633));
  AOI21_X1  g208(.A(new_n632), .B1(new_n633), .B2(new_n615), .ZN(G297));
  AOI21_X1  g209(.A(new_n632), .B1(new_n633), .B2(new_n615), .ZN(G280));
  INV_X1    g210(.A(G559), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n629), .B1(new_n636), .B2(G860), .ZN(G148));
  NAND2_X1  g212(.A1(new_n561), .A2(new_n567), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(new_n615), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n628), .A2(G559), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n639), .B1(new_n640), .B2(new_n615), .ZN(G323));
  XNOR2_X1  g216(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g217(.A1(new_n474), .A2(new_n476), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n643), .A2(new_n478), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT12), .Z(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT13), .Z(new_n646));
  INV_X1    g221(.A(G2100), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n482), .A2(G123), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n475), .A2(G111), .ZN(new_n651));
  OAI21_X1  g226(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n652));
  INV_X1    g227(.A(G135), .ZN(new_n653));
  OAI221_X1 g228(.A(new_n650), .B1(new_n651), .B2(new_n652), .C1(new_n653), .C2(new_n485), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(G2096), .Z(new_n655));
  NAND3_X1  g230(.A1(new_n648), .A2(new_n649), .A3(new_n655), .ZN(G156));
  INV_X1    g231(.A(KEYINPUT14), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2427), .B(G2438), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2430), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT15), .B(G2435), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n657), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n661), .B1(new_n660), .B2(new_n659), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2451), .B(G2454), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT16), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1341), .B(G1348), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n662), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2443), .B(G2446), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(G14), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n667), .A2(new_n668), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(G401));
  XNOR2_X1  g247(.A(G2067), .B(G2678), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT87), .ZN(new_n674));
  XOR2_X1   g249(.A(G2084), .B(G2090), .Z(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G2072), .B(G2078), .Z(new_n677));
  NOR3_X1   g252(.A1(new_n674), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT88), .B(KEYINPUT18), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n677), .B(KEYINPUT17), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n681), .A2(new_n675), .A3(new_n674), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n675), .B1(new_n674), .B2(new_n677), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n683), .A2(KEYINPUT89), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(KEYINPUT89), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n685), .B1(new_n674), .B2(new_n681), .ZN(new_n686));
  OAI211_X1 g261(.A(new_n680), .B(new_n682), .C1(new_n684), .C2(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G2096), .B(G2100), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(G227));
  XNOR2_X1  g264(.A(G1971), .B(G1976), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT19), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(G1956), .B(G2474), .Z(new_n693));
  XOR2_X1   g268(.A(G1961), .B(G1966), .Z(new_n694));
  AND2_X1   g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT20), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n693), .A2(new_n694), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  MUX2_X1   g275(.A(new_n700), .B(new_n699), .S(new_n692), .Z(new_n701));
  NOR2_X1   g276(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1991), .B(G1996), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(G1981), .B(G1986), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(G229));
  INV_X1    g284(.A(G29), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G33), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT25), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n478), .A2(G127), .ZN(new_n714));
  NAND2_X1  g289(.A1(G115), .A2(G2104), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n475), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  AOI211_X1 g291(.A(new_n713), .B(new_n716), .C1(G139), .C2(new_n486), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT97), .Z(new_n718));
  OAI21_X1  g293(.A(new_n711), .B1(new_n718), .B2(new_n710), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(new_n444), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n710), .A2(G27), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G164), .B2(new_n710), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(new_n445), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n710), .A2(G26), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT28), .Z(new_n725));
  NAND2_X1  g300(.A1(new_n482), .A2(G128), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT96), .Z(new_n727));
  NAND2_X1  g302(.A1(new_n486), .A2(G140), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n475), .A2(G116), .ZN(new_n729));
  OAI21_X1  g304(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n727), .B(new_n728), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n725), .B1(new_n731), .B2(G29), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G2067), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n720), .A2(new_n723), .A3(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(G29), .A2(G35), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G162), .B2(G29), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT29), .B(G2090), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n710), .A2(G32), .ZN(new_n739));
  AOI22_X1  g314(.A1(new_n486), .A2(G141), .B1(G129), .B2(new_n482), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n643), .A2(G105), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT98), .B(KEYINPUT26), .Z(new_n742));
  NAND3_X1  g317(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n740), .A2(new_n741), .A3(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n739), .B1(new_n746), .B2(new_n710), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT27), .B(G1996), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n480), .A2(G29), .ZN(new_n750));
  INV_X1    g325(.A(G2084), .ZN(new_n751));
  INV_X1    g326(.A(G34), .ZN(new_n752));
  AND2_X1   g327(.A1(new_n752), .A2(KEYINPUT24), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n752), .A2(KEYINPUT24), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n710), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  AND3_X1   g330(.A1(new_n750), .A2(new_n751), .A3(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n751), .B1(new_n750), .B2(new_n755), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT31), .B(G11), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT30), .ZN(new_n759));
  AND2_X1   g334(.A1(new_n759), .A2(G28), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n710), .B1(new_n759), .B2(G28), .ZN(new_n761));
  OAI221_X1 g336(.A(new_n758), .B1(new_n760), .B2(new_n761), .C1(new_n654), .C2(new_n710), .ZN(new_n762));
  NOR3_X1   g337(.A1(new_n756), .A2(new_n757), .A3(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(G16), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(G5), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G171), .B2(new_n764), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n749), .B(new_n763), .C1(G1961), .C2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n764), .A2(G20), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT23), .Z(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G299), .B2(G16), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(G1956), .Z(new_n771));
  NOR4_X1   g346(.A1(new_n734), .A2(new_n738), .A3(new_n767), .A4(new_n771), .ZN(new_n772));
  MUX2_X1   g347(.A(G19), .B(new_n638), .S(G16), .Z(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G1341), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n764), .A2(G4), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(new_n629), .B2(new_n764), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n774), .B1(G1348), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n764), .A2(G21), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G168), .B2(new_n764), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G1966), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G1961), .B2(new_n766), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n776), .A2(G1348), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n772), .A2(new_n777), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n764), .A2(G24), .ZN(new_n784));
  INV_X1    g359(.A(G290), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n784), .B1(new_n785), .B2(new_n764), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT92), .B(G1986), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n786), .B(new_n787), .Z(new_n788));
  NAND2_X1  g363(.A1(new_n482), .A2(G119), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n475), .A2(G107), .ZN(new_n790));
  OAI21_X1  g365(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n791));
  INV_X1    g366(.A(G131), .ZN(new_n792));
  OAI221_X1 g367(.A(new_n789), .B1(new_n790), .B2(new_n791), .C1(new_n792), .C2(new_n485), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT90), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  MUX2_X1   g370(.A(G25), .B(new_n795), .S(G29), .Z(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT35), .B(G1991), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT91), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n796), .B(new_n798), .Z(new_n799));
  NAND2_X1  g374(.A1(new_n764), .A2(G22), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G166), .B2(new_n764), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G1971), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n764), .A2(G23), .ZN(new_n803));
  INV_X1    g378(.A(G288), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n803), .B1(new_n804), .B2(new_n764), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT33), .B(G1976), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT94), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n805), .B(new_n807), .Z(new_n808));
  MUX2_X1   g383(.A(G6), .B(G305), .S(G16), .Z(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT32), .B(G1981), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT93), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n809), .B(new_n811), .Z(new_n812));
  NOR3_X1   g387(.A1(new_n802), .A2(new_n808), .A3(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n788), .B(new_n799), .C1(new_n814), .C2(KEYINPUT34), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT95), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n814), .A2(KEYINPUT34), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(KEYINPUT36), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT36), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n817), .A2(new_n821), .A3(new_n818), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n783), .B1(new_n820), .B2(new_n822), .ZN(G311));
  INV_X1    g398(.A(new_n783), .ZN(new_n824));
  INV_X1    g399(.A(new_n822), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n821), .B1(new_n817), .B2(new_n818), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(G150));
  NAND2_X1  g402(.A1(G80), .A2(G543), .ZN(new_n828));
  INV_X1    g403(.A(G67), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n828), .B1(new_n544), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(new_n547), .ZN(new_n831));
  INV_X1    g406(.A(G93), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n831), .B1(new_n832), .B2(new_n550), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n833), .B1(new_n537), .B2(G55), .ZN(new_n834));
  INV_X1    g409(.A(G860), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT37), .ZN(new_n837));
  OAI21_X1  g412(.A(G55), .B1(new_n562), .B2(new_n563), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n518), .A2(G93), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n838), .A2(new_n831), .A3(new_n839), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n561), .A2(new_n567), .A3(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n834), .B1(new_n554), .B2(new_n560), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT99), .ZN(new_n843));
  AND3_X1   g418(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n843), .B1(new_n841), .B2(new_n842), .ZN(new_n845));
  OR3_X1    g420(.A1(new_n844), .A2(new_n845), .A3(KEYINPUT38), .ZN(new_n846));
  OAI21_X1  g421(.A(KEYINPUT38), .B1(new_n844), .B2(new_n845), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n629), .A2(G559), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n849), .ZN(new_n851));
  AND3_X1   g426(.A1(new_n850), .A2(KEYINPUT39), .A3(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT100), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n850), .A2(new_n851), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n835), .B1(new_n855), .B2(KEYINPUT39), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n837), .B1(new_n853), .B2(new_n856), .ZN(G145));
  XNOR2_X1  g432(.A(new_n654), .B(new_n480), .ZN(new_n858));
  XNOR2_X1  g433(.A(G162), .B(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n504), .A2(new_n506), .ZN(new_n861));
  AND2_X1   g436(.A1(new_n498), .A2(new_n501), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n731), .B(new_n863), .ZN(new_n864));
  AOI22_X1  g439(.A1(new_n486), .A2(G142), .B1(G130), .B2(new_n482), .ZN(new_n865));
  OAI21_X1  g440(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT101), .ZN(new_n867));
  INV_X1    g442(.A(G118), .ZN(new_n868));
  AOI22_X1  g443(.A1(new_n866), .A2(new_n867), .B1(new_n868), .B2(G2105), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n869), .B1(new_n867), .B2(new_n866), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n865), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n864), .B(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n795), .B(KEYINPUT102), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n645), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n718), .B(new_n746), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n874), .A2(new_n875), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n872), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n878), .ZN(new_n880));
  INV_X1    g455(.A(new_n872), .ZN(new_n881));
  NOR3_X1   g456(.A1(new_n880), .A2(new_n876), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n860), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n881), .B1(new_n880), .B2(new_n876), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n877), .A2(new_n878), .A3(new_n872), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n884), .A2(new_n885), .A3(new_n859), .ZN(new_n886));
  INV_X1    g461(.A(G37), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n883), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g464(.A1(new_n840), .A2(new_n615), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n841), .A2(new_n842), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(KEYINPUT99), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n640), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  OAI22_X1  g469(.A1(new_n844), .A2(new_n845), .B1(new_n628), .B2(G559), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n626), .A2(KEYINPUT103), .A3(G299), .ZN(new_n896));
  NAND2_X1  g471(.A1(G299), .A2(KEYINPUT103), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n585), .A2(new_n586), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT103), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n898), .A2(new_n899), .A3(new_n581), .A4(new_n579), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n897), .A2(new_n900), .A3(new_n625), .A4(new_n624), .ZN(new_n901));
  AND3_X1   g476(.A1(new_n896), .A2(new_n901), .A3(KEYINPUT41), .ZN(new_n902));
  AOI21_X1  g477(.A(KEYINPUT41), .B1(new_n896), .B2(new_n901), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n894), .A2(new_n895), .A3(new_n904), .ZN(new_n905));
  OR2_X1    g480(.A1(new_n905), .A2(KEYINPUT104), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(KEYINPUT104), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n896), .A2(new_n901), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n908), .B1(new_n894), .B2(new_n895), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n906), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(G290), .B(G288), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT105), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n785), .A2(new_n804), .ZN(new_n914));
  NAND2_X1  g489(.A1(G290), .A2(G288), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n914), .A2(KEYINPUT105), .A3(new_n915), .ZN(new_n916));
  XOR2_X1   g491(.A(G303), .B(G305), .Z(new_n917));
  NAND3_X1  g492(.A1(new_n913), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  OR3_X1    g493(.A1(new_n911), .A2(new_n917), .A3(new_n912), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  XOR2_X1   g495(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n921));
  XNOR2_X1  g496(.A(new_n920), .B(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n910), .A2(KEYINPUT107), .A3(new_n922), .ZN(new_n923));
  AND2_X1   g498(.A1(new_n918), .A2(new_n919), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(new_n921), .ZN(new_n925));
  INV_X1    g500(.A(new_n921), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n920), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n925), .A2(KEYINPUT107), .A3(new_n927), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n928), .B(new_n906), .C1(new_n909), .C2(new_n907), .ZN(new_n929));
  OR2_X1    g504(.A1(new_n922), .A2(KEYINPUT107), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n923), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n890), .B1(new_n931), .B2(new_n615), .ZN(G295));
  OAI21_X1  g507(.A(new_n890), .B1(new_n931), .B2(new_n615), .ZN(G331));
  NAND2_X1  g508(.A1(G286), .A2(G171), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n532), .B(new_n538), .C1(new_n542), .C2(new_n551), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(new_n844), .B2(new_n845), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n934), .A2(new_n935), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n892), .A2(new_n893), .A3(new_n938), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n937), .A2(new_n939), .A3(new_n904), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n908), .B1(new_n937), .B2(new_n939), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n920), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n937), .A2(new_n939), .ZN(new_n943));
  INV_X1    g518(.A(new_n908), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n937), .A2(new_n939), .A3(new_n904), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n945), .A2(new_n924), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n942), .A2(new_n947), .A3(new_n887), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(KEYINPUT43), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n946), .B1(new_n941), .B2(KEYINPUT108), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n943), .A2(KEYINPUT108), .A3(new_n944), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n920), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n940), .A2(new_n941), .ZN(new_n953));
  AOI21_X1  g528(.A(G37), .B1(new_n953), .B2(new_n924), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n949), .B1(new_n955), .B2(KEYINPUT43), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT44), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT109), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT43), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n954), .A2(new_n959), .A3(new_n960), .A4(new_n942), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n942), .A2(new_n947), .A3(new_n960), .A4(new_n887), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT109), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n955), .A2(KEYINPUT110), .A3(KEYINPUT43), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n960), .B1(new_n952), .B2(new_n954), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT44), .B1(new_n967), .B2(KEYINPUT110), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n958), .B1(new_n966), .B2(new_n968), .ZN(G397));
  INV_X1    g544(.A(G1384), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n863), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT45), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n471), .A2(G40), .A3(new_n477), .A4(new_n479), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G1996), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  XOR2_X1   g552(.A(new_n977), .B(KEYINPUT111), .Z(new_n978));
  XOR2_X1   g553(.A(new_n975), .B(KEYINPUT112), .Z(new_n979));
  INV_X1    g554(.A(G2067), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n731), .B(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n981), .B1(new_n976), .B2(new_n746), .ZN(new_n982));
  AOI22_X1  g557(.A1(new_n978), .A2(new_n746), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n795), .A2(new_n798), .ZN(new_n984));
  AND2_X1   g559(.A1(new_n795), .A2(new_n798), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n979), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n983), .A2(new_n986), .ZN(new_n987));
  AND2_X1   g562(.A1(G290), .A2(G1986), .ZN(new_n988));
  NOR2_X1   g563(.A1(G290), .A2(G1986), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n975), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT113), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n991), .B(new_n992), .ZN(new_n993));
  OAI21_X1  g568(.A(KEYINPUT116), .B1(G164), .B2(G1384), .ZN(new_n994));
  INV_X1    g569(.A(new_n974), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT116), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n863), .A2(new_n996), .A3(new_n970), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n994), .A2(new_n995), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n804), .A2(G1976), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n998), .A2(G8), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(KEYINPUT52), .ZN(new_n1001));
  INV_X1    g576(.A(G1976), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT52), .B1(G288), .B2(new_n1002), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n998), .A2(G8), .A3(new_n999), .A4(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT49), .ZN(new_n1005));
  INV_X1    g580(.A(G1981), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1006), .B1(new_n603), .B2(KEYINPUT117), .ZN(new_n1007));
  AND2_X1   g582(.A1(G305), .A2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(G305), .A2(new_n1007), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1005), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  OR2_X1    g585(.A1(G305), .A2(new_n1007), .ZN(new_n1011));
  NAND2_X1  g586(.A1(G305), .A2(new_n1007), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1011), .A2(KEYINPUT49), .A3(new_n1012), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1010), .A2(new_n1013), .A3(G8), .A4(new_n998), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1001), .A2(new_n1004), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT118), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1001), .A2(new_n1014), .A3(KEYINPUT118), .A4(new_n1004), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  XOR2_X1   g594(.A(KEYINPUT114), .B(G1971), .Z(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n863), .A2(KEYINPUT45), .A3(new_n970), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(new_n995), .ZN(new_n1023));
  AOI21_X1  g598(.A(G1384), .B1(new_n861), .B2(new_n862), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1024), .A2(KEYINPUT45), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1021), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(KEYINPUT115), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n974), .B1(new_n1024), .B2(KEYINPUT45), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n973), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT115), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1029), .A2(new_n1030), .A3(new_n1021), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT50), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n994), .A2(new_n1032), .A3(new_n997), .ZN(new_n1033));
  INV_X1    g608(.A(G2090), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n974), .B1(new_n971), .B2(KEYINPUT50), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1027), .A2(new_n1031), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(G303), .A2(G8), .ZN(new_n1038));
  XOR2_X1   g613(.A(new_n1038), .B(KEYINPUT55), .Z(new_n1039));
  NAND3_X1  g614(.A1(new_n1037), .A2(new_n1039), .A3(G8), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1039), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n995), .B1(new_n971), .B2(KEYINPUT50), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n994), .A2(new_n997), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1042), .B1(KEYINPUT50), .B2(new_n1043), .ZN(new_n1044));
  AOI22_X1  g619(.A1(new_n1044), .A2(new_n1034), .B1(new_n1029), .B2(new_n1021), .ZN(new_n1045));
  INV_X1    g620(.A(G8), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1041), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1048));
  INV_X1    g623(.A(G1961), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1024), .A2(new_n996), .ZN(new_n1051));
  AOI211_X1 g626(.A(KEYINPUT116), .B(G1384), .C1(new_n861), .C2(new_n862), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n972), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1053), .A2(KEYINPUT53), .A3(new_n445), .A4(new_n1028), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1028), .A2(new_n973), .A3(new_n445), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1050), .A2(new_n1054), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n542), .ZN(new_n1059));
  INV_X1    g634(.A(new_n551), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1059), .A2(KEYINPUT54), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1062), .B1(new_n542), .B2(new_n551), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1029), .A2(G2078), .ZN(new_n1066));
  AOI22_X1  g641(.A1(new_n1066), .A2(KEYINPUT53), .B1(new_n1063), .B2(new_n1061), .ZN(new_n1067));
  AOI22_X1  g642(.A1(new_n1048), .A2(new_n1049), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1068));
  AOI22_X1  g643(.A1(new_n1058), .A2(new_n1065), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  AND4_X1   g644(.A1(new_n1019), .A2(new_n1040), .A3(new_n1047), .A4(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT125), .ZN(new_n1071));
  AOI21_X1  g646(.A(G1966), .B1(new_n1053), .B2(new_n1028), .ZN(new_n1072));
  AND3_X1   g647(.A1(new_n1033), .A2(new_n751), .A3(new_n1035), .ZN(new_n1073));
  OAI21_X1  g648(.A(G8), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n538), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n526), .A2(new_n529), .A3(new_n531), .ZN(new_n1076));
  OAI21_X1  g651(.A(G8), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1046), .B1(new_n532), .B2(new_n538), .ZN(new_n1078));
  OAI21_X1  g653(.A(KEYINPUT51), .B1(new_n1078), .B2(KEYINPUT124), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1074), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT51), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT124), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1081), .B1(new_n1077), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(G1966), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT45), .B1(new_n994), .B2(new_n997), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1084), .B1(new_n1085), .B2(new_n1023), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1033), .A2(new_n751), .A3(new_n1035), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  OAI211_X1 g663(.A(G8), .B(new_n1083), .C1(new_n1088), .C2(G286), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1080), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1077), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1071), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  AOI211_X1 g668(.A(KEYINPUT125), .B(new_n1091), .C1(new_n1080), .C2(new_n1089), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1070), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(KEYINPUT126), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT126), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1070), .B(new_n1097), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1044), .A2(G1956), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1029), .ZN(new_n1101));
  XNOR2_X1  g676(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n1102));
  XNOR2_X1  g677(.A(new_n1102), .B(G2072), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(G299), .A2(KEYINPUT120), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n1105), .B(KEYINPUT57), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1100), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1106), .B1(new_n1100), .B2(new_n1104), .ZN(new_n1108));
  INV_X1    g683(.A(G1348), .ZN(new_n1109));
  INV_X1    g684(.A(new_n998), .ZN(new_n1110));
  AOI22_X1  g685(.A1(new_n1109), .A2(new_n1048), .B1(new_n1110), .B2(new_n980), .ZN(new_n1111));
  OAI22_X1  g686(.A1(new_n1108), .A2(KEYINPUT122), .B1(new_n626), .B2(new_n1111), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1108), .A2(KEYINPUT122), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1107), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  XOR2_X1   g689(.A(KEYINPUT58), .B(G1341), .Z(new_n1115));
  AOI22_X1  g690(.A1(new_n1101), .A2(new_n976), .B1(new_n998), .B2(new_n1115), .ZN(new_n1116));
  OR3_X1    g691(.A1(new_n1116), .A2(KEYINPUT59), .A3(new_n638), .ZN(new_n1117));
  OAI21_X1  g692(.A(KEYINPUT59), .B1(new_n1116), .B2(new_n638), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n626), .A2(KEYINPUT60), .ZN(new_n1119));
  AOI22_X1  g694(.A1(new_n1117), .A2(new_n1118), .B1(new_n1111), .B2(new_n1119), .ZN(new_n1120));
  OR2_X1    g695(.A1(new_n1107), .A2(KEYINPUT61), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT60), .ZN(new_n1122));
  XOR2_X1   g697(.A(new_n1111), .B(new_n626), .Z(new_n1123));
  OAI211_X1 g698(.A(new_n1120), .B(new_n1121), .C1(new_n1122), .C2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1107), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1106), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1104), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1126), .B1(new_n1127), .B2(new_n1099), .ZN(new_n1128));
  OR2_X1    g703(.A1(new_n1128), .A2(KEYINPUT123), .ZN(new_n1129));
  AOI21_X1  g704(.A(KEYINPUT61), .B1(new_n1128), .B2(KEYINPUT123), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1125), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1114), .B1(new_n1124), .B2(new_n1131), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1096), .A2(new_n1098), .A3(new_n1132), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1014), .A2(new_n1002), .A3(new_n804), .ZN(new_n1134));
  NOR2_X1   g709(.A1(G305), .A2(G1981), .ZN(new_n1135));
  OAI211_X1 g710(.A(G8), .B(new_n998), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1136), .B1(new_n1015), .B2(new_n1040), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT119), .ZN(new_n1138));
  AND3_X1   g713(.A1(new_n1037), .A2(G8), .A3(new_n1039), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1039), .B1(new_n1037), .B2(G8), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1088), .A2(G8), .A3(G168), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1001), .A2(new_n1014), .A3(KEYINPUT63), .A4(new_n1004), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1138), .B1(new_n1141), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1037), .A2(G8), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(new_n1041), .ZN(new_n1147));
  AND4_X1   g722(.A1(new_n1138), .A2(new_n1144), .A3(new_n1147), .A4(new_n1040), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1145), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT63), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1019), .A2(new_n1040), .A3(new_n1047), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1150), .B1(new_n1151), .B2(new_n1142), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1137), .B1(new_n1149), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(KEYINPUT62), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1079), .B1(new_n1074), .B2(new_n1077), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1046), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1156));
  NOR3_X1   g731(.A1(new_n1156), .A2(new_n1083), .A3(new_n1078), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1092), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(KEYINPUT125), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT62), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1090), .A2(new_n1071), .A3(new_n1092), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1058), .A2(G171), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1151), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1154), .A2(new_n1162), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1153), .A2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n993), .B1(new_n1133), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(new_n981), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n979), .B1(new_n1168), .B2(new_n745), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT46), .ZN(new_n1170));
  AND2_X1   g745(.A1(new_n978), .A2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n978), .A2(new_n1170), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1169), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n1173), .B(KEYINPUT47), .ZN(new_n1174));
  AND2_X1   g749(.A1(new_n983), .A2(new_n984), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n731), .A2(G2067), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n979), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n989), .A2(new_n975), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1178), .B(KEYINPUT48), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n987), .A2(new_n1179), .ZN(new_n1180));
  AND3_X1   g755(.A1(new_n1174), .A2(new_n1177), .A3(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1167), .A2(new_n1181), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g757(.A(G319), .B1(new_n670), .B2(new_n671), .ZN(new_n1184));
  NOR2_X1   g758(.A1(new_n1184), .A2(G227), .ZN(new_n1185));
  NAND2_X1  g759(.A1(new_n708), .A2(new_n1185), .ZN(new_n1186));
  XNOR2_X1  g760(.A(new_n1186), .B(KEYINPUT127), .ZN(new_n1187));
  AND3_X1   g761(.A1(new_n1187), .A2(new_n888), .A3(new_n956), .ZN(G308));
  NAND3_X1  g762(.A1(new_n1187), .A2(new_n888), .A3(new_n956), .ZN(G225));
endmodule


