

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591;

  NAND2_X1 U322 ( .A1(n393), .A2(n392), .ZN(n487) );
  XNOR2_X1 U323 ( .A(n336), .B(n335), .ZN(n344) );
  XOR2_X1 U324 ( .A(KEYINPUT91), .B(n388), .Z(n520) );
  AND2_X1 U325 ( .A1(G228GAT), .A2(G233GAT), .ZN(n290) );
  XOR2_X1 U326 ( .A(n333), .B(n332), .Z(n291) );
  OR2_X1 U327 ( .A1(n480), .A2(n573), .ZN(n454) );
  XNOR2_X1 U328 ( .A(n441), .B(n290), .ZN(n327) );
  INV_X1 U329 ( .A(KEYINPUT112), .ZN(n469) );
  XNOR2_X1 U330 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U331 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U332 ( .A(n469), .B(KEYINPUT48), .ZN(n470) );
  XNOR2_X1 U333 ( .A(n334), .B(n291), .ZN(n335) );
  XNOR2_X1 U334 ( .A(n433), .B(n432), .ZN(n437) );
  XNOR2_X1 U335 ( .A(n471), .B(n470), .ZN(n532) );
  NOR2_X1 U336 ( .A1(n588), .A2(n411), .ZN(n412) );
  XNOR2_X1 U337 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U338 ( .A(KEYINPUT26), .B(n363), .ZN(n571) );
  XNOR2_X1 U339 ( .A(n445), .B(n444), .ZN(n579) );
  INV_X1 U340 ( .A(G43GAT), .ZN(n448) );
  XNOR2_X1 U341 ( .A(n447), .B(n446), .ZN(n506) );
  XNOR2_X1 U342 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U343 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U344 ( .A(n484), .B(n483), .ZN(G1349GAT) );
  XNOR2_X1 U345 ( .A(n451), .B(n450), .ZN(G1330GAT) );
  XOR2_X1 U346 ( .A(G176GAT), .B(KEYINPUT79), .Z(n293) );
  XNOR2_X1 U347 ( .A(G71GAT), .B(KEYINPUT20), .ZN(n292) );
  XNOR2_X1 U348 ( .A(n293), .B(n292), .ZN(n310) );
  XOR2_X1 U349 ( .A(G120GAT), .B(G127GAT), .Z(n295) );
  XNOR2_X1 U350 ( .A(G134GAT), .B(G99GAT), .ZN(n294) );
  XNOR2_X1 U351 ( .A(n295), .B(n294), .ZN(n297) );
  XOR2_X1 U352 ( .A(G43GAT), .B(G190GAT), .Z(n296) );
  XNOR2_X1 U353 ( .A(n297), .B(n296), .ZN(n306) );
  XNOR2_X1 U354 ( .A(G183GAT), .B(KEYINPUT78), .ZN(n298) );
  XNOR2_X1 U355 ( .A(n298), .B(KEYINPUT77), .ZN(n300) );
  XNOR2_X1 U356 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n299) );
  XNOR2_X1 U357 ( .A(n299), .B(KEYINPUT76), .ZN(n384) );
  XOR2_X1 U358 ( .A(n300), .B(n384), .Z(n304) );
  XOR2_X1 U359 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n302) );
  XNOR2_X1 U360 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n301) );
  XNOR2_X1 U361 ( .A(n302), .B(n301), .ZN(n353) );
  XNOR2_X1 U362 ( .A(G15GAT), .B(n353), .ZN(n303) );
  XNOR2_X1 U363 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U364 ( .A(n306), .B(n305), .ZN(n308) );
  NAND2_X1 U365 ( .A1(G227GAT), .A2(G233GAT), .ZN(n307) );
  XNOR2_X1 U366 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U367 ( .A(n310), .B(n309), .ZN(n361) );
  INV_X1 U368 ( .A(n361), .ZN(n535) );
  INV_X1 U369 ( .A(KEYINPUT38), .ZN(n447) );
  XOR2_X1 U370 ( .A(KEYINPUT73), .B(KEYINPUT11), .Z(n312) );
  NAND2_X1 U371 ( .A1(G232GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U372 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U373 ( .A(n313), .B(KEYINPUT9), .Z(n318) );
  XOR2_X1 U374 ( .A(G43GAT), .B(G50GAT), .Z(n315) );
  XNOR2_X1 U375 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n314) );
  XNOR2_X1 U376 ( .A(n315), .B(n314), .ZN(n422) );
  XNOR2_X1 U377 ( .A(G36GAT), .B(G190GAT), .ZN(n316) );
  XNOR2_X1 U378 ( .A(n316), .B(G218GAT), .ZN(n345) );
  XNOR2_X1 U379 ( .A(n422), .B(n345), .ZN(n317) );
  XNOR2_X1 U380 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U381 ( .A(KEYINPUT10), .B(G92GAT), .Z(n320) );
  XNOR2_X1 U382 ( .A(G162GAT), .B(G106GAT), .ZN(n319) );
  XNOR2_X1 U383 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U384 ( .A(n322), .B(n321), .Z(n324) );
  XOR2_X1 U385 ( .A(G29GAT), .B(G134GAT), .Z(n378) );
  XOR2_X1 U386 ( .A(G99GAT), .B(G85GAT), .Z(n440) );
  XNOR2_X1 U387 ( .A(n378), .B(n440), .ZN(n323) );
  XOR2_X1 U388 ( .A(n324), .B(n323), .Z(n557) );
  XNOR2_X1 U389 ( .A(KEYINPUT36), .B(n557), .ZN(n588) );
  XOR2_X1 U390 ( .A(KEYINPUT82), .B(G218GAT), .Z(n326) );
  XNOR2_X1 U391 ( .A(G50GAT), .B(G22GAT), .ZN(n325) );
  XNOR2_X1 U392 ( .A(n326), .B(n325), .ZN(n328) );
  XOR2_X1 U393 ( .A(G106GAT), .B(G78GAT), .Z(n441) );
  XOR2_X1 U394 ( .A(n329), .B(G155GAT), .Z(n336) );
  XOR2_X1 U395 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n331) );
  XNOR2_X1 U396 ( .A(G141GAT), .B(G162GAT), .ZN(n330) );
  XNOR2_X1 U397 ( .A(n331), .B(n330), .ZN(n383) );
  XNOR2_X1 U398 ( .A(n383), .B(KEYINPUT81), .ZN(n334) );
  XOR2_X1 U399 ( .A(KEYINPUT24), .B(KEYINPUT85), .Z(n333) );
  XNOR2_X1 U400 ( .A(G148GAT), .B(KEYINPUT86), .ZN(n332) );
  XOR2_X1 U401 ( .A(KEYINPUT84), .B(KEYINPUT83), .Z(n338) );
  XNOR2_X1 U402 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n337) );
  XNOR2_X1 U403 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U404 ( .A(G197GAT), .B(n339), .ZN(n356) );
  XOR2_X1 U405 ( .A(KEYINPUT22), .B(G204GAT), .Z(n341) );
  XNOR2_X1 U406 ( .A(KEYINPUT80), .B(KEYINPUT23), .ZN(n340) );
  XNOR2_X1 U407 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U408 ( .A(n356), .B(n342), .Z(n343) );
  XNOR2_X1 U409 ( .A(n344), .B(n343), .ZN(n476) );
  XOR2_X1 U410 ( .A(n345), .B(KEYINPUT92), .Z(n347) );
  NAND2_X1 U411 ( .A1(G226GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U412 ( .A(n347), .B(n346), .ZN(n350) );
  XOR2_X1 U413 ( .A(G8GAT), .B(G183GAT), .Z(n397) );
  XNOR2_X1 U414 ( .A(n397), .B(KEYINPUT94), .ZN(n348) );
  XNOR2_X1 U415 ( .A(n348), .B(KEYINPUT93), .ZN(n349) );
  XOR2_X1 U416 ( .A(n350), .B(n349), .Z(n355) );
  XOR2_X1 U417 ( .A(G64GAT), .B(G92GAT), .Z(n352) );
  XNOR2_X1 U418 ( .A(G176GAT), .B(G204GAT), .ZN(n351) );
  XNOR2_X1 U419 ( .A(n352), .B(n351), .ZN(n433) );
  XNOR2_X1 U420 ( .A(n353), .B(n433), .ZN(n354) );
  XNOR2_X1 U421 ( .A(n355), .B(n354), .ZN(n358) );
  INV_X1 U422 ( .A(n356), .ZN(n357) );
  XOR2_X1 U423 ( .A(n358), .B(n357), .Z(n364) );
  NAND2_X1 U424 ( .A1(n364), .A2(n361), .ZN(n359) );
  NAND2_X1 U425 ( .A1(n476), .A2(n359), .ZN(n360) );
  XOR2_X1 U426 ( .A(KEYINPUT25), .B(n360), .Z(n366) );
  NOR2_X1 U427 ( .A1(n476), .A2(n361), .ZN(n362) );
  XOR2_X1 U428 ( .A(KEYINPUT95), .B(n362), .Z(n363) );
  INV_X1 U429 ( .A(n364), .ZN(n523) );
  XOR2_X1 U430 ( .A(n523), .B(KEYINPUT27), .Z(n389) );
  NAND2_X1 U431 ( .A1(n571), .A2(n389), .ZN(n365) );
  NAND2_X1 U432 ( .A1(n366), .A2(n365), .ZN(n367) );
  XNOR2_X1 U433 ( .A(KEYINPUT96), .B(n367), .ZN(n387) );
  XOR2_X1 U434 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n369) );
  NAND2_X1 U435 ( .A1(G225GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U436 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U437 ( .A(n370), .B(KEYINPUT88), .Z(n374) );
  XNOR2_X1 U438 ( .A(G120GAT), .B(G148GAT), .ZN(n371) );
  XNOR2_X1 U439 ( .A(n371), .B(G57GAT), .ZN(n439) );
  XNOR2_X1 U440 ( .A(G1GAT), .B(G127GAT), .ZN(n372) );
  XNOR2_X1 U441 ( .A(n372), .B(G155GAT), .ZN(n396) );
  XNOR2_X1 U442 ( .A(n439), .B(n396), .ZN(n373) );
  XNOR2_X1 U443 ( .A(n374), .B(n373), .ZN(n382) );
  XOR2_X1 U444 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n376) );
  XNOR2_X1 U445 ( .A(KEYINPUT89), .B(KEYINPUT90), .ZN(n375) );
  XNOR2_X1 U446 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U447 ( .A(n377), .B(KEYINPUT87), .Z(n380) );
  XNOR2_X1 U448 ( .A(n378), .B(G85GAT), .ZN(n379) );
  XNOR2_X1 U449 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U450 ( .A(n382), .B(n381), .Z(n386) );
  XNOR2_X1 U451 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U452 ( .A(n386), .B(n385), .ZN(n388) );
  NAND2_X1 U453 ( .A1(n387), .A2(n388), .ZN(n393) );
  XNOR2_X1 U454 ( .A(n476), .B(KEYINPUT28), .ZN(n533) );
  AND2_X1 U455 ( .A1(n533), .A2(n535), .ZN(n391) );
  INV_X1 U456 ( .A(n389), .ZN(n390) );
  NOR2_X1 U457 ( .A1(n520), .A2(n390), .ZN(n530) );
  NAND2_X1 U458 ( .A1(n391), .A2(n530), .ZN(n392) );
  XOR2_X1 U459 ( .A(G64GAT), .B(G57GAT), .Z(n395) );
  XNOR2_X1 U460 ( .A(G211GAT), .B(G78GAT), .ZN(n394) );
  XNOR2_X1 U461 ( .A(n395), .B(n394), .ZN(n409) );
  XOR2_X1 U462 ( .A(n397), .B(n396), .Z(n399) );
  NAND2_X1 U463 ( .A1(G231GAT), .A2(G233GAT), .ZN(n398) );
  XNOR2_X1 U464 ( .A(n399), .B(n398), .ZN(n403) );
  XOR2_X1 U465 ( .A(KEYINPUT12), .B(KEYINPUT74), .Z(n401) );
  XNOR2_X1 U466 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n400) );
  XNOR2_X1 U467 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U468 ( .A(n403), .B(n402), .Z(n407) );
  XNOR2_X1 U469 ( .A(G22GAT), .B(G15GAT), .ZN(n404) );
  XNOR2_X1 U470 ( .A(n404), .B(KEYINPUT68), .ZN(n420) );
  XNOR2_X1 U471 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n405) );
  XNOR2_X1 U472 ( .A(n405), .B(KEYINPUT70), .ZN(n438) );
  XNOR2_X1 U473 ( .A(n420), .B(n438), .ZN(n406) );
  XNOR2_X1 U474 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U475 ( .A(n409), .B(n408), .Z(n584) );
  NAND2_X1 U476 ( .A1(n487), .A2(n584), .ZN(n410) );
  XOR2_X1 U477 ( .A(KEYINPUT101), .B(n410), .Z(n411) );
  XNOR2_X1 U478 ( .A(KEYINPUT37), .B(n412), .ZN(n519) );
  XOR2_X1 U479 ( .A(G1GAT), .B(G8GAT), .Z(n414) );
  XNOR2_X1 U480 ( .A(G169GAT), .B(G113GAT), .ZN(n413) );
  XNOR2_X1 U481 ( .A(n414), .B(n413), .ZN(n418) );
  XOR2_X1 U482 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n416) );
  XNOR2_X1 U483 ( .A(KEYINPUT69), .B(KEYINPUT66), .ZN(n415) );
  XNOR2_X1 U484 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U485 ( .A(n418), .B(n417), .ZN(n429) );
  XNOR2_X1 U486 ( .A(G197GAT), .B(G36GAT), .ZN(n419) );
  XNOR2_X1 U487 ( .A(n419), .B(G29GAT), .ZN(n421) );
  XOR2_X1 U488 ( .A(n421), .B(n420), .Z(n427) );
  XOR2_X1 U489 ( .A(n422), .B(KEYINPUT67), .Z(n424) );
  NAND2_X1 U490 ( .A1(G229GAT), .A2(G233GAT), .ZN(n423) );
  XNOR2_X1 U491 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U492 ( .A(n425), .B(G141GAT), .ZN(n426) );
  XNOR2_X1 U493 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U494 ( .A(n429), .B(n428), .Z(n573) );
  INV_X1 U495 ( .A(n573), .ZN(n559) );
  NAND2_X1 U496 ( .A1(G230GAT), .A2(G233GAT), .ZN(n431) );
  INV_X1 U497 ( .A(KEYINPUT33), .ZN(n430) );
  XOR2_X1 U498 ( .A(KEYINPUT31), .B(KEYINPUT72), .Z(n435) );
  XNOR2_X1 U499 ( .A(KEYINPUT32), .B(KEYINPUT71), .ZN(n434) );
  XNOR2_X1 U500 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U501 ( .A(n437), .B(n436), .ZN(n445) );
  XOR2_X1 U502 ( .A(n439), .B(n438), .Z(n443) );
  XNOR2_X1 U503 ( .A(n441), .B(n440), .ZN(n442) );
  NAND2_X1 U504 ( .A1(n559), .A2(n579), .ZN(n489) );
  NOR2_X1 U505 ( .A1(n519), .A2(n489), .ZN(n446) );
  NOR2_X1 U506 ( .A1(n535), .A2(n506), .ZN(n451) );
  XNOR2_X1 U507 ( .A(KEYINPUT104), .B(KEYINPUT40), .ZN(n449) );
  XNOR2_X1 U508 ( .A(n579), .B(KEYINPUT64), .ZN(n453) );
  INV_X1 U509 ( .A(KEYINPUT41), .ZN(n452) );
  XNOR2_X1 U510 ( .A(n453), .B(n452), .ZN(n480) );
  XNOR2_X1 U511 ( .A(n454), .B(KEYINPUT110), .ZN(n457) );
  INV_X1 U512 ( .A(n457), .ZN(n456) );
  INV_X1 U513 ( .A(KEYINPUT46), .ZN(n455) );
  NAND2_X1 U514 ( .A1(n456), .A2(n455), .ZN(n459) );
  NAND2_X1 U515 ( .A1(n457), .A2(KEYINPUT46), .ZN(n458) );
  NAND2_X1 U516 ( .A1(n459), .A2(n458), .ZN(n461) );
  XOR2_X1 U517 ( .A(KEYINPUT109), .B(n584), .Z(n563) );
  AND2_X1 U518 ( .A1(n563), .A2(n557), .ZN(n460) );
  AND2_X1 U519 ( .A1(n461), .A2(n460), .ZN(n462) );
  XNOR2_X1 U520 ( .A(n462), .B(KEYINPUT47), .ZN(n468) );
  NOR2_X1 U521 ( .A1(n588), .A2(n584), .ZN(n463) );
  XNOR2_X1 U522 ( .A(KEYINPUT45), .B(n463), .ZN(n464) );
  NAND2_X1 U523 ( .A1(n464), .A2(n579), .ZN(n465) );
  XNOR2_X1 U524 ( .A(n465), .B(KEYINPUT111), .ZN(n466) );
  NAND2_X1 U525 ( .A1(n466), .A2(n573), .ZN(n467) );
  NAND2_X1 U526 ( .A1(n468), .A2(n467), .ZN(n471) );
  XOR2_X1 U527 ( .A(n523), .B(KEYINPUT117), .Z(n472) );
  NOR2_X1 U528 ( .A1(n532), .A2(n472), .ZN(n473) );
  XNOR2_X1 U529 ( .A(n473), .B(KEYINPUT54), .ZN(n474) );
  NAND2_X1 U530 ( .A1(n474), .A2(n520), .ZN(n475) );
  XNOR2_X1 U531 ( .A(n475), .B(KEYINPUT65), .ZN(n572) );
  NAND2_X1 U532 ( .A1(n572), .A2(n476), .ZN(n478) );
  INV_X1 U533 ( .A(KEYINPUT55), .ZN(n477) );
  XNOR2_X1 U534 ( .A(n478), .B(n477), .ZN(n479) );
  NOR2_X1 U535 ( .A1(n535), .A2(n479), .ZN(n566) );
  INV_X1 U536 ( .A(n480), .ZN(n538) );
  NAND2_X1 U537 ( .A1(n566), .A2(n538), .ZN(n484) );
  XOR2_X1 U538 ( .A(KEYINPUT57), .B(KEYINPUT119), .Z(n482) );
  XOR2_X1 U539 ( .A(G176GAT), .B(KEYINPUT56), .Z(n481) );
  INV_X1 U540 ( .A(n557), .ZN(n565) );
  OR2_X1 U541 ( .A1(n584), .A2(n565), .ZN(n485) );
  XNOR2_X1 U542 ( .A(n485), .B(KEYINPUT16), .ZN(n486) );
  XNOR2_X1 U543 ( .A(n486), .B(KEYINPUT75), .ZN(n488) );
  NAND2_X1 U544 ( .A1(n488), .A2(n487), .ZN(n508) );
  OR2_X1 U545 ( .A1(n489), .A2(n508), .ZN(n498) );
  NOR2_X1 U546 ( .A1(n520), .A2(n498), .ZN(n491) );
  XNOR2_X1 U547 ( .A(KEYINPUT34), .B(KEYINPUT97), .ZN(n490) );
  XNOR2_X1 U548 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U549 ( .A(G1GAT), .B(n492), .ZN(G1324GAT) );
  NOR2_X1 U550 ( .A1(n523), .A2(n498), .ZN(n493) );
  XOR2_X1 U551 ( .A(G8GAT), .B(n493), .Z(G1325GAT) );
  NOR2_X1 U552 ( .A1(n498), .A2(n535), .ZN(n497) );
  XOR2_X1 U553 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n495) );
  XNOR2_X1 U554 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n494) );
  XNOR2_X1 U555 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U556 ( .A(n497), .B(n496), .ZN(G1326GAT) );
  NOR2_X1 U557 ( .A1(n533), .A2(n498), .ZN(n499) );
  XOR2_X1 U558 ( .A(G22GAT), .B(n499), .Z(G1327GAT) );
  XOR2_X1 U559 ( .A(KEYINPUT102), .B(KEYINPUT39), .Z(n501) );
  XNOR2_X1 U560 ( .A(G29GAT), .B(KEYINPUT100), .ZN(n500) );
  XNOR2_X1 U561 ( .A(n501), .B(n500), .ZN(n503) );
  NOR2_X1 U562 ( .A1(n520), .A2(n506), .ZN(n502) );
  XOR2_X1 U563 ( .A(n503), .B(n502), .Z(G1328GAT) );
  NOR2_X1 U564 ( .A1(n506), .A2(n523), .ZN(n505) );
  XNOR2_X1 U565 ( .A(G36GAT), .B(KEYINPUT103), .ZN(n504) );
  XNOR2_X1 U566 ( .A(n505), .B(n504), .ZN(G1329GAT) );
  NOR2_X1 U567 ( .A1(n506), .A2(n533), .ZN(n507) );
  XOR2_X1 U568 ( .A(G50GAT), .B(n507), .Z(G1331GAT) );
  NAND2_X1 U569 ( .A1(n538), .A2(n573), .ZN(n518) );
  OR2_X1 U570 ( .A1(n518), .A2(n508), .ZN(n515) );
  NOR2_X1 U571 ( .A1(n520), .A2(n515), .ZN(n510) );
  XNOR2_X1 U572 ( .A(KEYINPUT105), .B(KEYINPUT42), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U574 ( .A(G57GAT), .B(n511), .ZN(G1332GAT) );
  NOR2_X1 U575 ( .A1(n523), .A2(n515), .ZN(n512) );
  XOR2_X1 U576 ( .A(KEYINPUT106), .B(n512), .Z(n513) );
  XNOR2_X1 U577 ( .A(G64GAT), .B(n513), .ZN(G1333GAT) );
  NOR2_X1 U578 ( .A1(n535), .A2(n515), .ZN(n514) );
  XOR2_X1 U579 ( .A(G71GAT), .B(n514), .Z(G1334GAT) );
  NOR2_X1 U580 ( .A1(n533), .A2(n515), .ZN(n517) );
  XNOR2_X1 U581 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n517), .B(n516), .ZN(G1335GAT) );
  OR2_X1 U583 ( .A1(n519), .A2(n518), .ZN(n526) );
  NOR2_X1 U584 ( .A1(n520), .A2(n526), .ZN(n522) );
  XNOR2_X1 U585 ( .A(G85GAT), .B(KEYINPUT107), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n522), .B(n521), .ZN(G1336GAT) );
  NOR2_X1 U587 ( .A1(n523), .A2(n526), .ZN(n524) );
  XOR2_X1 U588 ( .A(G92GAT), .B(n524), .Z(G1337GAT) );
  NOR2_X1 U589 ( .A1(n535), .A2(n526), .ZN(n525) );
  XOR2_X1 U590 ( .A(G99GAT), .B(n525), .Z(G1338GAT) );
  NOR2_X1 U591 ( .A1(n533), .A2(n526), .ZN(n528) );
  XNOR2_X1 U592 ( .A(KEYINPUT108), .B(KEYINPUT44), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U594 ( .A(G106GAT), .B(n529), .Z(G1339GAT) );
  XOR2_X1 U595 ( .A(G113GAT), .B(KEYINPUT113), .Z(n537) );
  INV_X1 U596 ( .A(n530), .ZN(n531) );
  NOR2_X1 U597 ( .A1(n532), .A2(n531), .ZN(n549) );
  NAND2_X1 U598 ( .A1(n549), .A2(n533), .ZN(n534) );
  NOR2_X1 U599 ( .A1(n535), .A2(n534), .ZN(n546) );
  NAND2_X1 U600 ( .A1(n546), .A2(n559), .ZN(n536) );
  XNOR2_X1 U601 ( .A(n537), .B(n536), .ZN(G1340GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT114), .B(KEYINPUT49), .Z(n540) );
  NAND2_X1 U603 ( .A1(n546), .A2(n538), .ZN(n539) );
  XNOR2_X1 U604 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U605 ( .A(G120GAT), .B(n541), .ZN(G1341GAT) );
  INV_X1 U606 ( .A(n546), .ZN(n542) );
  NOR2_X1 U607 ( .A1(n563), .A2(n542), .ZN(n544) );
  XNOR2_X1 U608 ( .A(KEYINPUT115), .B(KEYINPUT50), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U610 ( .A(G127GAT), .B(n545), .ZN(G1342GAT) );
  XOR2_X1 U611 ( .A(G134GAT), .B(KEYINPUT51), .Z(n548) );
  NAND2_X1 U612 ( .A1(n546), .A2(n565), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n548), .B(n547), .ZN(G1343GAT) );
  NAND2_X1 U614 ( .A1(n549), .A2(n571), .ZN(n556) );
  NOR2_X1 U615 ( .A1(n573), .A2(n556), .ZN(n550) );
  XOR2_X1 U616 ( .A(G141GAT), .B(n550), .Z(n551) );
  XNOR2_X1 U617 ( .A(KEYINPUT116), .B(n551), .ZN(G1344GAT) );
  NOR2_X1 U618 ( .A1(n480), .A2(n556), .ZN(n553) );
  XNOR2_X1 U619 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(n554), .ZN(G1345GAT) );
  NOR2_X1 U622 ( .A1(n584), .A2(n556), .ZN(n555) );
  XOR2_X1 U623 ( .A(G155GAT), .B(n555), .Z(G1346GAT) );
  NOR2_X1 U624 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U625 ( .A(G162GAT), .B(n558), .Z(G1347GAT) );
  NAND2_X1 U626 ( .A1(n566), .A2(n559), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n560), .B(KEYINPUT118), .ZN(n561) );
  XNOR2_X1 U628 ( .A(G169GAT), .B(n561), .ZN(G1348GAT) );
  INV_X1 U629 ( .A(n566), .ZN(n562) );
  NOR2_X1 U630 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U631 ( .A(G183GAT), .B(n564), .Z(G1350GAT) );
  XNOR2_X1 U632 ( .A(G190GAT), .B(KEYINPUT120), .ZN(n570) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n568) );
  XOR2_X1 U634 ( .A(KEYINPUT121), .B(KEYINPUT58), .Z(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(G1351GAT) );
  NAND2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n587) );
  NOR2_X1 U638 ( .A1(n573), .A2(n587), .ZN(n578) );
  XOR2_X1 U639 ( .A(KEYINPUT60), .B(KEYINPUT123), .Z(n575) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT122), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(KEYINPUT59), .B(n576), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1352GAT) );
  NOR2_X1 U644 ( .A1(n587), .A2(n579), .ZN(n583) );
  XOR2_X1 U645 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n581) );
  XNOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT125), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1353GAT) );
  NOR2_X1 U649 ( .A1(n584), .A2(n587), .ZN(n585) );
  XOR2_X1 U650 ( .A(KEYINPUT126), .B(n585), .Z(n586) );
  XNOR2_X1 U651 ( .A(G211GAT), .B(n586), .ZN(G1354GAT) );
  NOR2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n590) );
  XNOR2_X1 U653 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

