//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 0 1 0 0 1 1 0 0 1 1 1 1 1 1 1 0 1 0 0 1 1 1 0 0 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 0 1 1 0 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n797, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n880, new_n881, new_n883, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n945, new_n946,
    new_n947, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n978, new_n979, new_n980, new_n981;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G64gat), .B(G92gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n202), .B(new_n203), .Z(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G226gat), .A2(G233gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT66), .ZN(new_n208));
  INV_X1    g007(.A(G169gat), .ZN(new_n209));
  INV_X1    g008(.A(G176gat), .ZN(new_n210));
  NAND4_X1  g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .A4(KEYINPUT26), .ZN(new_n211));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212));
  NOR3_X1   g011(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT26), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n211), .B(new_n212), .C1(new_n213), .C2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT67), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n219), .A2(new_n215), .A3(new_n214), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT67), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n220), .A2(new_n221), .A3(new_n212), .A4(new_n211), .ZN(new_n222));
  INV_X1    g021(.A(G183gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT27), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT27), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G183gat), .ZN(new_n226));
  INV_X1    g025(.A(G190gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n224), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT28), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(KEYINPUT65), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(KEYINPUT27), .B(G183gat), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n232), .A2(KEYINPUT65), .A3(new_n229), .A4(new_n227), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n218), .A2(new_n222), .A3(new_n231), .A4(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n209), .A2(new_n210), .A3(KEYINPUT23), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT23), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n236), .B1(G169gat), .B2(G176gat), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n235), .A2(new_n237), .A3(KEYINPUT25), .A4(new_n214), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT64), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n212), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT24), .ZN(new_n242));
  NAND3_X1  g041(.A1(KEYINPUT64), .A2(G183gat), .A3(G190gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  AND3_X1   g043(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n245));
  NOR2_X1   g044(.A1(G183gat), .A2(G190gat), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n239), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT25), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n251));
  NOR3_X1   g050(.A1(new_n245), .A2(new_n251), .A3(new_n246), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n235), .A2(new_n237), .A3(new_n214), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n250), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n249), .A2(new_n254), .ZN(new_n255));
  AND3_X1   g054(.A1(new_n234), .A2(new_n255), .A3(KEYINPUT73), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT73), .B1(new_n234), .B2(new_n255), .ZN(new_n257));
  OAI211_X1 g056(.A(KEYINPUT74), .B(new_n207), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n233), .B(new_n231), .C1(new_n217), .C2(KEYINPUT67), .ZN(new_n259));
  AND2_X1   g058(.A1(new_n217), .A2(KEYINPUT67), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n238), .B1(new_n247), .B2(new_n244), .ZN(new_n261));
  AND3_X1   g060(.A1(new_n235), .A2(new_n237), .A3(new_n214), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n212), .A2(new_n242), .ZN(new_n263));
  NAND3_X1  g062(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n263), .B(new_n264), .C1(G183gat), .C2(G190gat), .ZN(new_n265));
  AOI21_X1  g064(.A(KEYINPUT25), .B1(new_n262), .B2(new_n265), .ZN(new_n266));
  OAI22_X1  g065(.A1(new_n259), .A2(new_n260), .B1(new_n261), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT73), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n234), .A2(new_n255), .A3(KEYINPUT73), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n206), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT74), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT29), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n267), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n272), .B1(new_n274), .B2(new_n206), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n258), .B1(new_n271), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT75), .ZN(new_n277));
  XNOR2_X1  g076(.A(KEYINPUT72), .B(G197gat), .ZN(new_n278));
  INV_X1    g077(.A(G204gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT22), .ZN(new_n281));
  INV_X1    g080(.A(G211gat), .ZN(new_n282));
  INV_X1    g081(.A(G218gat), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n280), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G211gat), .B(G218gat), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n280), .A2(new_n286), .A3(new_n284), .ZN(new_n289));
  AND2_X1   g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n276), .A2(new_n277), .A3(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT76), .ZN(new_n292));
  INV_X1    g091(.A(new_n290), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n207), .B1(new_n256), .B2(new_n257), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT29), .B1(new_n234), .B2(new_n255), .ZN(new_n295));
  OAI21_X1  g094(.A(KEYINPUT74), .B1(new_n295), .B2(new_n207), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n293), .B1(new_n297), .B2(new_n258), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n267), .A2(new_n206), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n269), .A2(new_n270), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n207), .A2(KEYINPUT29), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(KEYINPUT75), .B1(new_n302), .B2(new_n290), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n291), .B(new_n292), .C1(new_n298), .C2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n276), .A2(new_n290), .ZN(new_n306));
  INV_X1    g105(.A(new_n299), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n256), .A2(new_n257), .ZN(new_n308));
  INV_X1    g107(.A(new_n301), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n277), .B1(new_n310), .B2(new_n293), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n292), .B1(new_n312), .B2(new_n291), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n205), .B1(new_n305), .B2(new_n313), .ZN(new_n314));
  XOR2_X1   g113(.A(G1gat), .B(G29gat), .Z(new_n315));
  XNOR2_X1  g114(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n315), .B(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G57gat), .B(G85gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n317), .B(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  XOR2_X1   g119(.A(KEYINPUT80), .B(G155gat), .Z(new_n321));
  INV_X1    g120(.A(G162gat), .ZN(new_n322));
  OAI21_X1  g121(.A(KEYINPUT2), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  XOR2_X1   g122(.A(G155gat), .B(G162gat), .Z(new_n324));
  XNOR2_X1  g123(.A(G141gat), .B(G148gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT78), .B1(G155gat), .B2(G162gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(G155gat), .B(G162gat), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n328), .B1(new_n329), .B2(KEYINPUT78), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT2), .ZN(new_n331));
  OR2_X1    g130(.A1(new_n331), .A2(KEYINPUT79), .ZN(new_n332));
  AOI22_X1  g131(.A1(new_n331), .A2(KEYINPUT79), .B1(G155gat), .B2(G162gat), .ZN(new_n333));
  AND2_X1   g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n330), .B1(new_n334), .B2(new_n325), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT3), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n327), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(G120gat), .ZN(new_n338));
  OAI21_X1  g137(.A(KEYINPUT69), .B1(new_n338), .B2(G113gat), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT69), .ZN(new_n340));
  INV_X1    g139(.A(G113gat), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n340), .A2(new_n341), .A3(G120gat), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n339), .B(new_n342), .C1(new_n341), .C2(G120gat), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT1), .ZN(new_n344));
  INV_X1    g143(.A(G134gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(G127gat), .ZN(new_n346));
  INV_X1    g145(.A(G127gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(G134gat), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n343), .A2(new_n344), .A3(new_n346), .A4(new_n348), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n341), .A2(G120gat), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n338), .A2(G113gat), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n344), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT68), .ZN(new_n353));
  AND3_X1   g152(.A1(new_n346), .A2(new_n348), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n353), .B1(new_n346), .B2(new_n348), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n352), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n349), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n337), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n336), .B1(new_n327), .B2(new_n335), .ZN(new_n359));
  OAI21_X1  g158(.A(KEYINPUT81), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n359), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT81), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n361), .A2(new_n362), .A3(new_n357), .A4(new_n337), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  AND2_X1   g163(.A1(new_n327), .A2(new_n335), .ZN(new_n365));
  INV_X1    g164(.A(new_n357), .ZN(new_n366));
  XOR2_X1   g165(.A(KEYINPUT82), .B(KEYINPUT4), .Z(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n365), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n327), .A2(new_n335), .A3(new_n356), .A4(new_n349), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT4), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AND3_X1   g171(.A1(new_n369), .A2(KEYINPUT84), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT84), .B1(new_n369), .B2(new_n372), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n364), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(G225gat), .A2(G233gat), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n377), .A2(KEYINPUT5), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n375), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n365), .A2(new_n366), .ZN(new_n381));
  INV_X1    g180(.A(new_n370), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n377), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(KEYINPUT5), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n376), .B1(new_n370), .B2(new_n371), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n385), .B1(new_n370), .B2(new_n367), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n384), .B1(new_n364), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n320), .B1(new_n380), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n364), .A2(new_n386), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n389), .A2(KEYINPUT5), .A3(new_n383), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n390), .B(new_n319), .C1(new_n375), .C2(new_n379), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT6), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n388), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  OAI211_X1 g192(.A(KEYINPUT6), .B(new_n320), .C1(new_n380), .C2(new_n387), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n205), .B1(new_n312), .B2(new_n291), .ZN(new_n396));
  OAI21_X1  g195(.A(KEYINPUT30), .B1(new_n396), .B2(KEYINPUT77), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n303), .A2(new_n298), .ZN(new_n398));
  AOI211_X1 g197(.A(KEYINPUT75), .B(new_n293), .C1(new_n297), .C2(new_n258), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n204), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT77), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT30), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n314), .A2(new_n395), .A3(new_n397), .A4(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(KEYINPUT31), .B(G50gat), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n337), .A2(new_n273), .ZN(new_n406));
  AOI22_X1  g205(.A1(new_n290), .A2(new_n406), .B1(G228gat), .B2(G233gat), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n327), .A2(new_n335), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT29), .B1(new_n288), .B2(new_n289), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n408), .B1(new_n409), .B2(KEYINPUT3), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(G228gat), .A2(G233gat), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n406), .A2(KEYINPUT85), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT85), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n337), .A2(new_n415), .A3(new_n273), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n414), .A2(new_n290), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n413), .B1(new_n410), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n405), .B1(new_n412), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n405), .ZN(new_n420));
  AND2_X1   g219(.A1(new_n410), .A2(new_n417), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n411), .B(new_n420), .C1(new_n421), .C2(new_n413), .ZN(new_n422));
  XNOR2_X1  g221(.A(G78gat), .B(G106gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n423), .B(G22gat), .ZN(new_n424));
  AND3_X1   g223(.A1(new_n419), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n424), .B1(new_n419), .B2(new_n422), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n404), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT36), .ZN(new_n430));
  AND3_X1   g229(.A1(new_n234), .A2(new_n255), .A3(new_n357), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n357), .B1(new_n234), .B2(new_n255), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(G227gat), .ZN(new_n434));
  INV_X1    g233(.A(G233gat), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT70), .B1(new_n433), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n267), .A2(new_n366), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n234), .A2(new_n255), .A3(new_n357), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n438), .A2(KEYINPUT70), .A3(new_n436), .A4(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(KEYINPUT32), .B1(new_n437), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT33), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n443), .B1(new_n437), .B2(new_n441), .ZN(new_n444));
  XNOR2_X1  g243(.A(G15gat), .B(G43gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(G71gat), .B(G99gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n445), .B(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n442), .A2(new_n444), .A3(new_n448), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n433), .A2(new_n436), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT34), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n436), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n451), .B(new_n453), .C1(new_n431), .C2(new_n432), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT32), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n438), .A2(new_n436), .A3(new_n439), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT70), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n457), .B1(new_n460), .B2(new_n440), .ZN(new_n461));
  AND2_X1   g260(.A1(new_n447), .A2(KEYINPUT71), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n447), .A2(KEYINPUT71), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n462), .A2(new_n463), .A3(new_n443), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  AND3_X1   g265(.A1(new_n449), .A2(new_n456), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n456), .B1(new_n449), .B2(new_n466), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n430), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n456), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT33), .B1(new_n460), .B2(new_n440), .ZN(new_n471));
  NOR3_X1   g270(.A1(new_n461), .A2(new_n471), .A3(new_n447), .ZN(new_n472));
  INV_X1    g271(.A(new_n466), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n470), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n449), .A2(new_n456), .A3(new_n466), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n474), .A2(KEYINPUT36), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n469), .A2(new_n476), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n429), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n314), .A2(new_n397), .A3(new_n403), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT39), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n381), .A2(new_n382), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n480), .B1(new_n481), .B2(new_n376), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT84), .ZN(new_n483));
  INV_X1    g282(.A(new_n372), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n370), .A2(new_n367), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n369), .A2(KEYINPUT84), .A3(new_n372), .ZN(new_n487));
  AOI22_X1  g286(.A1(new_n486), .A2(new_n487), .B1(new_n360), .B2(new_n363), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n482), .B1(new_n488), .B2(new_n376), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n375), .A2(new_n480), .A3(new_n377), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n489), .A2(new_n490), .A3(new_n319), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT40), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n491), .A2(new_n492), .ZN(new_n494));
  INV_X1    g293(.A(new_n388), .ZN(new_n495));
  NOR3_X1   g294(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n428), .B1(new_n479), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n395), .A2(new_n396), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT37), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT76), .B1(new_n398), .B2(new_n399), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n499), .B1(new_n500), .B2(new_n304), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n499), .B1(new_n398), .B2(new_n399), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n502), .A2(KEYINPUT38), .A3(new_n205), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n312), .A2(new_n291), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n204), .B1(new_n505), .B2(new_n499), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT86), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n302), .A2(new_n507), .A3(new_n290), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n276), .A2(new_n290), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT86), .B1(new_n310), .B2(new_n293), .ZN(new_n510));
  OAI211_X1 g309(.A(KEYINPUT37), .B(new_n508), .C1(new_n509), .C2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(KEYINPUT38), .B1(new_n506), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n498), .B1(new_n504), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n478), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n467), .A2(new_n468), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT87), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(new_n517), .A3(new_n427), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n404), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT35), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g320(.A(KEYINPUT35), .B1(new_n404), .B2(new_n518), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n515), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT92), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT18), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(G29gat), .A2(G36gat), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT14), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(G29gat), .A2(G36gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(G43gat), .B(G50gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT15), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT88), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n533), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT15), .ZN(new_n539));
  INV_X1    g338(.A(G43gat), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n540), .A2(KEYINPUT88), .A3(G50gat), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n538), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n531), .B(KEYINPUT89), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n530), .A2(new_n534), .A3(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n536), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(G15gat), .B(G22gat), .ZN(new_n547));
  OR2_X1    g346(.A1(new_n547), .A2(G1gat), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT16), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n547), .B1(new_n549), .B2(G1gat), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT90), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n548), .B(new_n550), .C1(new_n551), .C2(G8gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n548), .A2(new_n550), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n548), .A2(new_n551), .ZN(new_n554));
  INV_X1    g353(.A(G8gat), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n546), .A2(new_n552), .A3(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT17), .ZN(new_n559));
  OAI21_X1  g358(.A(KEYINPUT91), .B1(new_n546), .B2(new_n559), .ZN(new_n560));
  AND3_X1   g359(.A1(new_n530), .A2(new_n534), .A3(new_n544), .ZN(new_n561));
  AOI22_X1  g360(.A1(new_n561), .A2(new_n542), .B1(new_n532), .B2(new_n535), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT91), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n562), .A2(new_n563), .A3(KEYINPUT17), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  AOI22_X1  g364(.A1(new_n546), .A2(new_n559), .B1(new_n556), .B2(new_n552), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n558), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(G229gat), .A2(G233gat), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n527), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G113gat), .B(G141gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(G197gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(KEYINPUT11), .B(G169gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT12), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n556), .A2(new_n552), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(new_n546), .ZN(new_n578));
  XOR2_X1   g377(.A(new_n568), .B(KEYINPUT13), .Z(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  OR2_X1    g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n582), .A2(new_n527), .A3(new_n568), .A4(new_n557), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n570), .A2(new_n576), .A3(new_n581), .A4(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n581), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n575), .B1(new_n585), .B2(new_n569), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n524), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(G57gat), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n589), .A2(KEYINPUT93), .ZN(new_n590));
  INV_X1    g389(.A(G64gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G71gat), .A2(G78gat), .ZN(new_n593));
  OR2_X1    g392(.A1(G71gat), .A2(G78gat), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT9), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n589), .A2(new_n591), .ZN(new_n598));
  OAI21_X1  g397(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n599));
  OAI211_X1 g398(.A(new_n593), .B(new_n594), .C1(new_n598), .C2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n602), .A2(KEYINPUT21), .ZN(new_n603));
  XOR2_X1   g402(.A(KEYINPUT95), .B(KEYINPUT19), .Z(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n602), .A2(KEYINPUT21), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(new_n577), .ZN(new_n607));
  OR2_X1    g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n605), .A2(new_n607), .ZN(new_n609));
  XNOR2_X1  g408(.A(G127gat), .B(G155gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT20), .ZN(new_n611));
  NAND2_X1  g410(.A1(G231gat), .A2(G233gat), .ZN(new_n612));
  XOR2_X1   g411(.A(new_n612), .B(KEYINPUT94), .Z(new_n613));
  XNOR2_X1  g412(.A(new_n611), .B(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(G183gat), .B(G211gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  AND3_X1   g415(.A1(new_n608), .A2(new_n609), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n616), .B1(new_n608), .B2(new_n609), .ZN(new_n618));
  OR2_X1    g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AND2_X1   g418(.A1(G232gat), .A2(G233gat), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n620), .A2(KEYINPUT41), .ZN(new_n621));
  XNOR2_X1  g420(.A(G134gat), .B(G162gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n546), .A2(new_n559), .ZN(new_n625));
  NAND2_X1  g424(.A1(G99gat), .A2(G106gat), .ZN(new_n626));
  OR2_X1    g425(.A1(new_n626), .A2(KEYINPUT98), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT8), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n628), .B1(new_n626), .B2(KEYINPUT98), .ZN(new_n629));
  INV_X1    g428(.A(G85gat), .ZN(new_n630));
  INV_X1    g429(.A(G92gat), .ZN(new_n631));
  AOI22_X1  g430(.A1(new_n627), .A2(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT96), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT7), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(KEYINPUT96), .A2(KEYINPUT7), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n635), .A2(G85gat), .A3(G92gat), .A4(new_n636), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n633), .B(new_n634), .C1(new_n630), .C2(new_n631), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n637), .A2(KEYINPUT97), .A3(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(KEYINPUT97), .B1(new_n637), .B2(new_n638), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n632), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  XOR2_X1   g441(.A(G99gat), .B(G106gat), .Z(new_n643));
  NOR2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n643), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n637), .A2(new_n638), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT97), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(new_n639), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n645), .B1(new_n649), .B2(new_n632), .ZN(new_n650));
  OAI211_X1 g449(.A(new_n565), .B(new_n625), .C1(new_n644), .C2(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n644), .A2(new_n650), .ZN(new_n652));
  AOI22_X1  g451(.A1(new_n652), .A2(new_n546), .B1(KEYINPUT41), .B2(new_n620), .ZN(new_n653));
  XOR2_X1   g452(.A(G190gat), .B(G218gat), .Z(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n651), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n655), .B1(new_n651), .B2(new_n653), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n624), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n658), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n660), .A2(new_n623), .A3(new_n656), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n619), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(G230gat), .A2(G233gat), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n601), .B1(new_n644), .B2(new_n650), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT10), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n642), .A2(new_n643), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n649), .A2(new_n645), .A3(new_n632), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n668), .A2(new_n602), .A3(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n666), .A2(new_n667), .A3(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n652), .A2(KEYINPUT10), .A3(new_n602), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT99), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n665), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n671), .A2(KEYINPUT99), .A3(new_n672), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n666), .A2(new_n670), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(new_n665), .ZN(new_n679));
  XOR2_X1   g478(.A(G120gat), .B(G148gat), .Z(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT100), .ZN(new_n681));
  XNOR2_X1  g480(.A(G176gat), .B(G204gat), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n681), .B(new_n682), .Z(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n677), .A2(new_n679), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n665), .B1(new_n671), .B2(new_n672), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n679), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(new_n683), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n663), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n588), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n395), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(G1gat), .ZN(G1324gat));
  INV_X1    g495(.A(new_n479), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n588), .A2(new_n697), .A3(new_n692), .ZN(new_n698));
  XOR2_X1   g497(.A(KEYINPUT16), .B(G8gat), .Z(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n700), .B1(new_n555), .B2(new_n698), .ZN(new_n701));
  MUX2_X1   g500(.A(new_n700), .B(new_n701), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g501(.A(G15gat), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n693), .A2(new_n703), .A3(new_n516), .ZN(new_n704));
  AND3_X1   g503(.A1(new_n469), .A2(KEYINPUT101), .A3(new_n476), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT101), .B1(new_n469), .B2(new_n476), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT102), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n588), .A2(new_n692), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n704), .B1(new_n709), .B2(new_n703), .ZN(G1326gat));
  NAND2_X1  g509(.A1(new_n693), .A2(new_n428), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT103), .ZN(new_n712));
  XNOR2_X1  g511(.A(KEYINPUT43), .B(G22gat), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n712), .B(new_n713), .ZN(G1327gat));
  INV_X1    g513(.A(new_n662), .ZN(new_n715));
  INV_X1    g514(.A(new_n690), .ZN(new_n716));
  INV_X1    g515(.A(new_n619), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n587), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AND3_X1   g519(.A1(new_n524), .A2(new_n715), .A3(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(G29gat), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n721), .A2(new_n722), .A3(new_n694), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT45), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n662), .A2(KEYINPUT44), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT104), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n514), .A2(new_n726), .A3(new_n429), .A4(new_n707), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(new_n523), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n469), .A2(KEYINPUT101), .A3(new_n476), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT101), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n477), .A2(new_n730), .ZN(new_n731));
  AND3_X1   g530(.A1(new_n429), .A2(new_n729), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n726), .B1(new_n732), .B2(new_n514), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n725), .B1(new_n728), .B2(new_n733), .ZN(new_n734));
  AOI22_X1  g533(.A1(new_n478), .A2(new_n514), .B1(new_n521), .B2(new_n522), .ZN(new_n735));
  OAI21_X1  g534(.A(KEYINPUT44), .B1(new_n735), .B2(new_n662), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n720), .ZN(new_n738));
  OAI21_X1  g537(.A(G29gat), .B1(new_n738), .B2(new_n395), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n739), .ZN(G1328gat));
  OAI21_X1  g539(.A(G36gat), .B1(new_n738), .B2(new_n697), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n718), .A2(G36gat), .A3(new_n662), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n524), .A2(new_n587), .A3(new_n479), .A4(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  OR2_X1    g544(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g545(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n743), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n741), .A2(new_n746), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(KEYINPUT106), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT106), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n741), .A2(new_n751), .A3(new_n746), .A4(new_n748), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(G1329gat));
  INV_X1    g552(.A(KEYINPUT47), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n474), .A2(new_n475), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n755), .A2(G43gat), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n721), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT107), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n721), .A2(KEYINPUT107), .A3(new_n756), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n754), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(KEYINPUT108), .B1(new_n738), .B2(new_n707), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(G43gat), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n738), .A2(KEYINPUT108), .A3(new_n707), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n761), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n737), .A2(new_n720), .ZN(new_n766));
  INV_X1    g565(.A(new_n708), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n540), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  AND2_X1   g567(.A1(new_n759), .A2(new_n760), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n754), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n765), .A2(new_n770), .ZN(G1330gat));
  AOI21_X1  g570(.A(G50gat), .B1(new_n721), .B2(new_n428), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n428), .A2(G50gat), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n772), .B1(new_n766), .B2(new_n773), .ZN(new_n774));
  XOR2_X1   g573(.A(new_n774), .B(KEYINPUT48), .Z(G1331gat));
  AND2_X1   g574(.A1(new_n497), .A2(new_n513), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n429), .A2(new_n729), .A3(new_n731), .ZN(new_n777));
  OAI21_X1  g576(.A(KEYINPUT104), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n778), .A2(new_n523), .A3(new_n727), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  NOR4_X1   g579(.A1(new_n780), .A2(new_n587), .A3(new_n663), .A4(new_n716), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n694), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n479), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n784), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n785));
  XOR2_X1   g584(.A(KEYINPUT49), .B(G64gat), .Z(new_n786));
  OAI21_X1  g585(.A(new_n785), .B1(new_n784), .B2(new_n786), .ZN(G1333gat));
  NAND2_X1  g586(.A1(new_n781), .A2(new_n767), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(G71gat), .ZN(new_n789));
  INV_X1    g588(.A(G71gat), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n781), .A2(new_n790), .A3(new_n516), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT50), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n789), .A2(KEYINPUT50), .A3(new_n791), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(G1334gat));
  NAND2_X1  g595(.A1(new_n781), .A2(new_n428), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n797), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g597(.A1(new_n717), .A2(new_n719), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n799), .A2(new_n716), .ZN(new_n800));
  XOR2_X1   g599(.A(new_n800), .B(KEYINPUT109), .Z(new_n801));
  AOI21_X1  g600(.A(new_n801), .B1(new_n734), .B2(new_n736), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(G85gat), .B1(new_n803), .B2(new_n395), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n799), .A2(new_n662), .ZN(new_n805));
  OAI211_X1 g604(.A(KEYINPUT51), .B(new_n805), .C1(new_n728), .C2(new_n733), .ZN(new_n806));
  OR2_X1    g605(.A1(new_n806), .A2(KEYINPUT110), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(KEYINPUT110), .ZN(new_n808));
  AOI21_X1  g607(.A(KEYINPUT51), .B1(new_n779), .B2(new_n805), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n807), .A2(new_n808), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n690), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n694), .A2(new_n630), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n804), .B1(new_n812), .B2(new_n813), .ZN(G1336gat));
  NOR3_X1   g613(.A1(new_n697), .A2(G92gat), .A3(new_n716), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n816), .B1(new_n810), .B2(new_n806), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n631), .B1(new_n802), .B2(new_n479), .ZN(new_n818));
  OAI21_X1  g617(.A(KEYINPUT52), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n811), .A2(new_n815), .ZN(new_n820));
  OR2_X1    g619(.A1(new_n818), .A2(KEYINPUT52), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(G1337gat));
  XOR2_X1   g621(.A(KEYINPUT111), .B(G99gat), .Z(new_n823));
  OAI21_X1  g622(.A(new_n823), .B1(new_n803), .B2(new_n708), .ZN(new_n824));
  OR2_X1    g623(.A1(new_n755), .A2(new_n823), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n824), .B1(new_n812), .B2(new_n825), .ZN(G1338gat));
  AOI211_X1 g625(.A(new_n427), .B(new_n801), .C1(new_n734), .C2(new_n736), .ZN(new_n827));
  INV_X1    g626(.A(G106gat), .ZN(new_n828));
  OAI21_X1  g627(.A(KEYINPUT112), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n716), .A2(new_n427), .A3(G106gat), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n830), .B(KEYINPUT113), .ZN(new_n831));
  INV_X1    g630(.A(new_n806), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n831), .B1(new_n832), .B2(new_n809), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT114), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(new_n801), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n737), .A2(new_n428), .A3(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT112), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n837), .A2(new_n838), .A3(G106gat), .ZN(new_n839));
  OAI211_X1 g638(.A(KEYINPUT114), .B(new_n831), .C1(new_n832), .C2(new_n809), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n829), .A2(new_n835), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(KEYINPUT53), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n811), .A2(new_n830), .ZN(new_n843));
  AOI21_X1  g642(.A(KEYINPUT53), .B1(new_n837), .B2(G106gat), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n842), .A2(new_n845), .ZN(G1339gat));
  NOR3_X1   g645(.A1(new_n663), .A2(new_n587), .A3(new_n690), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT55), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n671), .A2(new_n665), .A3(new_n672), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(KEYINPUT54), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n850), .B1(new_n675), .B2(new_n676), .ZN(new_n851));
  XOR2_X1   g650(.A(KEYINPUT115), .B(KEYINPUT54), .Z(new_n852));
  AOI21_X1  g651(.A(new_n684), .B1(new_n686), .B2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n848), .B1(new_n851), .B2(new_n854), .ZN(new_n855));
  AND3_X1   g654(.A1(new_n671), .A2(KEYINPUT99), .A3(new_n672), .ZN(new_n856));
  AOI21_X1  g655(.A(KEYINPUT99), .B1(new_n671), .B2(new_n672), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n856), .A2(new_n857), .A3(new_n665), .ZN(new_n858));
  OAI211_X1 g657(.A(KEYINPUT55), .B(new_n853), .C1(new_n858), .C2(new_n850), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n582), .A2(new_n557), .ZN(new_n860));
  INV_X1    g659(.A(new_n568), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n578), .A2(new_n580), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n574), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n585), .A2(new_n569), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n864), .B1(new_n865), .B2(new_n576), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n855), .A2(new_n859), .A3(new_n866), .A4(new_n685), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n619), .B1(new_n867), .B2(new_n715), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n855), .A2(new_n859), .A3(new_n587), .A4(new_n685), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n690), .A2(new_n866), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n869), .A2(new_n662), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n847), .B1(new_n868), .B2(new_n871), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n872), .A2(new_n755), .A3(new_n428), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n479), .A2(new_n395), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n875), .A2(new_n719), .ZN(new_n876));
  XNOR2_X1  g675(.A(new_n876), .B(new_n341), .ZN(G1340gat));
  NOR2_X1   g676(.A1(new_n875), .A2(new_n716), .ZN(new_n878));
  XNOR2_X1  g677(.A(new_n878), .B(new_n338), .ZN(G1341gat));
  NOR2_X1   g678(.A1(new_n875), .A2(new_n717), .ZN(new_n880));
  XOR2_X1   g679(.A(KEYINPUT116), .B(G127gat), .Z(new_n881));
  XNOR2_X1  g680(.A(new_n880), .B(new_n881), .ZN(G1342gat));
  NOR2_X1   g681(.A1(new_n479), .A2(new_n662), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n873), .A2(new_n345), .A3(new_n694), .A4(new_n883), .ZN(new_n884));
  XOR2_X1   g683(.A(new_n884), .B(KEYINPUT56), .Z(new_n885));
  OAI21_X1  g684(.A(G134gat), .B1(new_n875), .B2(new_n662), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(G1343gat));
  XNOR2_X1  g686(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n872), .A2(new_n427), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n708), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n874), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n719), .A2(G141gat), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT118), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n888), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n889), .A2(KEYINPUT57), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT57), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n898), .B1(new_n872), .B2(new_n427), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n707), .A2(new_n874), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  OR3_X1    g702(.A1(new_n903), .A2(KEYINPUT120), .A3(new_n719), .ZN(new_n904));
  OAI21_X1  g703(.A(KEYINPUT120), .B1(new_n903), .B2(new_n719), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n904), .A2(G141gat), .A3(new_n905), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n896), .B(new_n906), .C1(new_n895), .C2(new_n894), .ZN(new_n907));
  AOI21_X1  g706(.A(KEYINPUT117), .B1(new_n900), .B2(new_n902), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT117), .ZN(new_n909));
  AOI211_X1 g708(.A(new_n909), .B(new_n901), .C1(new_n897), .C2(new_n899), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(new_n587), .ZN(new_n912));
  AOI22_X1  g711(.A1(new_n912), .A2(G141gat), .B1(new_n892), .B2(new_n893), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT58), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n907), .B1(new_n913), .B2(new_n914), .ZN(G1344gat));
  INV_X1    g714(.A(G148gat), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n892), .A2(new_n916), .A3(new_n690), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT59), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n428), .B1(new_n872), .B2(KEYINPUT121), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT121), .ZN(new_n920));
  AOI211_X1 g719(.A(new_n920), .B(new_n847), .C1(new_n868), .C2(new_n871), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n898), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT122), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OAI211_X1 g723(.A(KEYINPUT122), .B(new_n898), .C1(new_n919), .C2(new_n921), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n924), .A2(new_n897), .A3(new_n925), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n901), .A2(new_n716), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n918), .B1(new_n928), .B2(G148gat), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n918), .A2(G148gat), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n930), .B1(new_n911), .B2(new_n690), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n917), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(KEYINPUT123), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT123), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n934), .B(new_n917), .C1(new_n929), .C2(new_n931), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n933), .A2(new_n935), .ZN(G1345gat));
  NAND3_X1  g735(.A1(new_n892), .A2(new_n321), .A3(new_n619), .ZN(new_n937));
  INV_X1    g736(.A(new_n911), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n938), .A2(new_n717), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n937), .B1(new_n939), .B2(new_n321), .ZN(G1346gat));
  NAND4_X1  g739(.A1(new_n890), .A2(new_n322), .A3(new_n694), .A4(new_n883), .ZN(new_n941));
  XOR2_X1   g740(.A(new_n941), .B(KEYINPUT124), .Z(new_n942));
  OAI21_X1  g741(.A(G162gat), .B1(new_n938), .B2(new_n662), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(G1347gat));
  NOR2_X1   g743(.A1(new_n697), .A2(new_n694), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n873), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(new_n587), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g747(.A1(new_n946), .A2(new_n690), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g749(.A1(new_n946), .A2(new_n619), .ZN(new_n951));
  AOI21_X1  g750(.A(KEYINPUT126), .B1(new_n951), .B2(G183gat), .ZN(new_n952));
  INV_X1    g751(.A(new_n232), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n954), .A2(KEYINPUT125), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n954), .A2(KEYINPUT125), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n952), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n957), .B(KEYINPUT60), .ZN(G1350gat));
  NOR2_X1   g757(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n959), .B1(new_n946), .B2(new_n715), .ZN(new_n960));
  NAND2_X1  g759(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n961));
  XOR2_X1   g760(.A(new_n960), .B(new_n961), .Z(G1351gat));
  AND2_X1   g761(.A1(new_n708), .A2(new_n945), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n963), .A2(new_n889), .ZN(new_n964));
  AOI21_X1  g763(.A(G197gat), .B1(new_n964), .B2(new_n587), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n926), .A2(new_n963), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n587), .A2(G197gat), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n965), .B1(new_n966), .B2(new_n967), .ZN(G1352gat));
  NAND3_X1  g767(.A1(new_n964), .A2(new_n279), .A3(new_n690), .ZN(new_n969));
  XOR2_X1   g768(.A(new_n969), .B(KEYINPUT62), .Z(new_n970));
  AND2_X1   g769(.A1(new_n966), .A2(new_n690), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n970), .B1(new_n279), .B2(new_n971), .ZN(G1353gat));
  NAND3_X1  g771(.A1(new_n964), .A2(new_n282), .A3(new_n619), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n966), .A2(new_n619), .ZN(new_n974));
  AND3_X1   g773(.A1(new_n974), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n975));
  AOI21_X1  g774(.A(KEYINPUT63), .B1(new_n974), .B2(G211gat), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n973), .B1(new_n975), .B2(new_n976), .ZN(G1354gat));
  NAND3_X1  g776(.A1(new_n963), .A2(new_n715), .A3(new_n889), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n978), .A2(new_n283), .ZN(new_n979));
  XNOR2_X1  g778(.A(new_n979), .B(KEYINPUT127), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n662), .A2(new_n283), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n980), .B1(new_n966), .B2(new_n981), .ZN(G1355gat));
endmodule


