//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 0 1 0 1 1 0 1 0 1 1 1 0 0 0 1 0 0 0 1 1 0 1 1 0 1 0 1 0 0 1 1 0 1 1 0 0 1 1 0 0 1 1 1 1 0 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n757, new_n758,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n835,
    new_n836, new_n837, new_n838, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n982, new_n983, new_n984;
  XNOR2_X1  g000(.A(G127gat), .B(G155gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G211gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT94), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT91), .B(G57gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G64gat), .ZN(new_n207));
  INV_X1    g006(.A(G64gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G57gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n207), .A2(KEYINPUT92), .A3(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT92), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT91), .ZN(new_n212));
  INV_X1    g011(.A(G57gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(KEYINPUT91), .A2(G57gat), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n208), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n209), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n211), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G71gat), .A2(G78gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(G71gat), .A2(G78gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT9), .ZN(new_n221));
  AOI22_X1  g020(.A1(new_n210), .A2(new_n218), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n219), .B(KEYINPUT90), .ZN(new_n223));
  NOR2_X1   g022(.A1(KEYINPUT90), .A2(KEYINPUT9), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n213), .A2(G64gat), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n224), .B1(new_n209), .B2(new_n225), .ZN(new_n226));
  NOR3_X1   g025(.A1(new_n223), .A2(new_n226), .A3(new_n220), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n205), .B1(new_n222), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n221), .A2(new_n219), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT92), .B1(new_n207), .B2(new_n209), .ZN(new_n230));
  NOR3_X1   g029(.A1(new_n216), .A2(new_n211), .A3(new_n217), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n227), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n232), .A2(KEYINPUT94), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n228), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT21), .ZN(new_n236));
  INV_X1    g035(.A(G183gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(G15gat), .B(G22gat), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT16), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n238), .B1(new_n239), .B2(G1gat), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n240), .B1(G1gat), .B2(new_n238), .ZN(new_n241));
  INV_X1    g040(.A(G8gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n241), .B(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n236), .A2(new_n237), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n237), .B1(new_n236), .B2(new_n243), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n222), .A2(new_n227), .ZN(new_n247));
  XNOR2_X1  g046(.A(KEYINPUT93), .B(KEYINPUT21), .ZN(new_n248));
  OAI22_X1  g047(.A1(new_n245), .A2(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n246), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n247), .A2(new_n248), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n250), .A2(new_n244), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n204), .B1(new_n249), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n255));
  NAND2_X1  g054(.A1(G231gat), .A2(G233gat), .ZN(new_n256));
  XOR2_X1   g055(.A(new_n255), .B(new_n256), .Z(new_n257));
  NAND3_X1  g056(.A1(new_n249), .A2(new_n252), .A3(new_n204), .ZN(new_n258));
  AND3_X1   g057(.A1(new_n254), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n257), .B1(new_n254), .B2(new_n258), .ZN(new_n260));
  OR2_X1    g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(G232gat), .A2(G233gat), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n263), .A2(KEYINPUT41), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n264), .B(KEYINPUT95), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n265), .B(G190gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n266), .B(G218gat), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT88), .ZN(new_n269));
  XOR2_X1   g068(.A(G43gat), .B(G50gat), .Z(new_n270));
  INV_X1    g069(.A(KEYINPUT15), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G43gat), .B(G50gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT15), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT14), .ZN(new_n275));
  INV_X1    g074(.A(G29gat), .ZN(new_n276));
  INV_X1    g075(.A(G36gat), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n279));
  AOI22_X1  g078(.A1(new_n278), .A2(new_n279), .B1(G29gat), .B2(G36gat), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n272), .A2(new_n274), .A3(new_n280), .ZN(new_n281));
  AND2_X1   g080(.A1(new_n278), .A2(new_n279), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n276), .A2(new_n277), .ZN(new_n283));
  OAI211_X1 g082(.A(KEYINPUT15), .B(new_n273), .C1(new_n282), .C2(new_n283), .ZN(new_n284));
  AND2_X1   g083(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n269), .B1(new_n285), .B2(KEYINPUT87), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT17), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n281), .A2(new_n284), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n287), .B1(new_n288), .B2(KEYINPUT88), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n269), .B(new_n287), .C1(new_n285), .C2(KEYINPUT87), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT97), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n293), .A2(KEYINPUT7), .ZN(new_n294));
  NAND2_X1  g093(.A1(G85gat), .A2(G92gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(G99gat), .A2(G106gat), .ZN(new_n296));
  AOI22_X1  g095(.A1(new_n294), .A2(new_n295), .B1(KEYINPUT8), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT7), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT97), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n293), .A2(KEYINPUT7), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n299), .A2(new_n300), .A3(G85gat), .A4(G92gat), .ZN(new_n301));
  INV_X1    g100(.A(G85gat), .ZN(new_n302));
  INV_X1    g101(.A(G92gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n297), .A2(new_n301), .A3(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G99gat), .B(G106gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n297), .A2(new_n301), .A3(new_n306), .A4(new_n304), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AOI22_X1  g109(.A1(new_n292), .A2(new_n310), .B1(KEYINPUT41), .B2(new_n263), .ZN(new_n311));
  XNOR2_X1  g110(.A(G134gat), .B(G162gat), .ZN(new_n312));
  XOR2_X1   g111(.A(new_n312), .B(KEYINPUT96), .Z(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  AND2_X1   g113(.A1(new_n308), .A2(new_n309), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(new_n288), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n311), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n314), .B1(new_n311), .B2(new_n316), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n268), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n311), .A2(new_n316), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(new_n313), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n322), .A2(new_n267), .A3(new_n317), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n261), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(G176gat), .ZN(new_n326));
  AND2_X1   g125(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n328));
  OAI211_X1 g127(.A(KEYINPUT23), .B(new_n326), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(G183gat), .A2(G190gat), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT24), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n333));
  INV_X1    g132(.A(G190gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n237), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n332), .A2(new_n333), .A3(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(G169gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(new_n326), .ZN(new_n338));
  NAND2_X1  g137(.A1(G169gat), .A2(G176gat), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT23), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n338), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n329), .A2(new_n336), .A3(new_n342), .ZN(new_n343));
  XOR2_X1   g142(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n332), .A2(new_n333), .ZN(new_n346));
  XNOR2_X1  g145(.A(KEYINPUT66), .B(G183gat), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT67), .B1(new_n347), .B2(G190gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n237), .A2(KEYINPUT66), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT66), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(G183gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT67), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n352), .A2(new_n353), .A3(new_n334), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n346), .B1(new_n348), .B2(new_n354), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n342), .B(KEYINPUT25), .C1(new_n341), .C2(new_n338), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n345), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(KEYINPUT27), .B(G183gat), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n358), .A2(KEYINPUT28), .A3(new_n334), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n349), .A2(new_n351), .A3(KEYINPUT27), .ZN(new_n360));
  OR2_X1    g159(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n361));
  AOI21_X1  g160(.A(G190gat), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n359), .B1(new_n362), .B2(KEYINPUT28), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n338), .A2(KEYINPUT26), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n364), .A2(new_n340), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n338), .A2(KEYINPUT26), .ZN(new_n366));
  AOI22_X1  g165(.A1(new_n365), .A2(new_n366), .B1(G183gat), .B2(G190gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n363), .A2(new_n367), .ZN(new_n368));
  XOR2_X1   g167(.A(G127gat), .B(G134gat), .Z(new_n369));
  OR2_X1    g168(.A1(KEYINPUT68), .A2(KEYINPUT1), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G113gat), .B(G120gat), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n372), .A2(KEYINPUT1), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n369), .B(new_n370), .C1(KEYINPUT1), .C2(new_n372), .ZN(new_n375));
  AND2_X1   g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n357), .A2(new_n368), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT69), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n357), .A2(new_n368), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n374), .A2(new_n375), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(G227gat), .A2(G233gat), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT69), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n357), .A2(new_n368), .A3(new_n383), .A4(new_n376), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n378), .A2(new_n381), .A3(new_n382), .A4(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n385), .B(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT32), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n378), .A2(new_n381), .A3(new_n384), .ZN(new_n390));
  INV_X1    g189(.A(new_n382), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n389), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT33), .ZN(new_n393));
  XNOR2_X1  g192(.A(G15gat), .B(G43gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n394), .B(G71gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n395), .B(G99gat), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n392), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n390), .A2(new_n391), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT32), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n393), .ZN(new_n401));
  INV_X1    g200(.A(new_n396), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT70), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n396), .B1(new_n399), .B2(KEYINPUT32), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT70), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n405), .A2(new_n406), .A3(new_n401), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n398), .B1(new_n404), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n388), .B1(new_n408), .B2(KEYINPUT72), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT33), .B1(new_n390), .B2(new_n391), .ZN(new_n410));
  NOR4_X1   g209(.A1(new_n392), .A2(new_n410), .A3(KEYINPUT70), .A4(new_n396), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n406), .B1(new_n405), .B2(new_n401), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n397), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT72), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n413), .A2(new_n414), .A3(new_n387), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n409), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT36), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT36), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n404), .A2(new_n407), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n387), .B1(new_n419), .B2(new_n397), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n397), .B(new_n387), .C1(new_n411), .C2(new_n412), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n418), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n417), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(G228gat), .A2(G233gat), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  XOR2_X1   g225(.A(G141gat), .B(G148gat), .Z(new_n427));
  INV_X1    g226(.A(KEYINPUT2), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  OR2_X1    g228(.A1(G155gat), .A2(G162gat), .ZN(new_n430));
  NAND2_X1  g229(.A1(G155gat), .A2(G162gat), .ZN(new_n431));
  AND2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n431), .B1(new_n430), .B2(KEYINPUT2), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT78), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n434), .A2(new_n427), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n435), .B1(new_n434), .B2(new_n427), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n433), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT3), .ZN(new_n440));
  INV_X1    g239(.A(G218gat), .ZN(new_n441));
  INV_X1    g240(.A(G197gat), .ZN(new_n442));
  INV_X1    g241(.A(G204gat), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(G197gat), .A2(G204gat), .ZN(new_n445));
  OR2_X1    g244(.A1(KEYINPUT73), .A2(G211gat), .ZN(new_n446));
  NAND2_X1  g245(.A1(KEYINPUT73), .A2(G211gat), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n446), .A2(G218gat), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT22), .ZN(new_n449));
  AOI221_X4 g248(.A(G211gat), .B1(new_n444), .B2(new_n445), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(G211gat), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n448), .A2(new_n449), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n444), .A2(new_n445), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n441), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  AND2_X1   g254(.A1(KEYINPUT73), .A2(G211gat), .ZN(new_n456));
  NOR2_X1   g255(.A1(KEYINPUT73), .A2(G211gat), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(KEYINPUT22), .B1(new_n458), .B2(G218gat), .ZN(new_n459));
  INV_X1    g258(.A(new_n453), .ZN(new_n460));
  OAI21_X1  g259(.A(G211gat), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n452), .A2(new_n451), .A3(new_n453), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n461), .A2(new_n462), .A3(G218gat), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT29), .B1(new_n455), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT82), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n440), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AOI211_X1 g265(.A(KEYINPUT82), .B(KEYINPUT29), .C1(new_n455), .C2(new_n463), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n439), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n455), .A2(new_n463), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT29), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n434), .A2(new_n427), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT78), .ZN(new_n472));
  AOI22_X1  g271(.A1(new_n472), .A2(new_n436), .B1(new_n429), .B2(new_n432), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(new_n440), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n469), .B1(new_n470), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n426), .B1(new_n468), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n464), .A2(new_n439), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n439), .A2(KEYINPUT3), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n476), .A2(new_n478), .A3(new_n479), .A4(new_n426), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(G22gat), .B1(new_n477), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(G22gat), .ZN(new_n483));
  NOR3_X1   g282(.A1(new_n450), .A2(new_n454), .A3(new_n441), .ZN(new_n484));
  AOI21_X1  g283(.A(G218gat), .B1(new_n461), .B2(new_n462), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n470), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT82), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n464), .A2(new_n465), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n487), .A2(new_n440), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n475), .B1(new_n489), .B2(new_n439), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n483), .B(new_n480), .C1(new_n490), .C2(new_n426), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n482), .A2(new_n491), .A3(KEYINPUT84), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT84), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n493), .B(G22gat), .C1(new_n477), .C2(new_n481), .ZN(new_n494));
  XNOR2_X1  g293(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(G50gat), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n496), .B(G78gat), .ZN(new_n497));
  INV_X1    g296(.A(G106gat), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n497), .B(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n492), .A2(new_n494), .A3(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT83), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n491), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT3), .B1(new_n486), .B2(KEYINPUT82), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n473), .B1(new_n504), .B2(new_n488), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n425), .B1(new_n505), .B2(new_n475), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n506), .A2(KEYINPUT83), .A3(new_n483), .A4(new_n480), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n503), .A2(new_n482), .A3(new_n499), .A4(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n501), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT80), .ZN(new_n510));
  NOR3_X1   g309(.A1(new_n439), .A2(KEYINPUT4), .A3(new_n380), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT4), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n512), .B1(new_n473), .B2(new_n376), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n510), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT4), .B1(new_n439), .B2(new_n380), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n473), .A2(new_n376), .A3(new_n512), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(new_n516), .A3(KEYINPUT80), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT5), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n474), .A2(new_n479), .A3(new_n380), .ZN(new_n520));
  NAND2_X1  g319(.A1(G225gat), .A2(G233gat), .ZN(new_n521));
  AND2_X1   g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n518), .A2(new_n519), .A3(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n439), .B(new_n380), .ZN(new_n524));
  INV_X1    g323(.A(new_n521), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT79), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n527), .B(KEYINPUT4), .C1(new_n439), .C2(new_n380), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n520), .A2(new_n521), .A3(new_n528), .ZN(new_n529));
  AND3_X1   g328(.A1(new_n515), .A2(new_n516), .A3(KEYINPUT79), .ZN(new_n530));
  OAI211_X1 g329(.A(KEYINPUT5), .B(new_n526), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n523), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(KEYINPUT0), .B(G57gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(G85gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(G1gat), .B(G29gat), .ZN(new_n535));
  XOR2_X1   g334(.A(new_n534), .B(new_n535), .Z(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n532), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT6), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n523), .A2(new_n531), .A3(new_n536), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n532), .A2(KEYINPUT6), .A3(new_n537), .ZN(new_n542));
  AND2_X1   g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(G226gat), .A2(G233gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(KEYINPUT74), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n357), .A2(new_n368), .A3(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n379), .ZN(new_n547));
  OR2_X1    g346(.A1(new_n545), .A2(KEYINPUT29), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n469), .B(new_n546), .C1(new_n547), .C2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n469), .ZN(new_n550));
  AND3_X1   g349(.A1(new_n357), .A2(new_n368), .A3(new_n545), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n548), .B1(new_n357), .B2(new_n368), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G8gat), .B(G36gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(G92gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(KEYINPUT75), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(new_n208), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n554), .A2(KEYINPUT30), .A3(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n560), .B1(new_n554), .B2(new_n559), .ZN(new_n561));
  AND3_X1   g360(.A1(new_n554), .A2(KEYINPUT76), .A3(new_n559), .ZN(new_n562));
  AOI21_X1  g361(.A(KEYINPUT76), .B1(new_n554), .B2(new_n559), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(KEYINPUT77), .B(KEYINPUT30), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n561), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n509), .B1(new_n543), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT37), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n559), .B1(new_n554), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n549), .A2(new_n553), .A3(KEYINPUT37), .ZN(new_n571));
  AND2_X1   g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT85), .ZN(new_n573));
  AOI21_X1  g372(.A(KEYINPUT38), .B1(new_n570), .B2(new_n573), .ZN(new_n574));
  AOI211_X1 g373(.A(new_n563), .B(new_n562), .C1(new_n572), .C2(new_n574), .ZN(new_n575));
  OAI211_X1 g374(.A(new_n543), .B(new_n575), .C1(new_n574), .C2(new_n572), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n518), .A2(new_n520), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(new_n525), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n578), .B(KEYINPUT39), .C1(new_n525), .C2(new_n524), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT39), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n577), .A2(new_n580), .A3(new_n525), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n579), .A2(new_n536), .A3(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT40), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n579), .A2(KEYINPUT40), .A3(new_n536), .A4(new_n581), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n584), .A2(new_n567), .A3(new_n538), .A4(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n483), .B1(new_n506), .B2(new_n480), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n587), .B1(new_n502), .B2(new_n491), .ZN(new_n588));
  AND2_X1   g387(.A1(new_n507), .A2(new_n499), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n499), .B1(new_n587), .B2(new_n493), .ZN(new_n590));
  AOI22_X1  g389(.A1(new_n588), .A2(new_n589), .B1(new_n590), .B2(new_n492), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n576), .A2(new_n586), .A3(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n424), .A2(new_n568), .A3(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT35), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n509), .B1(new_n415), .B2(new_n409), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n543), .A2(new_n567), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n413), .A2(new_n388), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n598), .A2(new_n501), .A3(new_n508), .A4(new_n421), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n541), .A2(new_n542), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n600), .A2(new_n594), .A3(new_n566), .ZN(new_n601));
  OAI21_X1  g400(.A(KEYINPUT86), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n420), .A2(new_n422), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT86), .ZN(new_n604));
  AND3_X1   g403(.A1(new_n600), .A2(new_n594), .A3(new_n566), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n603), .A2(new_n604), .A3(new_n591), .A4(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n593), .B1(new_n597), .B2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n243), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(new_n288), .ZN(new_n610));
  NAND2_X1  g409(.A1(G229gat), .A2(G233gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT89), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT87), .ZN(new_n613));
  AOI211_X1 g412(.A(KEYINPUT88), .B(KEYINPUT17), .C1(new_n288), .C2(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n614), .B1(new_n286), .B2(new_n289), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n610), .B(new_n612), .C1(new_n615), .C2(new_n609), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT18), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n609), .B(new_n285), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n612), .B(KEYINPUT13), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n292), .A2(new_n243), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n622), .A2(KEYINPUT18), .A3(new_n610), .A4(new_n612), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n618), .A2(new_n621), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT11), .B(G169gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(G197gat), .ZN(new_n626));
  XOR2_X1   g425(.A(G113gat), .B(G141gat), .Z(new_n627));
  XOR2_X1   g426(.A(new_n626), .B(new_n627), .Z(new_n628));
  XOR2_X1   g427(.A(new_n628), .B(KEYINPUT12), .Z(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n624), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n618), .A2(new_n623), .A3(new_n629), .A4(new_n621), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(G120gat), .B(G148gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(new_n326), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(new_n443), .ZN(new_n636));
  NAND2_X1  g435(.A1(G230gat), .A2(G233gat), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n637), .B(KEYINPUT99), .Z(new_n638));
  NAND3_X1  g437(.A1(new_n235), .A2(KEYINPUT10), .A3(new_n315), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n307), .A2(KEYINPUT98), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n232), .A2(new_n233), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(new_n310), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n315), .A2(new_n232), .A3(new_n233), .A4(new_n640), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT10), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n638), .B1(new_n639), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n638), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n647), .B1(new_n642), .B2(new_n643), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n636), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT100), .ZN(new_n651));
  NOR3_X1   g450(.A1(new_n646), .A2(new_n648), .A3(new_n636), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n652), .ZN(new_n655));
  AOI21_X1  g454(.A(KEYINPUT100), .B1(new_n655), .B2(new_n649), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  AND4_X1   g458(.A1(new_n325), .A2(new_n608), .A3(new_n633), .A4(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(new_n543), .ZN(new_n661));
  XNOR2_X1  g460(.A(KEYINPUT101), .B(G1gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(G1324gat));
  AND2_X1   g462(.A1(new_n660), .A2(new_n567), .ZN(new_n664));
  NAND2_X1  g463(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n239), .A2(new_n242), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT42), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n668), .ZN(new_n670));
  OAI211_X1 g469(.A(new_n669), .B(new_n670), .C1(new_n242), .C2(new_n664), .ZN(G1325gat));
  AOI21_X1  g470(.A(G15gat), .B1(new_n660), .B2(new_n603), .ZN(new_n672));
  INV_X1    g471(.A(new_n424), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n660), .A2(G15gat), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n672), .B1(new_n673), .B2(new_n674), .ZN(G1326gat));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n509), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT43), .B(G22gat), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(G1327gat));
  AND2_X1   g477(.A1(new_n608), .A2(new_n324), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n259), .A2(new_n260), .ZN(new_n680));
  INV_X1    g479(.A(new_n633), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n680), .A2(new_n681), .A3(new_n658), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n683), .A2(new_n276), .A3(new_n543), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT45), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n324), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(KEYINPUT102), .B1(new_n597), .B2(new_n607), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n416), .A2(new_n596), .A3(new_n591), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(KEYINPUT35), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT102), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n690), .A2(new_n691), .A3(new_n602), .A4(new_n606), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n688), .A2(new_n593), .A3(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT103), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n688), .A2(KEYINPUT103), .A3(new_n593), .A4(new_n692), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n687), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n679), .A2(new_n686), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n699), .A2(new_n543), .A3(new_n682), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n685), .B1(new_n701), .B2(new_n276), .ZN(G1328gat));
  NAND3_X1  g501(.A1(new_n699), .A2(new_n567), .A3(new_n682), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT104), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n699), .A2(KEYINPUT104), .A3(new_n567), .A4(new_n682), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n705), .A2(G36gat), .A3(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n683), .A2(new_n277), .A3(new_n567), .ZN(new_n708));
  XOR2_X1   g507(.A(new_n708), .B(KEYINPUT46), .Z(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n709), .ZN(G1329gat));
  OAI211_X1 g509(.A(new_n673), .B(new_n682), .C1(new_n697), .C2(new_n698), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(G43gat), .ZN(new_n712));
  INV_X1    g511(.A(G43gat), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n683), .A2(new_n713), .A3(new_n603), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT105), .ZN(new_n716));
  AOI21_X1  g515(.A(KEYINPUT47), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n715), .B(new_n717), .ZN(G1330gat));
  INV_X1    g517(.A(KEYINPUT106), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n699), .A2(new_n719), .A3(new_n509), .A4(new_n682), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n509), .B(new_n682), .C1(new_n697), .C2(new_n698), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(KEYINPUT106), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n720), .A2(G50gat), .A3(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(G50gat), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n683), .A2(new_n724), .A3(new_n509), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n725), .A2(KEYINPUT48), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n721), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n725), .B1(new_n728), .B2(new_n724), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT48), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n727), .A2(new_n731), .ZN(G1331gat));
  NAND2_X1  g531(.A1(new_n695), .A2(new_n696), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n658), .A2(new_n681), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n733), .A2(new_n325), .A3(new_n735), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n600), .B(KEYINPUT107), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(new_n206), .ZN(G1332gat));
  AND3_X1   g538(.A1(new_n733), .A2(new_n325), .A3(new_n735), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n567), .ZN(new_n741));
  OR2_X1    g540(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XOR2_X1   g542(.A(KEYINPUT49), .B(G64gat), .Z(new_n744));
  NOR2_X1   g543(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(KEYINPUT108), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n741), .A2(new_n742), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT108), .ZN(new_n748));
  OAI211_X1 g547(.A(new_n747), .B(new_n748), .C1(new_n741), .C2(new_n744), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n746), .A2(new_n749), .ZN(G1333gat));
  INV_X1    g549(.A(G71gat), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n740), .A2(new_n751), .A3(new_n603), .ZN(new_n752));
  OAI21_X1  g551(.A(G71gat), .B1(new_n736), .B2(new_n424), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT50), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n754), .B(new_n755), .ZN(G1334gat));
  NOR2_X1   g555(.A1(new_n736), .A2(new_n591), .ZN(new_n757));
  XNOR2_X1  g556(.A(KEYINPUT109), .B(G78gat), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n757), .B(new_n758), .ZN(G1335gat));
  NOR2_X1   g558(.A1(new_n680), .A2(new_n734), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n699), .A2(new_n760), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n761), .A2(new_n302), .A3(new_n600), .ZN(new_n762));
  INV_X1    g561(.A(new_n324), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n680), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n693), .A2(new_n681), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(KEYINPUT51), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT51), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n693), .A2(new_n767), .A3(new_n681), .A4(new_n764), .ZN(new_n768));
  AND2_X1   g567(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n769), .A2(new_n543), .A3(new_n658), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n762), .B1(new_n302), .B2(new_n770), .ZN(G1336gat));
  NAND4_X1  g570(.A1(new_n769), .A2(new_n303), .A3(new_n658), .A4(new_n567), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n567), .B(new_n760), .C1(new_n697), .C2(new_n698), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n772), .B1(new_n774), .B2(new_n303), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(KEYINPUT52), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT52), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n772), .B(new_n777), .C1(new_n774), .C2(new_n303), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(G1337gat));
  OAI21_X1  g578(.A(G99gat), .B1(new_n761), .B2(new_n424), .ZN(new_n780));
  INV_X1    g579(.A(G99gat), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n769), .A2(new_n781), .A3(new_n658), .A4(new_n603), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(G1338gat));
  INV_X1    g582(.A(KEYINPUT111), .ZN(new_n784));
  OR2_X1    g583(.A1(new_n784), .A2(KEYINPUT53), .ZN(new_n785));
  AND4_X1   g584(.A1(new_n498), .A2(new_n766), .A3(new_n658), .A4(new_n768), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n509), .B(new_n760), .C1(new_n697), .C2(new_n698), .ZN(new_n787));
  XOR2_X1   g586(.A(KEYINPUT110), .B(G106gat), .Z(new_n788));
  AOI22_X1  g587(.A1(new_n509), .A2(new_n786), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n784), .A2(KEYINPUT53), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n785), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n769), .A2(new_n498), .A3(new_n658), .A4(new_n509), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n787), .A2(new_n788), .ZN(new_n793));
  AND4_X1   g592(.A1(new_n785), .A2(new_n792), .A3(new_n793), .A4(new_n790), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n791), .A2(new_n794), .ZN(G1339gat));
  NAND2_X1  g594(.A1(new_n639), .A2(new_n645), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n647), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n639), .A2(new_n645), .A3(new_n638), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n797), .A2(KEYINPUT54), .A3(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n636), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n800), .B1(new_n646), .B2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n799), .A2(KEYINPUT55), .A3(new_n802), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n803), .A2(new_n655), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n799), .A2(new_n802), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n633), .A2(new_n804), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n619), .A2(new_n620), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n622), .A2(new_n610), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n809), .B1(new_n810), .B2(new_n612), .ZN(new_n811));
  INV_X1    g610(.A(new_n628), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n632), .B(new_n813), .C1(new_n653), .C2(new_n656), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n324), .B1(new_n808), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n324), .A2(new_n804), .A3(new_n807), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n813), .A2(new_n632), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n261), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n658), .A2(new_n633), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n680), .A2(new_n820), .A3(new_n763), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n822), .A2(new_n591), .A3(new_n603), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n543), .A2(new_n566), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(G113gat), .B1(new_n826), .B2(new_n681), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n737), .B1(new_n819), .B2(new_n821), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n595), .ZN(new_n829));
  OR3_X1    g628(.A1(new_n829), .A2(G113gat), .A3(new_n567), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n827), .B1(new_n830), .B2(new_n681), .ZN(G1340gat));
  OAI21_X1  g630(.A(G120gat), .B1(new_n826), .B2(new_n659), .ZN(new_n832));
  OR3_X1    g631(.A1(new_n829), .A2(G120gat), .A3(new_n567), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n832), .B1(new_n833), .B2(new_n659), .ZN(G1341gat));
  INV_X1    g633(.A(new_n829), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n835), .A2(new_n680), .A3(new_n566), .ZN(new_n836));
  INV_X1    g635(.A(G127gat), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n261), .A2(new_n837), .ZN(new_n838));
  AOI22_X1  g637(.A1(new_n836), .A2(new_n837), .B1(new_n825), .B2(new_n838), .ZN(G1342gat));
  INV_X1    g638(.A(G134gat), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n324), .A2(new_n566), .ZN(new_n841));
  XOR2_X1   g640(.A(new_n841), .B(KEYINPUT112), .Z(new_n842));
  NAND3_X1  g641(.A1(new_n835), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  XOR2_X1   g642(.A(new_n843), .B(KEYINPUT56), .Z(new_n844));
  OAI21_X1  g643(.A(G134gat), .B1(new_n826), .B2(new_n763), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(G1343gat));
  NOR2_X1   g645(.A1(new_n673), .A2(new_n591), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n828), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n848), .A2(new_n567), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n850), .A2(G141gat), .A3(new_n681), .ZN(new_n851));
  INV_X1    g650(.A(new_n821), .ZN(new_n852));
  INV_X1    g651(.A(new_n818), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n805), .A2(KEYINPUT113), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT114), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT113), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n799), .A2(new_n856), .A3(new_n802), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n854), .A2(new_n855), .A3(new_n806), .A4(new_n857), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n858), .A2(new_n633), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n803), .A2(new_n655), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n854), .A2(new_n806), .A3(new_n857), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n860), .B1(new_n861), .B2(KEYINPUT114), .ZN(new_n862));
  INV_X1    g661(.A(new_n817), .ZN(new_n863));
  AOI22_X1  g662(.A1(new_n859), .A2(new_n862), .B1(new_n658), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n853), .B1(new_n864), .B2(new_n324), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n852), .B1(new_n865), .B2(new_n261), .ZN(new_n866));
  OAI21_X1  g665(.A(KEYINPUT57), .B1(new_n866), .B2(new_n591), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n424), .A2(new_n543), .A3(new_n566), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n591), .B1(new_n819), .B2(new_n821), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT57), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n867), .A2(new_n633), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n851), .B1(G141gat), .B2(new_n872), .ZN(new_n873));
  XOR2_X1   g672(.A(KEYINPUT116), .B(KEYINPUT58), .Z(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT115), .ZN(new_n876));
  AND3_X1   g675(.A1(new_n799), .A2(new_n856), .A3(new_n802), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n856), .B1(new_n799), .B2(new_n802), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n877), .A2(new_n878), .A3(KEYINPUT55), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n804), .B1(new_n879), .B2(new_n855), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n858), .A2(new_n633), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n814), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n818), .B1(new_n882), .B2(new_n763), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n821), .B1(new_n883), .B2(new_n680), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n870), .B1(new_n884), .B2(new_n509), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n886));
  INV_X1    g685(.A(new_n868), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n876), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n862), .A2(new_n633), .A3(new_n858), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n324), .B1(new_n890), .B2(new_n814), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n261), .B1(new_n891), .B2(new_n818), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n591), .B1(new_n892), .B2(new_n821), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n871), .B(KEYINPUT115), .C1(new_n893), .C2(new_n870), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n889), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(new_n633), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n851), .B1(new_n896), .B2(G141gat), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT58), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n875), .B1(new_n897), .B2(new_n898), .ZN(G1344gat));
  XNOR2_X1  g698(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n816), .B(KEYINPUT119), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n891), .B1(new_n863), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n821), .B1(new_n903), .B2(new_n680), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n904), .A2(new_n870), .A3(new_n509), .ZN(new_n905));
  OR2_X1    g704(.A1(new_n869), .A2(new_n870), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n905), .A2(new_n658), .A3(new_n887), .A4(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n901), .B1(new_n907), .B2(G148gat), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT117), .ZN(new_n910));
  INV_X1    g709(.A(new_n894), .ZN(new_n911));
  AOI21_X1  g710(.A(KEYINPUT115), .B1(new_n867), .B2(new_n871), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n658), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(G148gat), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n914), .A2(KEYINPUT59), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n910), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n659), .B1(new_n889), .B2(new_n894), .ZN(new_n917));
  INV_X1    g716(.A(new_n915), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n917), .A2(KEYINPUT117), .A3(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n909), .B1(new_n916), .B2(new_n919), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n850), .A2(G148gat), .A3(new_n659), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n920), .A2(KEYINPUT120), .A3(new_n922), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT120), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n913), .A2(new_n910), .A3(new_n915), .ZN(new_n925));
  OAI21_X1  g724(.A(KEYINPUT117), .B1(new_n917), .B2(new_n918), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n908), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n924), .B1(new_n927), .B2(new_n921), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n923), .A2(new_n928), .ZN(G1345gat));
  AOI21_X1  g728(.A(G155gat), .B1(new_n849), .B2(new_n680), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n680), .A2(G155gat), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(KEYINPUT121), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n930), .B1(new_n895), .B2(new_n932), .ZN(G1346gat));
  AOI21_X1  g732(.A(new_n763), .B1(new_n889), .B2(new_n894), .ZN(new_n934));
  INV_X1    g733(.A(G162gat), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n842), .A2(new_n935), .ZN(new_n936));
  OAI22_X1  g735(.A1(new_n934), .A2(new_n935), .B1(new_n848), .B2(new_n936), .ZN(G1347gat));
  NAND2_X1  g736(.A1(new_n737), .A2(new_n567), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n823), .A2(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(new_n939), .ZN(new_n940));
  OAI21_X1  g739(.A(G169gat), .B1(new_n940), .B2(new_n681), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n543), .B1(new_n819), .B2(new_n821), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n942), .A2(new_n567), .A3(new_n595), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n633), .B1(new_n328), .B2(new_n327), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n941), .B1(new_n943), .B2(new_n944), .ZN(G1348gat));
  NAND3_X1  g744(.A1(new_n939), .A2(G176gat), .A3(new_n658), .ZN(new_n946));
  XOR2_X1   g745(.A(new_n946), .B(KEYINPUT122), .Z(new_n947));
  INV_X1    g746(.A(new_n943), .ZN(new_n948));
  AOI21_X1  g747(.A(G176gat), .B1(new_n948), .B2(new_n658), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n947), .A2(new_n949), .ZN(G1349gat));
  OAI21_X1  g749(.A(new_n347), .B1(new_n940), .B2(new_n261), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n948), .A2(new_n680), .A3(new_n358), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT60), .ZN(new_n953));
  AOI22_X1  g752(.A1(new_n951), .A2(new_n952), .B1(KEYINPUT123), .B2(new_n953), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n953), .A2(KEYINPUT123), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n954), .B(new_n955), .ZN(G1350gat));
  AOI21_X1  g755(.A(new_n334), .B1(new_n939), .B2(new_n324), .ZN(new_n957));
  XOR2_X1   g756(.A(new_n957), .B(KEYINPUT61), .Z(new_n958));
  NAND3_X1  g757(.A1(new_n948), .A2(new_n334), .A3(new_n324), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(G1351gat));
  NAND3_X1  g759(.A1(new_n847), .A2(new_n567), .A3(new_n942), .ZN(new_n961));
  NOR3_X1   g760(.A1(new_n961), .A2(G197gat), .A3(new_n681), .ZN(new_n962));
  XOR2_X1   g761(.A(new_n962), .B(KEYINPUT124), .Z(new_n963));
  NOR2_X1   g762(.A1(new_n673), .A2(new_n938), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n905), .A2(new_n906), .A3(new_n964), .ZN(new_n965));
  OAI21_X1  g764(.A(G197gat), .B1(new_n965), .B2(new_n681), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n963), .A2(new_n966), .ZN(G1352gat));
  AND3_X1   g766(.A1(new_n905), .A2(new_n658), .A3(new_n906), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n443), .B1(new_n968), .B2(new_n964), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n961), .A2(G204gat), .A3(new_n659), .ZN(new_n970));
  XOR2_X1   g769(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n971));
  XNOR2_X1  g770(.A(new_n970), .B(new_n971), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n969), .A2(new_n972), .ZN(new_n973));
  XOR2_X1   g772(.A(new_n973), .B(KEYINPUT126), .Z(G1353gat));
  OR3_X1    g773(.A1(new_n961), .A2(new_n261), .A3(new_n458), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n965), .A2(new_n261), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n976), .A2(new_n451), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(KEYINPUT63), .ZN(new_n978));
  INV_X1    g777(.A(new_n978), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n977), .A2(KEYINPUT63), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n975), .B1(new_n979), .B2(new_n980), .ZN(G1354gat));
  NOR3_X1   g780(.A1(new_n965), .A2(new_n441), .A3(new_n763), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n441), .B1(new_n961), .B2(new_n763), .ZN(new_n983));
  XNOR2_X1  g782(.A(new_n983), .B(KEYINPUT127), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n982), .A2(new_n984), .ZN(G1355gat));
endmodule


