//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 0 1 0 1 1 0 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 0 0 1 0 1 0 1 1 1 1 1 0 1 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:11 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1198, new_n1199, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G50), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT64), .Z(new_n205));
  INV_X1    g0005(.A(G77), .ZN(new_n206));
  AND2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0008(.A(G250), .ZN(new_n209));
  INV_X1    g0009(.A(KEYINPUT65), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  OAI21_X1  g0011(.A(new_n210), .B1(new_n211), .B2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(G13), .ZN(new_n213));
  NAND4_X1  g0013(.A1(new_n213), .A2(KEYINPUT65), .A3(G1), .A4(G20), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G257), .ZN(new_n217));
  INV_X1    g0017(.A(G264), .ZN(new_n218));
  AOI211_X1 g0018(.A(new_n209), .B(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  INV_X1    g0020(.A(G20), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n203), .A2(G50), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(new_n219), .A2(KEYINPUT0), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n225), .B1(KEYINPUT0), .B2(new_n219), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n227));
  INV_X1    g0027(.A(G244), .ZN(new_n228));
  INV_X1    g0028(.A(G107), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n227), .B1(new_n206), .B2(new_n228), .C1(new_n229), .C2(new_n218), .ZN(new_n230));
  AOI22_X1  g0030(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  INV_X1    g0032(.A(G97), .ZN(new_n233));
  OAI221_X1 g0033(.A(new_n231), .B1(new_n201), .B2(new_n232), .C1(new_n233), .C2(new_n217), .ZN(new_n234));
  OAI21_X1  g0034(.A(new_n211), .B1(new_n230), .B2(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT1), .ZN(new_n236));
  NOR2_X1   g0036(.A1(new_n226), .A2(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(new_n232), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT2), .B(G226), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G264), .B(G270), .Z(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XOR2_X1   g0047(.A(new_n246), .B(new_n247), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT66), .ZN(new_n249));
  XOR2_X1   g0049(.A(G68), .B(G77), .Z(new_n250));
  XNOR2_X1  g0050(.A(G50), .B(G58), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n250), .B(new_n251), .Z(new_n252));
  XOR2_X1   g0052(.A(new_n249), .B(new_n252), .Z(G351));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n220), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n205), .A2(new_n221), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n201), .A2(KEYINPUT8), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT8), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G58), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(G20), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G150), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G20), .A2(G33), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  OAI22_X1  g0067(.A1(new_n261), .A2(new_n264), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n255), .B1(new_n256), .B2(new_n268), .ZN(new_n269));
  NOR3_X1   g0069(.A1(new_n213), .A2(new_n221), .A3(G1), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n270), .A2(new_n255), .ZN(new_n271));
  INV_X1    g0071(.A(G50), .ZN(new_n272));
  INV_X1    g0072(.A(G1), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n272), .B1(new_n273), .B2(G20), .ZN(new_n274));
  AOI22_X1  g0074(.A1(new_n271), .A2(new_n274), .B1(new_n272), .B2(new_n270), .ZN(new_n275));
  AND3_X1   g0075(.A1(new_n269), .A2(KEYINPUT9), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(KEYINPUT9), .B1(new_n269), .B2(new_n275), .ZN(new_n277));
  INV_X1    g0077(.A(G41), .ZN(new_n278));
  OAI211_X1 g0078(.A(G1), .B(G13), .C1(new_n262), .C2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G45), .ZN(new_n280));
  AOI21_X1  g0080(.A(G1), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n279), .A2(G274), .A3(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n273), .B1(G41), .B2(G45), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n279), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n283), .B1(G226), .B2(new_n286), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT3), .B(G33), .ZN(new_n288));
  NOR2_X1   g0088(.A1(G222), .A2(G1698), .ZN(new_n289));
  INV_X1    g0089(.A(G1698), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n290), .A2(G223), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n288), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n220), .B1(G33), .B2(G41), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n292), .B(new_n293), .C1(G77), .C2(new_n288), .ZN(new_n294));
  AND2_X1   g0094(.A1(new_n287), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G190), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NOR3_X1   g0098(.A1(new_n276), .A2(new_n277), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(KEYINPUT67), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT10), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n296), .A2(G200), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n299), .A2(new_n303), .ZN(new_n304));
  XOR2_X1   g0104(.A(new_n302), .B(new_n304), .Z(new_n305));
  NAND2_X1  g0105(.A1(new_n269), .A2(new_n275), .ZN(new_n306));
  INV_X1    g0106(.A(G179), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n295), .A2(new_n307), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n306), .B(new_n308), .C1(G169), .C2(new_n295), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n305), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G226), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n290), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n232), .A2(G1698), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n288), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(G33), .A2(G97), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n279), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G238), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n282), .B1(new_n285), .B2(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(KEYINPUT13), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  NOR3_X1   g0121(.A1(new_n317), .A2(new_n319), .A3(KEYINPUT13), .ZN(new_n322));
  NOR3_X1   g0122(.A1(new_n321), .A2(new_n322), .A3(new_n307), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT69), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n320), .A2(new_n325), .ZN(new_n326));
  OAI211_X1 g0126(.A(KEYINPUT69), .B(KEYINPUT13), .C1(new_n317), .C2(new_n319), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n317), .A2(new_n319), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT13), .ZN(new_n329));
  AOI21_X1  g0129(.A(KEYINPUT68), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT68), .ZN(new_n331));
  NOR4_X1   g0131(.A1(new_n317), .A2(new_n319), .A3(new_n331), .A4(KEYINPUT13), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n326), .B(new_n327), .C1(new_n330), .C2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n333), .A2(KEYINPUT14), .A3(G169), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(KEYINPUT14), .B1(new_n333), .B2(G169), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n324), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n266), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n338), .B1(new_n264), .B2(new_n206), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n255), .ZN(new_n340));
  XOR2_X1   g0140(.A(new_n340), .B(KEYINPUT11), .Z(new_n341));
  NAND2_X1  g0141(.A1(new_n270), .A2(new_n202), .ZN(new_n342));
  XNOR2_X1  g0142(.A(new_n342), .B(KEYINPUT12), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n273), .A2(G20), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n271), .A2(G68), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n341), .B1(KEYINPUT70), .B2(new_n346), .ZN(new_n347));
  OR2_X1    g0147(.A1(new_n346), .A2(KEYINPUT70), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n337), .A2(new_n349), .ZN(new_n350));
  NOR3_X1   g0150(.A1(new_n321), .A2(new_n322), .A3(new_n297), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n333), .A2(G200), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n271), .A2(G77), .A3(new_n344), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n213), .A2(G1), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(G20), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n355), .B1(G77), .B2(new_n357), .ZN(new_n358));
  AND2_X1   g0158(.A1(new_n254), .A2(new_n220), .ZN(new_n359));
  XOR2_X1   g0159(.A(KEYINPUT15), .B(G87), .Z(new_n360));
  AOI22_X1  g0160(.A1(new_n360), .A2(new_n263), .B1(G20), .B2(G77), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n260), .A2(new_n266), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n359), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n358), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n288), .A2(G238), .A3(G1698), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n365), .B1(new_n229), .B2(new_n288), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT3), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(G33), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  NOR3_X1   g0170(.A1(new_n370), .A2(new_n232), .A3(G1698), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n293), .B1(new_n366), .B2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n283), .B1(G244), .B2(new_n286), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(G169), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n364), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n376), .B1(G179), .B2(new_n374), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n374), .A2(G200), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n378), .B(new_n364), .C1(new_n297), .C2(new_n374), .ZN(new_n379));
  AND3_X1   g0179(.A1(new_n354), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  AND3_X1   g0180(.A1(new_n311), .A2(new_n350), .A3(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT74), .ZN(new_n382));
  NAND2_X1  g0182(.A1(G58), .A2(G68), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n203), .A2(new_n383), .ZN(new_n384));
  AOI22_X1  g0184(.A1(new_n384), .A2(G20), .B1(G159), .B2(new_n266), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  XNOR2_X1  g0186(.A(KEYINPUT71), .B(KEYINPUT3), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n369), .B1(new_n387), .B2(G33), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT7), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n389), .A2(G20), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT72), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n368), .A2(G33), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n221), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n392), .B1(new_n395), .B2(new_n389), .ZN(new_n396));
  AOI21_X1  g0196(.A(G20), .B1(new_n367), .B2(new_n369), .ZN(new_n397));
  NOR3_X1   g0197(.A1(new_n397), .A2(KEYINPUT72), .A3(KEYINPUT7), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n391), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(G68), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n386), .B1(new_n400), .B2(KEYINPUT73), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT73), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n399), .A2(new_n402), .A3(G68), .ZN(new_n403));
  AOI21_X1  g0203(.A(KEYINPUT16), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n368), .A2(KEYINPUT71), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT71), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(KEYINPUT3), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n405), .A2(new_n407), .A3(G33), .ZN(new_n408));
  AOI21_X1  g0208(.A(G20), .B1(new_n408), .B2(new_n367), .ZN(new_n409));
  OAI21_X1  g0209(.A(G68), .B1(new_n409), .B2(new_n389), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n393), .B1(new_n387), .B2(G33), .ZN(new_n411));
  NOR3_X1   g0211(.A1(new_n411), .A2(KEYINPUT7), .A3(G20), .ZN(new_n412));
  OAI211_X1 g0212(.A(KEYINPUT16), .B(new_n385), .C1(new_n410), .C2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n255), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n382), .B1(new_n404), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(KEYINPUT72), .B1(new_n397), .B2(KEYINPUT7), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n392), .B(new_n389), .C1(new_n288), .C2(G20), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n416), .A2(new_n417), .B1(new_n388), .B2(new_n390), .ZN(new_n418));
  OAI21_X1  g0218(.A(KEYINPUT73), .B1(new_n418), .B2(new_n202), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n403), .A2(new_n419), .A3(new_n385), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT16), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n414), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(KEYINPUT74), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n359), .A2(new_n357), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n260), .A2(new_n344), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n424), .B1(KEYINPUT75), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(KEYINPUT75), .B2(new_n425), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n261), .A2(new_n270), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  XNOR2_X1  g0229(.A(new_n429), .B(KEYINPUT76), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n408), .A2(new_n367), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n312), .A2(G1698), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n432), .B1(G223), .B2(G1698), .ZN(new_n433));
  INV_X1    g0233(.A(G87), .ZN(new_n434));
  OAI22_X1  g0234(.A1(new_n431), .A2(new_n433), .B1(new_n262), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n293), .ZN(new_n436));
  XNOR2_X1  g0236(.A(new_n436), .B(KEYINPUT77), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n282), .B1(new_n285), .B2(new_n232), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n438), .A2(G190), .ZN(new_n439));
  INV_X1    g0239(.A(G200), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n438), .B1(new_n435), .B2(new_n293), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n437), .A2(new_n439), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n415), .A2(new_n423), .A3(new_n430), .A4(new_n444), .ZN(new_n445));
  XNOR2_X1  g0245(.A(KEYINPUT78), .B(KEYINPUT17), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT79), .ZN(new_n449));
  AND2_X1   g0249(.A1(new_n427), .A2(new_n428), .ZN(new_n450));
  XNOR2_X1  g0250(.A(new_n450), .B(KEYINPUT76), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n420), .A2(new_n421), .ZN(new_n452));
  INV_X1    g0252(.A(new_n414), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n451), .B1(new_n382), .B2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT17), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n456), .A2(KEYINPUT78), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n455), .A2(new_n423), .A3(new_n444), .A4(new_n458), .ZN(new_n459));
  AND3_X1   g0259(.A1(new_n448), .A2(new_n449), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n449), .B1(new_n448), .B2(new_n459), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n438), .A2(G179), .ZN(new_n462));
  AOI22_X1  g0262(.A1(new_n437), .A2(new_n462), .B1(new_n375), .B2(new_n442), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n430), .B1(new_n422), .B2(KEYINPUT74), .ZN(new_n464));
  AOI211_X1 g0264(.A(new_n382), .B(new_n414), .C1(new_n420), .C2(new_n421), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT18), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT18), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n468), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NOR3_X1   g0270(.A1(new_n460), .A2(new_n461), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n381), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n273), .A2(G33), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n271), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(G116), .ZN(new_n476));
  OAI21_X1  g0276(.A(KEYINPUT84), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT84), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n271), .A2(new_n478), .A3(G116), .A4(new_n474), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(G33), .A2(G283), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n481), .B(new_n221), .C1(G33), .C2(new_n233), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n221), .A2(G116), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n482), .A2(new_n484), .A3(new_n255), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT20), .ZN(new_n486));
  OR2_X1    g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n486), .ZN(new_n488));
  AOI22_X1  g0288(.A1(new_n487), .A2(new_n488), .B1(new_n356), .B2(new_n483), .ZN(new_n489));
  XNOR2_X1  g0289(.A(KEYINPUT5), .B(G41), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n280), .A2(G1), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n279), .A2(G274), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(G270), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n492), .A2(new_n279), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(G257), .A2(G1698), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n499), .B1(new_n218), .B2(G1698), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n500), .A2(new_n408), .A3(new_n367), .ZN(new_n501));
  INV_X1    g0301(.A(G303), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n501), .B1(new_n502), .B2(new_n288), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n279), .B1(new_n503), .B2(KEYINPUT83), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT83), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n501), .B(new_n505), .C1(new_n502), .C2(new_n288), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n498), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n480), .B(new_n489), .C1(new_n507), .C2(new_n440), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n508), .B1(G190), .B2(new_n507), .ZN(new_n509));
  NOR2_X1   g0309(.A1(KEYINPUT85), .A2(KEYINPUT21), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n489), .A2(new_n480), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(G169), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n510), .B1(new_n512), .B2(new_n507), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n504), .A2(new_n506), .ZN(new_n514));
  INV_X1    g0314(.A(new_n498), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n510), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n516), .A2(G169), .A3(new_n517), .A4(new_n511), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n507), .A2(new_n511), .A3(G179), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n513), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n509), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n270), .A2(KEYINPUT25), .A3(new_n229), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(KEYINPUT25), .B1(new_n270), .B2(new_n229), .ZN(new_n524));
  OAI22_X1  g0324(.A1(new_n475), .A2(new_n229), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n221), .A2(G87), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT22), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n408), .A2(new_n529), .A3(new_n367), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n528), .B1(new_n370), .B2(new_n527), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT23), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n532), .B1(new_n221), .B2(G107), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n229), .A2(KEYINPUT23), .A3(G20), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n262), .A2(new_n476), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n533), .A2(new_n534), .B1(new_n535), .B2(new_n221), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n530), .A2(new_n531), .A3(new_n536), .ZN(new_n537));
  OR2_X1    g0337(.A1(new_n537), .A2(KEYINPUT86), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(KEYINPUT86), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n538), .A2(KEYINPUT24), .A3(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n255), .B1(new_n539), .B2(KEYINPUT24), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n526), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(KEYINPUT87), .B1(new_n497), .B2(new_n218), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n293), .B1(new_n491), .B2(new_n490), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT87), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n545), .A2(new_n546), .A3(G264), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n217), .A2(G1698), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(G250), .B2(G1698), .ZN(new_n550));
  INV_X1    g0350(.A(G294), .ZN(new_n551));
  OAI22_X1  g0351(.A1(new_n431), .A2(new_n550), .B1(new_n262), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n293), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n548), .A2(new_n495), .A3(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n554), .A2(KEYINPUT88), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT88), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n544), .A2(new_n547), .B1(new_n552), .B2(new_n293), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n556), .B1(new_n557), .B2(new_n495), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n297), .B1(new_n555), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n554), .A2(new_n440), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n543), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n542), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n525), .B1(new_n562), .B2(new_n540), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n554), .A2(KEYINPUT88), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n557), .A2(new_n556), .A3(new_n495), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n564), .A2(G169), .A3(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n557), .A2(G179), .A3(new_n495), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n563), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n561), .A2(new_n568), .ZN(new_n569));
  NOR3_X1   g0369(.A1(new_n293), .A2(new_n209), .A3(new_n491), .ZN(new_n570));
  INV_X1    g0370(.A(new_n491), .ZN(new_n571));
  OAI21_X1  g0371(.A(KEYINPUT80), .B1(new_n493), .B2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT80), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n279), .A2(new_n573), .A3(G274), .A4(new_n491), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n570), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(G238), .A2(G1698), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n576), .B1(new_n228), .B2(G1698), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n577), .A2(new_n408), .A3(new_n367), .ZN(new_n578));
  INV_X1    g0378(.A(new_n535), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n293), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n575), .A2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT81), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n575), .A2(new_n581), .A3(KEYINPUT81), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n584), .A2(new_n307), .A3(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n360), .A2(new_n357), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT19), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n263), .A2(new_n588), .A3(G97), .ZN(new_n589));
  NOR2_X1   g0389(.A1(G97), .A2(G107), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n590), .A2(new_n434), .B1(new_n316), .B2(new_n221), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n589), .B1(new_n591), .B2(new_n588), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n221), .A2(G68), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n592), .B1(new_n431), .B2(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n587), .B1(new_n594), .B2(new_n255), .ZN(new_n595));
  XNOR2_X1  g0395(.A(new_n360), .B(KEYINPUT82), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n595), .B1(new_n475), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n586), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(G169), .B1(new_n584), .B2(new_n585), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n584), .A2(G190), .A3(new_n585), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n271), .A2(G87), .A3(new_n474), .ZN(new_n601));
  AND2_X1   g0401(.A1(new_n595), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n440), .B1(new_n584), .B2(new_n585), .ZN(new_n604));
  OAI22_X1  g0404(.A1(new_n598), .A2(new_n599), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n494), .B1(G257), .B2(new_n545), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n288), .A2(G250), .A3(G1698), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT4), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n608), .A2(new_n228), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n288), .A2(new_n290), .A3(new_n609), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n607), .A2(new_n610), .A3(new_n481), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n290), .A2(G244), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n608), .B1(new_n431), .B2(new_n612), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  OAI211_X1 g0414(.A(G190), .B(new_n606), .C1(new_n614), .C2(new_n279), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n229), .A2(KEYINPUT6), .A3(G97), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n233), .A2(new_n229), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n617), .A2(new_n590), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n616), .B1(new_n618), .B2(KEYINPUT6), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n619), .A2(G20), .B1(G77), .B2(new_n266), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n620), .B1(new_n418), .B2(new_n229), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n255), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n279), .B1(new_n611), .B2(new_n613), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n495), .B1(new_n217), .B2(new_n497), .ZN(new_n624));
  OAI21_X1  g0424(.A(G200), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  MUX2_X1   g0425(.A(new_n357), .B(new_n475), .S(G97), .Z(new_n626));
  NAND4_X1  g0426(.A1(new_n615), .A2(new_n622), .A3(new_n625), .A4(new_n626), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n622), .A2(new_n626), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n375), .B1(new_n623), .B2(new_n624), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n606), .B1(new_n614), .B2(new_n279), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n629), .B1(new_n630), .B2(G179), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n627), .B1(new_n628), .B2(new_n631), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n605), .A2(new_n632), .ZN(new_n633));
  AND4_X1   g0433(.A1(new_n473), .A2(new_n521), .A3(new_n569), .A4(new_n633), .ZN(G372));
  NAND2_X1  g0434(.A1(new_n448), .A2(new_n459), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(KEYINPUT79), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n448), .A2(new_n459), .A3(new_n449), .ZN(new_n637));
  INV_X1    g0437(.A(new_n354), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n350), .B1(new_n638), .B2(new_n377), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n636), .A2(new_n637), .A3(new_n639), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n467), .A2(new_n469), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n305), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n642), .A2(new_n310), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n643), .A2(KEYINPUT92), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT92), .ZN(new_n645));
  NOR3_X1   g0445(.A1(new_n642), .A2(new_n645), .A3(new_n310), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n628), .A2(new_n631), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT26), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n605), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT91), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n582), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n586), .B(new_n597), .C1(G169), .C2(new_n655), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n600), .B(new_n602), .C1(new_n440), .C2(new_n655), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n649), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n651), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n654), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n657), .A2(new_n656), .ZN(new_n661));
  OR3_X1    g0461(.A1(new_n561), .A2(new_n661), .A3(new_n632), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n520), .A2(KEYINPUT89), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT89), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n513), .A2(new_n518), .A3(new_n664), .A4(new_n519), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n568), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(KEYINPUT90), .B1(new_n662), .B2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT90), .ZN(new_n668));
  NOR3_X1   g0468(.A1(new_n561), .A2(new_n661), .A3(new_n632), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n663), .A2(new_n665), .ZN(new_n670));
  OAI211_X1 g0470(.A(new_n668), .B(new_n669), .C1(new_n670), .C2(new_n568), .ZN(new_n671));
  INV_X1    g0471(.A(new_n656), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n672), .B1(new_n652), .B2(new_n653), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n660), .A2(new_n667), .A3(new_n671), .A4(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n473), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n648), .A2(new_n675), .ZN(G369));
  NAND2_X1  g0476(.A1(new_n356), .A2(new_n221), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n678), .B(KEYINPUT93), .ZN(new_n679));
  OAI21_X1  g0479(.A(G213), .B1(new_n677), .B2(KEYINPUT27), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(G343), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(new_n511), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n684), .B(KEYINPUT94), .ZN(new_n685));
  MUX2_X1   g0485(.A(new_n670), .B(new_n521), .S(new_n685), .Z(new_n686));
  AND2_X1   g0486(.A1(new_n686), .A2(G330), .ZN(new_n687));
  INV_X1    g0487(.A(new_n683), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n569), .B1(new_n563), .B2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n568), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n689), .B1(new_n690), .B2(new_n688), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n687), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n520), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(new_n683), .ZN(new_n695));
  AOI22_X1  g0495(.A1(new_n695), .A2(new_n569), .B1(new_n568), .B2(new_n688), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n693), .A2(new_n696), .ZN(G399));
  NOR2_X1   g0497(.A1(new_n216), .A2(G41), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n590), .A2(new_n434), .A3(new_n476), .ZN(new_n699));
  NOR3_X1   g0499(.A1(new_n698), .A2(new_n273), .A3(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n700), .B1(new_n224), .B2(new_n698), .ZN(new_n701));
  XOR2_X1   g0501(.A(new_n701), .B(KEYINPUT28), .Z(new_n702));
  OAI21_X1  g0502(.A(new_n669), .B1(new_n520), .B2(new_n568), .ZN(new_n703));
  OR3_X1    g0503(.A1(new_n605), .A2(new_n650), .A3(KEYINPUT26), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n672), .B1(new_n658), .B2(KEYINPUT26), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n703), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  AND3_X1   g0506(.A1(new_n706), .A2(KEYINPUT29), .A3(new_n688), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n674), .A2(new_n688), .ZN(new_n708));
  XOR2_X1   g0508(.A(KEYINPUT97), .B(KEYINPUT29), .Z(new_n709));
  AOI21_X1  g0509(.A(new_n707), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(G330), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n633), .A2(new_n569), .A3(new_n521), .A4(new_n688), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(KEYINPUT31), .ZN(new_n713));
  NOR3_X1   g0513(.A1(new_n516), .A2(new_n630), .A3(new_n307), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n584), .A2(new_n557), .A3(new_n585), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(KEYINPUT95), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT95), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n584), .A2(new_n585), .A3(new_n717), .A4(new_n557), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n714), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT30), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n714), .A2(new_n716), .A3(KEYINPUT30), .A4(new_n718), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n655), .A2(G179), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n723), .A2(new_n554), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n724), .A2(KEYINPUT96), .A3(new_n516), .A4(new_n630), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT96), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n723), .A2(new_n554), .A3(new_n630), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n726), .B1(new_n727), .B2(new_n507), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n721), .A2(new_n722), .A3(new_n725), .A4(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(new_n683), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n713), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT31), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n727), .A2(new_n507), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n733), .B1(new_n719), .B2(new_n720), .ZN(new_n734));
  AOI211_X1 g0534(.A(new_n732), .B(new_n688), .C1(new_n734), .C2(new_n722), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n711), .B1(new_n731), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n710), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n702), .B1(new_n738), .B2(G1), .ZN(G364));
  NOR2_X1   g0539(.A1(new_n686), .A2(G330), .ZN(new_n740));
  INV_X1    g0540(.A(new_n698), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n213), .A2(G20), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n273), .B1(new_n742), .B2(G45), .ZN(new_n743));
  AOI211_X1 g0543(.A(new_n740), .B(new_n687), .C1(new_n741), .C2(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n220), .B1(G20), .B2(new_n375), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n297), .A2(G179), .A3(G200), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(new_n221), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n221), .A2(G179), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G190), .A2(G200), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g0552(.A(KEYINPUT99), .B(G159), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT32), .ZN(new_n755));
  AOI22_X1  g0555(.A1(G97), .A2(new_n749), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n221), .A2(new_n307), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G200), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n297), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n750), .A2(new_n297), .A3(G200), .ZN(new_n761));
  OAI221_X1 g0561(.A(new_n756), .B1(new_n272), .B2(new_n760), .C1(new_n229), .C2(new_n761), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n750), .A2(G190), .A3(G200), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G87), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n758), .A2(G190), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  OAI221_X1 g0567(.A(new_n765), .B1(new_n755), .B2(new_n754), .C1(new_n767), .C2(new_n202), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n757), .A2(new_n751), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n757), .A2(G190), .A3(new_n440), .ZN(new_n770));
  OAI221_X1 g0570(.A(new_n288), .B1(new_n769), .B2(new_n206), .C1(new_n201), .C2(new_n770), .ZN(new_n771));
  OR3_X1    g0571(.A1(new_n762), .A2(new_n768), .A3(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G322), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(G311), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n370), .B1(new_n769), .B2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n752), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n774), .B(new_n776), .C1(G329), .C2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n764), .A2(G303), .ZN(new_n779));
  XNOR2_X1  g0579(.A(KEYINPUT33), .B(G317), .ZN(new_n780));
  INV_X1    g0580(.A(new_n761), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n766), .A2(new_n780), .B1(new_n781), .B2(G283), .ZN(new_n782));
  AOI22_X1  g0582(.A1(G294), .A2(new_n749), .B1(new_n759), .B2(G326), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n778), .A2(new_n779), .A3(new_n782), .A4(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n746), .B1(new_n772), .B2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n743), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n698), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n216), .A2(new_n411), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n790), .B1(new_n280), .B2(new_n224), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n792), .A2(KEYINPUT98), .B1(G45), .B2(new_n252), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n793), .B1(KEYINPUT98), .B2(new_n792), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n216), .A2(new_n370), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n795), .A2(G355), .B1(new_n476), .B2(new_n216), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(G13), .A2(G33), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(G20), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(new_n745), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n785), .B(new_n788), .C1(new_n797), .C2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n800), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n802), .B1(new_n686), .B2(new_n803), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT100), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n744), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(G396));
  OAI21_X1  g0607(.A(new_n379), .B1(new_n688), .B2(new_n364), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(new_n377), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n377), .A2(new_n683), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n708), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n674), .A2(new_n688), .A3(new_n812), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n737), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(new_n787), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n814), .A2(new_n737), .A3(new_n815), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n745), .A2(new_n798), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n788), .B1(new_n206), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n769), .ZN(new_n822));
  AOI22_X1  g0622(.A1(G116), .A2(new_n822), .B1(new_n777), .B2(G311), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n823), .B(new_n370), .C1(new_n551), .C2(new_n770), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n759), .A2(G303), .B1(new_n781), .B2(G87), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(new_n229), .B2(new_n763), .ZN(new_n826));
  INV_X1    g0626(.A(G283), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n767), .A2(new_n827), .B1(new_n233), .B2(new_n748), .ZN(new_n828));
  NOR3_X1   g0628(.A1(new_n824), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n770), .ZN(new_n830));
  INV_X1    g0630(.A(new_n753), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n830), .A2(G143), .B1(new_n822), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(G137), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n832), .B1(new_n767), .B2(new_n265), .C1(new_n833), .C2(new_n760), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n834), .B(KEYINPUT34), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n781), .A2(G68), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n836), .B1(new_n272), .B2(new_n763), .C1(new_n201), .C2(new_n748), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n431), .B(new_n837), .C1(G132), .C2(new_n777), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n829), .B1(new_n835), .B2(new_n838), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n821), .B1(new_n746), .B2(new_n839), .C1(new_n812), .C2(new_n799), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n819), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(G384));
  OR2_X1    g0642(.A1(new_n619), .A2(KEYINPUT35), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n619), .A2(KEYINPUT35), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n843), .A2(G116), .A3(new_n222), .A4(new_n844), .ZN(new_n845));
  XOR2_X1   g0645(.A(new_n845), .B(KEYINPUT36), .Z(new_n846));
  NAND3_X1  g0646(.A1(new_n224), .A2(G77), .A3(new_n383), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n272), .A2(G68), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n273), .B(G13), .C1(new_n847), .C2(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  NOR3_X1   g0650(.A1(new_n464), .A2(new_n465), .A3(new_n443), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n385), .B1(new_n410), .B2(new_n412), .ZN(new_n852));
  AND2_X1   g0652(.A1(new_n852), .A2(new_n421), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n450), .B1(new_n853), .B2(new_n414), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n463), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n681), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(KEYINPUT37), .B1(new_n851), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n856), .B1(new_n464), .B2(new_n465), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT37), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n466), .A2(new_n860), .A3(new_n445), .A4(new_n861), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  OAI211_X1 g0664(.A(KEYINPUT38), .B(new_n864), .C1(new_n471), .C2(new_n857), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT106), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n636), .A2(new_n641), .A3(new_n637), .ZN(new_n868));
  INV_X1    g0668(.A(new_n857), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n870), .A2(KEYINPUT106), .A3(KEYINPUT38), .A4(new_n864), .ZN(new_n871));
  XNOR2_X1  g0671(.A(KEYINPUT105), .B(KEYINPUT39), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n466), .A2(new_n860), .A3(new_n445), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(KEYINPUT37), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n862), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n470), .B1(new_n448), .B2(new_n459), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n875), .B1(new_n876), .B2(new_n860), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT38), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n872), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n867), .A2(new_n871), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(KEYINPUT107), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT107), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n867), .A2(new_n879), .A3(new_n882), .A4(new_n871), .ZN(new_n883));
  AOI21_X1  g0683(.A(KEYINPUT38), .B1(new_n870), .B2(new_n864), .ZN(new_n884));
  AOI211_X1 g0684(.A(new_n878), .B(new_n863), .C1(new_n868), .C2(new_n869), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT39), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n881), .A2(new_n883), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n333), .A2(G169), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT14), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n323), .B1(new_n890), .B2(new_n334), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n347), .A2(new_n348), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT102), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT102), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n337), .A2(new_n894), .A3(new_n349), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n688), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n887), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n470), .A2(new_n681), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n884), .A2(new_n885), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT104), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n811), .B(KEYINPUT101), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n815), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n892), .A2(new_n688), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n905), .B1(new_n352), .B2(new_n353), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n893), .A2(new_n906), .A3(new_n895), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT103), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n893), .A2(new_n906), .A3(new_n895), .A4(KEYINPUT103), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n354), .A2(new_n891), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n909), .A2(new_n910), .B1(new_n905), .B2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n904), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n901), .B1(new_n902), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n902), .B2(new_n914), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n899), .A2(new_n900), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n473), .A2(new_n710), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n648), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n917), .B(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n877), .A2(new_n878), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n867), .A2(new_n871), .A3(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n729), .A2(KEYINPUT31), .A3(new_n683), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT108), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n729), .A2(KEYINPUT108), .A3(KEYINPUT31), .A4(new_n683), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n925), .A2(new_n926), .B1(new_n713), .B2(new_n730), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT40), .ZN(new_n928));
  NOR4_X1   g0728(.A1(new_n912), .A2(new_n927), .A3(new_n928), .A4(new_n813), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n922), .A2(new_n929), .ZN(new_n930));
  NOR3_X1   g0730(.A1(new_n912), .A2(new_n927), .A3(new_n813), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n884), .B2(new_n885), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n928), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n472), .A2(new_n927), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n711), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n934), .B2(new_n935), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n920), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n273), .B2(new_n742), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n920), .A2(new_n937), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n850), .B1(new_n939), .B2(new_n940), .ZN(G367));
  NOR2_X1   g0741(.A1(new_n693), .A2(KEYINPUT110), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n650), .B(new_n627), .C1(new_n628), .C2(new_n688), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n649), .A2(new_n683), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n696), .A2(new_n945), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n946), .B(KEYINPUT45), .Z(new_n947));
  NOR2_X1   g0747(.A1(new_n696), .A2(new_n945), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT44), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n942), .B(new_n950), .Z(new_n951));
  NAND2_X1  g0751(.A1(new_n695), .A2(new_n569), .ZN(new_n952));
  OAI221_X1 g0752(.A(new_n952), .B1(new_n691), .B2(new_n695), .C1(new_n687), .C2(KEYINPUT111), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n687), .A2(KEYINPUT111), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n953), .B(new_n954), .Z(new_n955));
  NAND3_X1  g0755(.A1(new_n951), .A2(new_n738), .A3(new_n955), .ZN(new_n956));
  AND2_X1   g0756(.A1(new_n956), .A2(new_n738), .ZN(new_n957));
  XOR2_X1   g0757(.A(KEYINPUT109), .B(KEYINPUT41), .Z(new_n958));
  XNOR2_X1  g0758(.A(new_n698), .B(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n743), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n945), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n961), .A2(new_n952), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n963), .A2(KEYINPUT42), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n650), .B1(new_n943), .B2(new_n690), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n963), .A2(KEYINPUT42), .B1(new_n688), .B2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n688), .A2(new_n602), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n661), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n672), .A2(new_n967), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n964), .A2(new_n966), .B1(KEYINPUT43), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n970), .A2(KEYINPUT43), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n971), .B(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n692), .A2(new_n945), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n973), .B(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n960), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n216), .A2(new_n360), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n801), .B(new_n977), .C1(new_n790), .C2(new_n244), .ZN(new_n978));
  AND2_X1   g0778(.A1(new_n978), .A2(new_n787), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n749), .A2(G68), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n980), .B1(new_n201), .B2(new_n763), .C1(new_n767), .C2(new_n753), .ZN(new_n981));
  AOI22_X1  g0781(.A1(G50), .A2(new_n822), .B1(new_n777), .B2(G137), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n982), .B(new_n288), .C1(new_n265), .C2(new_n770), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n759), .A2(G143), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n984), .B1(new_n206), .B2(new_n761), .ZN(new_n985));
  OR3_X1    g0785(.A1(new_n981), .A2(new_n983), .A3(new_n985), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n551), .A2(new_n767), .B1(new_n760), .B2(new_n775), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(G97), .B2(new_n781), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n770), .A2(new_n502), .B1(new_n769), .B2(new_n827), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(G317), .B2(new_n777), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n411), .B1(new_n749), .B2(G107), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n988), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n763), .A2(new_n476), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT46), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n986), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT47), .Z(new_n996));
  OAI221_X1 g0796(.A(new_n979), .B1(new_n746), .B2(new_n996), .C1(new_n970), .C2(new_n803), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n976), .A2(new_n997), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(KEYINPUT112), .Z(G387));
  AOI21_X1  g0799(.A(new_n741), .B1(new_n955), .B2(new_n738), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n738), .B2(new_n955), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n830), .A2(G317), .B1(new_n822), .B2(G303), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n1002), .B1(new_n767), .B2(new_n775), .C1(new_n773), .C2(new_n760), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT113), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT48), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n749), .A2(G283), .B1(new_n764), .B2(G294), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1010), .A2(KEYINPUT49), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n411), .B1(G326), .B2(new_n777), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n476), .B2(new_n761), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT114), .Z(new_n1014));
  INV_X1    g0814(.A(KEYINPUT49), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1014), .B1(new_n1009), .B2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n763), .A2(new_n206), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(G159), .B2(new_n759), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n261), .B2(new_n767), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n596), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(new_n749), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n769), .A2(new_n202), .B1(new_n752), .B2(new_n265), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(G50), .B2(new_n830), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n431), .B1(G97), .B2(new_n781), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1021), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n1011), .A2(new_n1016), .B1(new_n1019), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT115), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n746), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n1027), .B2(new_n1026), .ZN(new_n1029));
  OR2_X1    g0829(.A1(new_n691), .A2(new_n803), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n241), .A2(new_n280), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n1031), .A2(new_n789), .B1(new_n699), .B2(new_n795), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n260), .A2(new_n272), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT50), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n280), .B1(new_n202), .B2(new_n206), .ZN(new_n1035));
  NOR3_X1   g0835(.A1(new_n1034), .A2(new_n699), .A3(new_n1035), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n1032), .A2(new_n1036), .B1(G107), .B2(new_n215), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n788), .B1(new_n1037), .B2(new_n801), .ZN(new_n1038));
  AND3_X1   g0838(.A1(new_n1029), .A2(new_n1030), .A3(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(new_n955), .B2(new_n786), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1001), .A2(new_n1040), .ZN(G393));
  OAI221_X1 g0841(.A(new_n801), .B1(new_n233), .B2(new_n215), .C1(new_n248), .C2(new_n790), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n787), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(G317), .A2(new_n759), .B1(new_n830), .B2(G311), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT52), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n370), .B1(new_n752), .B2(new_n773), .C1(new_n551), .C2(new_n769), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n229), .A2(new_n761), .B1(new_n763), .B2(new_n827), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n767), .A2(new_n502), .B1(new_n476), .B2(new_n748), .ZN(new_n1048));
  OR4_X1    g0848(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(G150), .A2(new_n759), .B1(new_n830), .B2(G159), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT116), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(KEYINPUT51), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n260), .A2(new_n822), .B1(new_n777), .B2(G143), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n748), .A2(new_n206), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n202), .A2(new_n763), .B1(new_n761), .B2(new_n434), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n1054), .B(new_n1055), .C1(G50), .C2(new_n766), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n1052), .A2(new_n411), .A3(new_n1053), .A4(new_n1056), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1051), .A2(KEYINPUT51), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1049), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1043), .B1(new_n1059), .B2(new_n745), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n945), .B2(new_n803), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n950), .B(new_n692), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n955), .A2(new_n738), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n1062), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n956), .A2(new_n698), .A3(new_n1064), .ZN(new_n1065));
  AND2_X1   g0865(.A1(new_n1065), .A2(KEYINPUT117), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1065), .A2(KEYINPUT117), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1061), .B1(new_n743), .B2(new_n1062), .C1(new_n1066), .C2(new_n1067), .ZN(G390));
  NAND2_X1  g0868(.A1(new_n914), .A2(new_n897), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n881), .A2(new_n883), .A3(new_n886), .A4(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n706), .A2(new_n688), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1071), .A2(new_n810), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1072), .A2(new_n811), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n922), .B(new_n897), .C1(new_n1073), .C2(new_n912), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1070), .A2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n912), .A2(new_n813), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n927), .A2(new_n711), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1075), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n737), .A2(new_n812), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1070), .B(new_n1074), .C1(new_n912), .C2(new_n1081), .ZN(new_n1082));
  AND2_X1   g0882(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n473), .A2(new_n1077), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n648), .A2(new_n918), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1081), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n811), .B(new_n1072), .C1(new_n1086), .C2(new_n913), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1077), .A2(new_n812), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n912), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1078), .B1(new_n1086), .B2(new_n913), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n1087), .A2(new_n1089), .B1(new_n1090), .B2(new_n904), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1085), .A2(new_n1091), .ZN(new_n1092));
  OR2_X1    g0892(.A1(new_n1083), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1080), .A2(new_n1082), .A3(new_n1092), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1093), .A2(new_n698), .A3(new_n1094), .ZN(new_n1095));
  OR2_X1    g0895(.A1(new_n887), .A2(new_n799), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n820), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n787), .B1(new_n260), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(G132), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n770), .A2(new_n1099), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(KEYINPUT54), .B(G143), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n288), .B1(new_n769), .B2(new_n1101), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n1100), .B(new_n1102), .C1(G125), .C2(new_n777), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n763), .A2(new_n265), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT53), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(G159), .A2(new_n749), .B1(new_n766), .B2(G137), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n759), .A2(G128), .B1(new_n781), .B2(G50), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1103), .A2(new_n1105), .A3(new_n1106), .A4(new_n1107), .ZN(new_n1108));
  OR2_X1    g0908(.A1(new_n1108), .A2(KEYINPUT118), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(KEYINPUT118), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1054), .B1(G283), .B2(new_n759), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n229), .B2(new_n767), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n770), .A2(new_n476), .B1(new_n752), .B2(new_n551), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n288), .B(new_n1113), .C1(G97), .C2(new_n822), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1114), .A2(new_n765), .A3(new_n836), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1109), .B(new_n1110), .C1(new_n1112), .C2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1098), .B1(new_n1116), .B2(new_n745), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n1083), .A2(new_n786), .B1(new_n1096), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1095), .A2(new_n1118), .ZN(G378));
  INV_X1    g0919(.A(new_n1085), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1094), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n930), .A2(new_n933), .A3(G330), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(KEYINPUT121), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT121), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n930), .A2(new_n933), .A3(new_n1124), .A4(G330), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n306), .A2(new_n856), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n311), .B(new_n1126), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1127), .B(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1123), .A2(new_n1125), .A3(new_n1130), .ZN(new_n1131));
  AND2_X1   g0931(.A1(new_n916), .A2(new_n900), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n934), .A2(new_n1124), .A3(G330), .A4(new_n1129), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1131), .A2(new_n899), .A3(new_n1132), .A4(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n917), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1121), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT57), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT122), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1121), .A2(new_n1136), .A3(KEYINPUT57), .A4(new_n1134), .ZN(new_n1142));
  AND2_X1   g0942(.A1(new_n1142), .A2(new_n698), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1137), .A2(KEYINPUT122), .A3(new_n1138), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1141), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n787), .B1(G50), .B2(new_n1097), .ZN(new_n1146));
  AOI211_X1 g0946(.A(G33), .B(G41), .C1(new_n777), .C2(G124), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1147), .B1(new_n761), .B2(new_n753), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n766), .A2(G132), .B1(new_n822), .B2(G137), .ZN(new_n1149));
  XOR2_X1   g0949(.A(new_n1149), .B(KEYINPUT120), .Z(new_n1150));
  AOI22_X1  g0950(.A1(G125), .A2(new_n759), .B1(new_n830), .B2(G128), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n1151), .B1(new_n265), .B2(new_n748), .C1(new_n763), .C2(new_n1101), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1148), .B1(new_n1154), .B2(KEYINPUT59), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1155), .B1(KEYINPUT59), .B2(new_n1154), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n411), .A2(G41), .ZN(new_n1157));
  AOI211_X1 g0957(.A(G50), .B(new_n1157), .C1(new_n262), .C2(new_n278), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1020), .A2(new_n822), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n830), .A2(G107), .B1(new_n777), .B2(G283), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1159), .A2(new_n980), .A3(new_n1157), .A4(new_n1160), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n761), .A2(new_n201), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n233), .A2(new_n767), .B1(new_n760), .B2(new_n476), .ZN(new_n1163));
  NOR4_X1   g0963(.A1(new_n1161), .A2(new_n1017), .A3(new_n1162), .A4(new_n1163), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1158), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1156), .B(new_n1166), .C1(new_n1165), .C2(new_n1164), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1146), .B1(new_n1167), .B2(new_n745), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1168), .B1(new_n1130), .B2(new_n799), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  AND2_X1   g0970(.A1(new_n1136), .A2(new_n1134), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1170), .B1(new_n1171), .B2(new_n786), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1145), .A2(new_n1172), .ZN(G375));
  INV_X1    g0973(.A(new_n1091), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n912), .A2(new_n798), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n787), .B1(G68), .B2(new_n1097), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n766), .A2(G116), .B1(new_n822), .B2(G107), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT123), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n760), .A2(new_n551), .B1(new_n761), .B2(new_n206), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(G97), .B2(new_n764), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n370), .B1(new_n770), .B2(new_n827), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(G303), .B2(new_n777), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1178), .A2(new_n1180), .A3(new_n1021), .A4(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(G159), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n201), .A2(new_n761), .B1(new_n763), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n777), .A2(G128), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1186), .B(new_n411), .C1(new_n265), .C2(new_n769), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1185), .B(new_n1187), .C1(G50), .C2(new_n749), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT124), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n759), .A2(G132), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n1190), .B1(new_n833), .B2(new_n770), .C1(new_n767), .C2(new_n1101), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1183), .B1(new_n1189), .B2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1176), .B1(new_n1192), .B2(new_n745), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n1174), .A2(new_n786), .B1(new_n1175), .B2(new_n1193), .ZN(new_n1194));
  OR2_X1    g0994(.A1(new_n1092), .A2(new_n959), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1120), .A2(new_n1174), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1194), .B1(new_n1195), .B2(new_n1196), .ZN(G381));
  NAND3_X1  g0997(.A1(new_n1001), .A2(new_n806), .A3(new_n1040), .ZN(new_n1198));
  OR4_X1    g0998(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1198), .ZN(new_n1199));
  OR4_X1    g0999(.A1(G387), .A2(new_n1199), .A3(G375), .A4(G378), .ZN(G407));
  INV_X1    g1000(.A(new_n1172), .ZN(new_n1201));
  AOI21_X1  g1001(.A(KEYINPUT122), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1142), .A2(new_n698), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1201), .B1(new_n1204), .B2(new_n1144), .ZN(new_n1205));
  INV_X1    g1005(.A(G378), .ZN(new_n1206));
  INV_X1    g1006(.A(G213), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1207), .A2(G343), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1205), .A2(new_n1206), .A3(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(G407), .A2(G213), .A3(new_n1209), .ZN(G409));
  NAND3_X1  g1010(.A1(new_n1145), .A2(G378), .A3(new_n1172), .ZN(new_n1211));
  OR2_X1    g1011(.A1(new_n1137), .A2(new_n959), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(new_n1172), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1206), .A2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1208), .B1(new_n1211), .B2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT60), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n1085), .A2(new_n1091), .A3(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1216), .B1(new_n1085), .B2(new_n1091), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n698), .B1(new_n1085), .B2(new_n1091), .C1(new_n1217), .C2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(new_n1194), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(new_n841), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1219), .A2(G384), .A3(new_n1194), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1208), .ZN(new_n1223));
  INV_X1    g1023(.A(G2897), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  AND3_X1   g1025(.A1(new_n1221), .A2(new_n1222), .A3(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1225), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1227));
  NOR3_X1   g1027(.A1(new_n1226), .A2(new_n1227), .A3(KEYINPUT125), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT125), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1222), .ZN(new_n1230));
  AOI21_X1  g1030(.A(G384), .B1(new_n1219), .B2(new_n1194), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n1230), .A2(new_n1231), .B1(new_n1224), .B2(new_n1223), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1221), .A2(new_n1222), .A3(new_n1225), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1229), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1228), .A2(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(KEYINPUT126), .B1(new_n1215), .B2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT126), .ZN(new_n1237));
  OAI21_X1  g1037(.A(KEYINPUT125), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1232), .A2(new_n1233), .A3(new_n1229), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(G378), .B1(new_n1172), .B2(new_n1212), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n1205), .B2(G378), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1237), .B(new_n1240), .C1(new_n1242), .C2(new_n1208), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1236), .A2(new_n1243), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1215), .A2(KEYINPUT63), .A3(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(G393), .A2(G396), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n1198), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT127), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1247), .A2(KEYINPUT127), .A3(new_n1198), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(G390), .ZN(new_n1253));
  AOI21_X1  g1053(.A(KEYINPUT112), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1253), .B1(G390), .B2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n998), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT61), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1253), .B(new_n998), .C1(G390), .C2(new_n1254), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1257), .A2(new_n1258), .A3(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1211), .A2(new_n1214), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1261), .A2(new_n1223), .A3(new_n1245), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT63), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1260), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1244), .A2(new_n1246), .A3(new_n1264), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1262), .A2(KEYINPUT62), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1258), .B1(new_n1215), .B2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT62), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1269), .B1(new_n1215), .B2(new_n1245), .ZN(new_n1270));
  NOR3_X1   g1070(.A1(new_n1266), .A2(new_n1268), .A3(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1257), .A2(new_n1259), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1265), .B1(new_n1271), .B2(new_n1273), .ZN(G405));
  NAND2_X1  g1074(.A1(G375), .A2(new_n1206), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(new_n1211), .ZN(new_n1276));
  OR2_X1    g1076(.A1(new_n1276), .A2(new_n1245), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1245), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n1272), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1277), .A2(new_n1273), .A3(new_n1278), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(G402));
endmodule


