//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 1 1 1 0 1 1 0 0 1 0 0 0 0 1 0 1 1 1 0 1 1 0 1 1 0 0 1 1 0 0 1 1 0 0 0 1 1 0 1 0 1 0 0 1 0 1 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:29 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1242, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1307, new_n1308, new_n1309;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0005(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G107), .A2(G264), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G87), .A2(G250), .ZN(new_n208));
  NAND3_X1  g0008(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(G97), .ZN(new_n210));
  INV_X1    g0010(.A(G257), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(G77), .ZN(new_n213));
  INV_X1    g0013(.A(G244), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G58), .ZN(new_n216));
  INV_X1    g0016(.A(G232), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NOR4_X1   g0018(.A1(new_n209), .A2(new_n212), .A3(new_n215), .A4(new_n218), .ZN(new_n219));
  XOR2_X1   g0019(.A(KEYINPUT64), .B(G68), .Z(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(G238), .ZN(new_n221));
  AOI22_X1  g0021(.A1(new_n219), .A2(new_n221), .B1(G1), .B2(G20), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT1), .Z(new_n223));
  INV_X1    g0023(.A(G1), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR3_X1   g0025(.A1(new_n224), .A2(new_n225), .A3(G13), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT0), .Z(new_n228));
  OAI21_X1  g0028(.A(G50), .B1(G58), .B2(G68), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NOR3_X1   g0030(.A1(new_n229), .A2(new_n225), .A3(new_n230), .ZN(new_n231));
  NOR3_X1   g0031(.A1(new_n223), .A2(new_n228), .A3(new_n231), .ZN(G361));
  XOR2_X1   g0032(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n233));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G226), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  INV_X1    g0038(.A(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT66), .B(G264), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n237), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT3), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(KEYINPUT7), .A3(new_n225), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT76), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT7), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT3), .B(G33), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n259), .B1(new_n260), .B2(G20), .ZN(new_n261));
  NAND4_X1  g0061(.A1(new_n255), .A2(KEYINPUT76), .A3(KEYINPUT7), .A4(new_n225), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n258), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G68), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G20), .A2(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G159), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n201), .B1(new_n220), .B2(G58), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n266), .B1(new_n267), .B2(new_n225), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n264), .A2(KEYINPUT16), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(new_n230), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT16), .ZN(new_n273));
  INV_X1    g0073(.A(new_n220), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n253), .A2(KEYINPUT77), .A3(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n252), .ZN(new_n276));
  AOI21_X1  g0076(.A(KEYINPUT77), .B1(new_n253), .B2(G33), .ZN(new_n277));
  OAI211_X1 g0077(.A(KEYINPUT7), .B(new_n225), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n274), .B1(new_n278), .B2(new_n261), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n273), .B1(new_n268), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n270), .A2(new_n272), .A3(new_n280), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n225), .A2(G1), .ZN(new_n282));
  XNOR2_X1  g0082(.A(new_n282), .B(KEYINPUT70), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT8), .B(G58), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  AND2_X1   g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n224), .A2(G13), .A3(G20), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n288), .A2(new_n272), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n286), .A2(new_n289), .B1(new_n288), .B2(new_n284), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n281), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G169), .ZN(new_n292));
  AND2_X1   g0092(.A1(G1), .A2(G13), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT69), .ZN(new_n294));
  INV_X1    g0094(.A(G41), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n293), .B(new_n294), .C1(new_n251), .C2(new_n295), .ZN(new_n296));
  AND2_X1   g0096(.A1(G33), .A2(G41), .ZN(new_n297));
  OAI21_X1  g0097(.A(KEYINPUT69), .B1(new_n297), .B2(new_n230), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(G33), .A2(G87), .ZN(new_n301));
  INV_X1    g0101(.A(G1698), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n302), .A2(G226), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n260), .B(new_n303), .C1(G223), .C2(G1698), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n300), .B1(new_n301), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n293), .B1(new_n251), .B2(new_n295), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n224), .B1(G41), .B2(G45), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n306), .A2(G232), .A3(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G45), .ZN(new_n309));
  AOI21_X1  g0109(.A(G1), .B1(new_n295), .B2(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(KEYINPUT67), .B1(new_n310), .B2(G274), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n224), .B(G274), .C1(G41), .C2(G45), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT67), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n308), .B1(new_n311), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n292), .B1(new_n305), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT78), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n304), .A2(new_n301), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n299), .ZN(new_n320));
  INV_X1    g0120(.A(G179), .ZN(new_n321));
  XNOR2_X1  g0121(.A(new_n312), .B(new_n313), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n322), .A2(KEYINPUT78), .A3(new_n308), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n318), .A2(new_n320), .A3(new_n321), .A4(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n316), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(KEYINPUT18), .B1(new_n291), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT18), .ZN(new_n328));
  AOI211_X1 g0128(.A(new_n328), .B(new_n325), .C1(new_n281), .C2(new_n290), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n290), .ZN(new_n331));
  INV_X1    g0131(.A(new_n272), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n268), .B1(G68), .B2(new_n263), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n332), .B1(new_n333), .B2(KEYINPUT16), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n331), .B1(new_n334), .B2(new_n280), .ZN(new_n335));
  INV_X1    g0135(.A(G200), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n336), .B1(new_n305), .B2(new_n315), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n318), .A2(new_n320), .A3(new_n323), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n337), .B1(new_n338), .B2(G190), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n335), .A2(KEYINPUT17), .A3(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n281), .A2(new_n290), .A3(new_n339), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT17), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT68), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n345), .B1(new_n255), .B2(new_n302), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n260), .A2(KEYINPUT68), .A3(G1698), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n346), .A2(G238), .A3(new_n347), .ZN(new_n348));
  AND3_X1   g0148(.A1(new_n252), .A2(new_n254), .A3(new_n302), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n349), .A2(G232), .B1(G107), .B2(new_n255), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n299), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n297), .A2(new_n230), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n353), .A2(new_n310), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(G244), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n352), .A2(new_n322), .A3(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n356), .A2(G179), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT74), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n287), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n224), .A2(KEYINPUT74), .A3(G13), .A4(G20), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n362), .A2(new_n272), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n363), .A2(G77), .A3(new_n283), .ZN(new_n364));
  INV_X1    g0164(.A(new_n362), .ZN(new_n365));
  AND2_X1   g0165(.A1(KEYINPUT15), .A2(G87), .ZN(new_n366));
  NOR2_X1   g0166(.A1(KEYINPUT15), .A2(G87), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n225), .A2(G33), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  OR2_X1    g0171(.A1(new_n371), .A2(KEYINPUT73), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(KEYINPUT73), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n265), .ZN(new_n375));
  OAI22_X1  g0175(.A1(new_n284), .A2(new_n375), .B1(new_n225), .B2(new_n213), .ZN(new_n376));
  AND2_X1   g0176(.A1(new_n376), .A2(KEYINPUT72), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n376), .A2(KEYINPUT72), .ZN(new_n378));
  NOR3_X1   g0178(.A1(new_n374), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  OAI221_X1 g0179(.A(new_n364), .B1(G77), .B2(new_n365), .C1(new_n379), .C2(new_n332), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n356), .A2(new_n292), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n358), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  OR3_X1    g0183(.A1(new_n330), .A2(new_n344), .A3(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n346), .A2(G223), .A3(new_n347), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n349), .A2(G222), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n385), .B(new_n386), .C1(new_n213), .C2(new_n260), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n299), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n354), .A2(G226), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(new_n322), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(G200), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n203), .A2(G20), .ZN(new_n392));
  INV_X1    g0192(.A(G150), .ZN(new_n393));
  OAI221_X1 g0193(.A(new_n392), .B1(new_n393), .B2(new_n375), .C1(new_n369), .C2(new_n284), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n272), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n288), .A2(new_n202), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n283), .A2(G50), .A3(new_n289), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  XNOR2_X1  g0198(.A(new_n398), .B(KEYINPUT9), .ZN(new_n399));
  INV_X1    g0199(.A(G190), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n391), .B(new_n399), .C1(new_n400), .C2(new_n390), .ZN(new_n401));
  XNOR2_X1  g0201(.A(new_n401), .B(KEYINPUT10), .ZN(new_n402));
  OR2_X1    g0202(.A1(new_n390), .A2(G179), .ZN(new_n403));
  OR2_X1    g0203(.A1(new_n403), .A2(KEYINPUT71), .ZN(new_n404));
  INV_X1    g0204(.A(new_n398), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n405), .B1(new_n390), .B2(new_n292), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n403), .A2(KEYINPUT71), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n404), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n402), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT14), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n354), .A2(G238), .ZN(new_n411));
  NOR2_X1   g0211(.A1(G226), .A2(G1698), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n412), .B1(new_n217), .B2(G1698), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n413), .A2(new_n260), .B1(G33), .B2(G97), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n411), .B(new_n322), .C1(new_n300), .C2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT13), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n413), .A2(new_n260), .ZN(new_n417));
  NAND2_X1  g0217(.A1(G33), .A2(G97), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n299), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT13), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n420), .A2(new_n421), .A3(new_n411), .A4(new_n322), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n416), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n410), .B1(new_n423), .B2(G169), .ZN(new_n424));
  AOI211_X1 g0224(.A(KEYINPUT14), .B(new_n292), .C1(new_n416), .C2(new_n422), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n423), .A2(new_n321), .ZN(new_n426));
  NOR3_X1   g0226(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n220), .A2(new_n225), .ZN(new_n428));
  OAI22_X1  g0228(.A1(new_n375), .A2(new_n202), .B1(new_n369), .B2(new_n213), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n272), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  XNOR2_X1  g0230(.A(new_n430), .B(KEYINPUT11), .ZN(new_n431));
  OR2_X1    g0231(.A1(new_n288), .A2(KEYINPUT12), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n363), .A2(new_n283), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(KEYINPUT12), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(G68), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n274), .A2(new_n362), .A3(KEYINPUT12), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n431), .A2(new_n432), .A3(new_n435), .A4(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n427), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n416), .A2(new_n422), .A3(KEYINPUT75), .A4(G190), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n423), .A2(G200), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT75), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(new_n423), .B2(new_n400), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n438), .A2(new_n441), .A3(new_n442), .A4(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n440), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n356), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(G190), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n365), .A2(G77), .ZN(new_n449));
  INV_X1    g0249(.A(new_n379), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n449), .B1(new_n450), .B2(new_n272), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n356), .A2(G200), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n448), .A2(new_n451), .A3(new_n364), .A4(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g0254(.A1(new_n384), .A2(new_n409), .A3(new_n446), .A4(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(G116), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n456), .B1(new_n224), .B2(G33), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n363), .A2(new_n457), .ZN(new_n458));
  OR2_X1    g0258(.A1(KEYINPUT81), .A2(G116), .ZN(new_n459));
  NAND2_X1  g0259(.A1(KEYINPUT81), .A2(G116), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n362), .A2(KEYINPUT87), .A3(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(KEYINPUT87), .B1(new_n362), .B2(new_n461), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n458), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n461), .A2(G20), .ZN(new_n466));
  AOI21_X1  g0266(.A(G20), .B1(G33), .B2(G283), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n251), .A2(G97), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n469), .A2(KEYINPUT88), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT88), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n471), .B1(new_n467), .B2(new_n468), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n272), .B(new_n466), .C1(new_n470), .C2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT20), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g0275(.A(new_n469), .B(KEYINPUT88), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n476), .A2(KEYINPUT20), .A3(new_n272), .A4(new_n466), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n465), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n260), .A2(G257), .A3(new_n302), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n260), .A2(G264), .A3(G1698), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n255), .A2(G303), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n299), .ZN(new_n483));
  XOR2_X1   g0283(.A(KEYINPUT5), .B(G41), .Z(new_n484));
  NOR2_X1   g0284(.A1(new_n309), .A2(G1), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n306), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(KEYINPUT86), .B1(new_n487), .B2(new_n239), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n485), .A2(G274), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  XNOR2_X1  g0291(.A(KEYINPUT5), .B(G41), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n353), .B1(new_n492), .B2(new_n485), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT86), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n493), .A2(new_n494), .A3(G270), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n483), .A2(new_n488), .A3(new_n491), .A4(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G169), .ZN(new_n497));
  OAI21_X1  g0297(.A(KEYINPUT89), .B1(new_n478), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT21), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n477), .A2(new_n475), .ZN(new_n500));
  INV_X1    g0300(.A(new_n464), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n501), .A2(new_n462), .B1(new_n363), .B2(new_n457), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT89), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n503), .A2(new_n504), .A3(G169), .A4(new_n496), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n498), .A2(new_n499), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n490), .B1(new_n482), .B2(new_n299), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n507), .A2(G179), .A3(new_n488), .A4(new_n495), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n508), .B1(new_n497), .B2(new_n499), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n503), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n496), .A2(G200), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n478), .B(new_n511), .C1(new_n400), .C2(new_n496), .ZN(new_n512));
  AND3_X1   g0312(.A1(new_n506), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n252), .A2(new_n254), .A3(G257), .A4(G1698), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n252), .A2(new_n254), .A3(G250), .A4(new_n302), .ZN(new_n515));
  NAND2_X1  g0315(.A1(G33), .A2(G294), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n299), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n493), .A2(G264), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n518), .A2(new_n519), .A3(new_n491), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G169), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT90), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AND2_X1   g0323(.A1(new_n518), .A2(new_n519), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n524), .A2(G179), .A3(new_n491), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n520), .A2(KEYINPUT90), .A3(G169), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n523), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n252), .A2(new_n254), .A3(new_n225), .A4(G87), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(KEYINPUT22), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT22), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n260), .A2(new_n530), .A3(new_n225), .A4(G87), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n461), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n370), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n225), .A2(G107), .ZN(new_n535));
  XNOR2_X1  g0335(.A(new_n535), .B(KEYINPUT23), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n532), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT24), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n532), .A2(KEYINPUT24), .A3(new_n534), .A4(new_n536), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n539), .A2(new_n272), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n224), .A2(G33), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n287), .A2(new_n542), .A3(new_n230), .A4(new_n271), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(G107), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n287), .A2(G107), .ZN(new_n546));
  XNOR2_X1  g0346(.A(new_n546), .B(KEYINPUT25), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n541), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n527), .A2(new_n548), .ZN(new_n549));
  OR2_X1    g0349(.A1(G238), .A2(G1698), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n214), .A2(G1698), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n252), .A2(new_n550), .A3(new_n254), .A4(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n459), .A2(G33), .A3(new_n460), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(KEYINPUT82), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT82), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n552), .A2(new_n556), .A3(new_n553), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n555), .A2(new_n299), .A3(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n353), .A2(new_n485), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(G250), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n560), .A2(new_n489), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n558), .A2(new_n321), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(G169), .B1(new_n558), .B2(new_n561), .ZN(new_n563));
  OAI21_X1  g0363(.A(KEYINPUT83), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n368), .B1(new_n360), .B2(new_n361), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT19), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n225), .B1(new_n418), .B2(new_n566), .ZN(new_n567));
  NOR2_X1   g0367(.A1(G97), .A2(G107), .ZN(new_n568));
  INV_X1    g0368(.A(G87), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n252), .A2(new_n254), .A3(new_n225), .A4(G68), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n225), .A2(G33), .A3(G97), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n566), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n571), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n565), .B1(new_n575), .B2(new_n272), .ZN(new_n576));
  INV_X1    g0376(.A(new_n368), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n577), .A2(new_n543), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT84), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n576), .A2(KEYINPUT84), .A3(new_n579), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n558), .A2(new_n561), .A3(new_n321), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT83), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n582), .A2(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n564), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n558), .A2(new_n561), .A3(G190), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT85), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n558), .A2(new_n561), .A3(KEYINPUT85), .A4(G190), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n544), .A2(G87), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n576), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n558), .A2(new_n561), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n594), .B1(new_n595), .B2(G200), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n520), .A2(new_n336), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n598), .B1(G190), .B2(new_n520), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n599), .A2(new_n545), .A3(new_n547), .A4(new_n541), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n549), .A2(new_n587), .A3(new_n597), .A4(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n287), .A2(G97), .ZN(new_n603));
  INV_X1    g0403(.A(G107), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n604), .B1(new_n278), .B2(new_n261), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n375), .A2(new_n213), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT6), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n210), .A2(new_n604), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n607), .B1(new_n608), .B2(new_n568), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n604), .A2(KEYINPUT6), .A3(G97), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n225), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  OR3_X1    g0411(.A1(new_n605), .A2(new_n606), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n603), .B1(new_n612), .B2(new_n272), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n252), .A2(new_n254), .A3(G244), .A4(new_n302), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT80), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT4), .ZN(new_n616));
  NOR3_X1   g0416(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n614), .A2(new_n616), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(KEYINPUT79), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT79), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n614), .A2(new_n620), .A3(new_n616), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n617), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n615), .B1(new_n614), .B2(new_n616), .ZN(new_n623));
  NAND2_X1  g0423(.A1(G33), .A2(G283), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n260), .A2(G250), .A3(G1698), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n300), .B1(new_n622), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n490), .B1(new_n493), .B2(G257), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(G200), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n544), .A2(G97), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n349), .A2(KEYINPUT80), .A3(KEYINPUT4), .A4(G244), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n614), .A2(new_n620), .A3(new_n616), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n620), .B1(new_n614), .B2(new_n616), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n299), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n637), .A2(G190), .A3(new_n628), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n613), .A2(new_n630), .A3(new_n631), .A4(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n292), .B1(new_n627), .B2(new_n629), .ZN(new_n640));
  INV_X1    g0440(.A(new_n603), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n605), .A2(new_n606), .A3(new_n611), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n641), .B(new_n631), .C1(new_n642), .C2(new_n332), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n637), .A2(new_n321), .A3(new_n628), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n640), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n639), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n455), .A2(new_n513), .A3(new_n602), .A4(new_n647), .ZN(new_n648));
  XOR2_X1   g0448(.A(new_n648), .B(KEYINPUT91), .Z(G372));
  INV_X1    g0449(.A(KEYINPUT92), .ZN(new_n650));
  INV_X1    g0450(.A(new_n594), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n560), .A2(new_n489), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n552), .A2(new_n556), .A3(new_n553), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n556), .B1(new_n552), .B2(new_n553), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n652), .B1(new_n655), .B2(new_n299), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n651), .B1(new_n656), .B2(new_n336), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n657), .B1(new_n590), .B2(new_n591), .ZN(new_n658));
  AOI21_X1  g0458(.A(KEYINPUT84), .B1(new_n576), .B2(new_n579), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n567), .A2(new_n570), .B1(new_n566), .B2(new_n573), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n332), .B1(new_n660), .B2(new_n572), .ZN(new_n661));
  NOR4_X1   g0461(.A1(new_n661), .A2(new_n578), .A3(new_n581), .A4(new_n565), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  NOR3_X1   g0463(.A1(new_n663), .A2(new_n562), .A3(new_n563), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n650), .B1(new_n658), .B2(new_n664), .ZN(new_n665));
  OAI221_X1 g0465(.A(new_n584), .B1(new_n659), .B2(new_n662), .C1(G169), .C2(new_n656), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n597), .A2(new_n666), .A3(KEYINPUT92), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT93), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n645), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n640), .A2(new_n643), .A3(KEYINPUT93), .A4(new_n644), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT26), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n668), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n639), .A2(new_n600), .A3(new_n645), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n506), .A2(new_n510), .A3(new_n549), .ZN(new_n676));
  AOI21_X1  g0476(.A(KEYINPUT92), .B1(new_n597), .B2(new_n666), .ZN(new_n677));
  AND3_X1   g0477(.A1(new_n597), .A2(new_n666), .A3(KEYINPUT92), .ZN(new_n678));
  OAI211_X1 g0478(.A(new_n675), .B(new_n676), .C1(new_n677), .C2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n645), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n680), .A2(new_n597), .A3(new_n587), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(KEYINPUT26), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n674), .A2(new_n679), .A3(new_n666), .A4(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n455), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n408), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n439), .B1(new_n445), .B2(new_n383), .ZN(new_n686));
  OAI22_X1  g0486(.A1(new_n686), .A2(new_n344), .B1(new_n327), .B2(new_n329), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n685), .B1(new_n687), .B2(new_n402), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n684), .A2(new_n688), .ZN(G369));
  INV_X1    g0489(.A(G13), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(G20), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(new_n224), .ZN(new_n692));
  OR2_X1    g0492(.A1(new_n692), .A2(KEYINPUT27), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(KEYINPUT27), .ZN(new_n694));
  AND3_X1   g0494(.A1(new_n693), .A2(G213), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(G343), .ZN(new_n696));
  XNOR2_X1  g0496(.A(new_n696), .B(KEYINPUT94), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n513), .B1(new_n478), .B2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT95), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n506), .A2(new_n510), .ZN(new_n700));
  INV_X1    g0500(.A(new_n697), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(new_n503), .A3(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n698), .A2(new_n699), .A3(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n699), .B1(new_n698), .B2(new_n702), .ZN(new_n705));
  OAI21_X1  g0505(.A(G330), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n701), .A2(new_n548), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n549), .A2(new_n600), .ZN(new_n709));
  OAI22_X1  g0509(.A1(new_n708), .A2(new_n709), .B1(new_n549), .B2(new_n697), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n549), .A2(new_n701), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n701), .B1(new_n506), .B2(new_n510), .ZN(new_n713));
  INV_X1    g0513(.A(new_n709), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n712), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n711), .A2(new_n715), .ZN(G399));
  NAND2_X1  g0516(.A1(new_n226), .A2(new_n295), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(G1), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n568), .A2(new_n569), .A3(new_n456), .ZN(new_n719));
  OAI22_X1  g0519(.A1(new_n718), .A2(new_n719), .B1(new_n229), .B2(new_n717), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT28), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT99), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n673), .B1(new_n668), .B2(new_n672), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n666), .B1(new_n681), .B2(KEYINPUT26), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n722), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n587), .A2(new_n597), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(new_n645), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n664), .B1(new_n727), .B2(new_n673), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n670), .A2(new_n671), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n729), .B1(new_n665), .B2(new_n667), .ZN(new_n730));
  OAI211_X1 g0530(.A(new_n728), .B(KEYINPUT99), .C1(new_n730), .C2(new_n673), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n725), .A2(new_n679), .A3(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n732), .A2(KEYINPUT29), .A3(new_n697), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT98), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n683), .A2(new_n697), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT29), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  AOI211_X1 g0537(.A(KEYINPUT98), .B(KEYINPUT29), .C1(new_n683), .C2(new_n697), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n733), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(KEYINPUT96), .A2(KEYINPUT30), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n637), .A2(new_n656), .A3(new_n524), .A4(new_n628), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n740), .B1(new_n741), .B2(new_n508), .ZN(new_n742));
  AOI21_X1  g0542(.A(G179), .B1(new_n637), .B2(new_n628), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n743), .A2(new_n496), .A3(new_n520), .A4(new_n595), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n627), .A2(new_n629), .ZN(new_n745));
  INV_X1    g0545(.A(new_n508), .ZN(new_n746));
  INV_X1    g0546(.A(new_n740), .ZN(new_n747));
  AND3_X1   g0547(.A1(new_n524), .A2(new_n561), .A3(new_n558), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n745), .A2(new_n746), .A3(new_n747), .A4(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n742), .A2(new_n744), .A3(new_n749), .ZN(new_n750));
  AND3_X1   g0550(.A1(new_n750), .A2(KEYINPUT31), .A3(new_n701), .ZN(new_n751));
  AOI21_X1  g0551(.A(KEYINPUT31), .B1(new_n750), .B2(new_n701), .ZN(new_n752));
  OAI21_X1  g0552(.A(KEYINPUT97), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n750), .A2(new_n701), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT31), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT97), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n750), .A2(KEYINPUT31), .A3(new_n701), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n756), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n513), .A2(new_n602), .A3(new_n647), .A4(new_n697), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n753), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G330), .ZN(new_n762));
  AND2_X1   g0562(.A1(new_n739), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n721), .B1(new_n763), .B2(G1), .ZN(G364));
  NOR2_X1   g0564(.A1(G13), .A2(G33), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G20), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n698), .A2(new_n702), .A3(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n225), .A2(G190), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n769), .A2(G179), .A3(new_n336), .ZN(new_n770));
  INV_X1    g0570(.A(G311), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n769), .A2(G179), .A3(G200), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  XNOR2_X1  g0574(.A(KEYINPUT33), .B(G317), .ZN(new_n775));
  NOR2_X1   g0575(.A1(G179), .A2(G200), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n225), .B1(new_n776), .B2(G190), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n774), .A2(new_n775), .B1(new_n778), .B2(G294), .ZN(new_n779));
  INV_X1    g0579(.A(G283), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n336), .A2(G179), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n769), .A2(new_n781), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n779), .B(new_n255), .C1(new_n780), .C2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n769), .A2(new_n776), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n772), .B(new_n783), .C1(G329), .C2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n225), .A2(new_n400), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n787), .A2(G179), .A3(new_n336), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G322), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n787), .A2(new_n781), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G303), .ZN(new_n793));
  NOR4_X1   g0593(.A1(new_n225), .A2(new_n321), .A3(new_n400), .A4(new_n336), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G326), .ZN(new_n795));
  NAND4_X1  g0595(.A1(new_n786), .A2(new_n790), .A3(new_n793), .A4(new_n795), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT102), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n777), .A2(new_n210), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n792), .A2(G87), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n799), .B(new_n260), .C1(new_n216), .C2(new_n788), .ZN(new_n800));
  INV_X1    g0600(.A(new_n782), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n798), .B(new_n800), .C1(G107), .C2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n794), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(new_n202), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n785), .A2(G159), .ZN(new_n805));
  INV_X1    g0605(.A(G68), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n805), .A2(KEYINPUT32), .B1(new_n806), .B2(new_n773), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n804), .B(new_n807), .C1(KEYINPUT32), .C2(new_n805), .ZN(new_n808));
  OR2_X1    g0608(.A1(new_n770), .A2(KEYINPUT101), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n770), .A2(KEYINPUT101), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n802), .B(new_n808), .C1(new_n213), .C2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n797), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n230), .B1(G20), .B2(new_n292), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n718), .B1(G45), .B2(new_n691), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n255), .A2(new_n226), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(KEYINPUT100), .ZN(new_n818));
  INV_X1    g0618(.A(new_n229), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(new_n309), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n818), .B(new_n820), .C1(new_n309), .C2(new_n249), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n260), .A2(new_n226), .A3(G355), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n821), .B(new_n822), .C1(G116), .C2(new_n226), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n767), .A2(new_n814), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n768), .A2(new_n815), .A3(new_n816), .A4(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n816), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n706), .A2(new_n827), .ZN(new_n828));
  NOR3_X1   g0628(.A1(new_n704), .A2(G330), .A3(new_n705), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n826), .B1(new_n828), .B2(new_n829), .ZN(G396));
  NOR2_X1   g0630(.A1(new_n382), .A2(new_n701), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n701), .A2(new_n380), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n453), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n831), .B1(new_n382), .B2(new_n833), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n735), .B(new_n834), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(new_n762), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n827), .ZN(new_n837));
  OR2_X1    g0637(.A1(new_n834), .A2(new_n766), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n255), .B1(new_n791), .B2(new_n604), .C1(new_n780), .C2(new_n773), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n798), .B(new_n839), .C1(G294), .C2(new_n789), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n801), .A2(G87), .ZN(new_n841));
  INV_X1    g0641(.A(new_n811), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n533), .ZN(new_n843));
  AOI22_X1  g0643(.A1(G303), .A2(new_n794), .B1(new_n785), .B2(G311), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n840), .A2(new_n841), .A3(new_n843), .A4(new_n844), .ZN(new_n845));
  AOI22_X1  g0645(.A1(G143), .A2(new_n789), .B1(new_n774), .B2(G150), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n794), .A2(G137), .ZN(new_n847));
  INV_X1    g0647(.A(G159), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n846), .B(new_n847), .C1(new_n811), .C2(new_n848), .ZN(new_n849));
  XNOR2_X1  g0649(.A(KEYINPUT103), .B(KEYINPUT34), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n849), .A2(new_n850), .B1(new_n216), .B2(new_n777), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n851), .B1(G50), .B2(new_n792), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n801), .A2(G68), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n849), .A2(new_n850), .B1(G132), .B2(new_n785), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n845), .B1(new_n855), .B2(new_n255), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n814), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n814), .A2(new_n765), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n213), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n838), .A2(new_n816), .A3(new_n857), .A4(new_n859), .ZN(new_n860));
  XOR2_X1   g0660(.A(new_n860), .B(KEYINPUT104), .Z(new_n861));
  NAND2_X1  g0661(.A1(new_n837), .A2(new_n861), .ZN(G384));
  AND2_X1   g0662(.A1(new_n609), .A2(new_n610), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT35), .ZN(new_n864));
  AOI211_X1 g0664(.A(new_n225), .B(new_n230), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n865), .B(G116), .C1(new_n864), .C2(new_n863), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n866), .B(KEYINPUT36), .ZN(new_n867));
  AOI211_X1 g0667(.A(new_n213), .B(new_n229), .C1(new_n220), .C2(G58), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n868), .B(KEYINPUT105), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n806), .A2(G50), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n870), .B(KEYINPUT106), .ZN(new_n871));
  OAI211_X1 g0671(.A(G1), .B(new_n690), .C1(new_n869), .C2(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n751), .A2(new_n752), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n760), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n701), .A2(new_n437), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n445), .B(new_n875), .C1(new_n427), .C2(new_n438), .ZN(new_n876));
  OR2_X1    g0676(.A1(new_n427), .A2(new_n875), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n878), .A2(new_n834), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n334), .B1(KEYINPUT16), .B2(new_n333), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n290), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n695), .B(new_n881), .C1(new_n330), .C2(new_n344), .ZN(new_n882));
  INV_X1    g0682(.A(new_n695), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n880), .A2(new_n290), .B1(new_n325), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n341), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT37), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n291), .A2(new_n326), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n291), .A2(new_n695), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT37), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n887), .A2(new_n888), .A3(new_n889), .A4(new_n341), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  AND3_X1   g0691(.A1(new_n882), .A2(KEYINPUT38), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT38), .B1(new_n882), .B2(new_n891), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n874), .B(new_n879), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT40), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n887), .A2(new_n888), .A3(new_n341), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(KEYINPUT37), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n890), .ZN(new_n899));
  INV_X1    g0699(.A(new_n888), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n900), .B1(new_n330), .B2(new_n344), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT38), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n892), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n879), .A2(new_n874), .A3(KEYINPUT40), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT107), .ZN(new_n905));
  NOR3_X1   g0705(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n879), .A2(new_n874), .A3(KEYINPUT40), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n899), .A2(new_n901), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT38), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n882), .A2(KEYINPUT38), .A3(new_n891), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT107), .B1(new_n907), .B2(new_n912), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n896), .B(G330), .C1(new_n906), .C2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n455), .A2(G330), .A3(new_n874), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n905), .B1(new_n903), .B2(new_n904), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n907), .A2(KEYINPUT107), .A3(new_n912), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n917), .A2(new_n918), .B1(new_n895), .B2(new_n894), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n919), .A2(new_n455), .A3(new_n874), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n916), .A2(new_n920), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n733), .B(new_n455), .C1(new_n737), .C2(new_n738), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n688), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n921), .B(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT39), .ZN(new_n925));
  NOR3_X1   g0725(.A1(new_n892), .A2(new_n893), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT39), .B1(new_n910), .B2(new_n911), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n440), .A2(new_n701), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n878), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n683), .A2(new_n697), .A3(new_n834), .ZN(new_n932));
  INV_X1    g0732(.A(new_n831), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OR2_X1    g0734(.A1(new_n892), .A2(new_n893), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n330), .A2(new_n883), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n930), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n924), .B(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n691), .A2(new_n224), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n867), .B(new_n872), .C1(new_n939), .C2(new_n940), .ZN(G367));
  OAI21_X1  g0741(.A(new_n668), .B1(new_n651), .B2(new_n697), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n664), .A2(new_n594), .A3(new_n701), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n767), .ZN(new_n946));
  INV_X1    g0746(.A(new_n818), .ZN(new_n947));
  OAI221_X1 g0747(.A(new_n824), .B1(new_n226), .B2(new_n577), .C1(new_n242), .C2(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n777), .A2(new_n604), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n792), .A2(KEYINPUT46), .A3(G116), .ZN(new_n950));
  INV_X1    g0750(.A(G317), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n950), .B(new_n255), .C1(new_n951), .C2(new_n784), .ZN(new_n952));
  AOI211_X1 g0752(.A(new_n949), .B(new_n952), .C1(G303), .C2(new_n789), .ZN(new_n953));
  AOI21_X1  g0753(.A(KEYINPUT46), .B1(new_n792), .B2(new_n533), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n801), .A2(G97), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n803), .B2(new_n771), .ZN(new_n956));
  AOI211_X1 g0756(.A(new_n954), .B(new_n956), .C1(G294), .C2(new_n774), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n953), .B(new_n957), .C1(new_n780), .C2(new_n811), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n260), .B1(new_n811), .B2(new_n202), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n777), .A2(new_n806), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n788), .A2(new_n393), .B1(new_n782), .B2(new_n213), .ZN(new_n961));
  NOR3_X1   g0761(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n794), .A2(G143), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n848), .A2(new_n773), .B1(new_n791), .B2(new_n216), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(G137), .B2(new_n785), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n962), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n958), .A2(new_n966), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT47), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n814), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n946), .A2(new_n816), .A3(new_n948), .A4(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n224), .B1(new_n691), .B2(G45), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT45), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT112), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n697), .B1(new_n613), .B2(new_n631), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n646), .A2(new_n975), .B1(new_n645), .B2(new_n697), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT109), .ZN(new_n977));
  AND2_X1   g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n976), .A2(new_n977), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n715), .B(new_n974), .C1(new_n978), .C2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n976), .B(new_n977), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n974), .B1(new_n982), .B2(new_n715), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n973), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n978), .A2(new_n979), .ZN(new_n985));
  INV_X1    g0785(.A(new_n715), .ZN(new_n986));
  OAI21_X1  g0786(.A(KEYINPUT112), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n987), .A2(KEYINPUT45), .A3(new_n980), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT44), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n982), .B2(new_n715), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n985), .A2(KEYINPUT44), .A3(new_n986), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n984), .A2(new_n988), .A3(new_n992), .ZN(new_n993));
  AND2_X1   g0793(.A1(new_n707), .A2(new_n710), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n711), .A2(new_n992), .A3(new_n984), .A4(new_n988), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n710), .A2(new_n713), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT113), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n997), .B(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n713), .A2(new_n714), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT114), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1000), .B(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT115), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1003), .B1(new_n707), .B2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n706), .A2(KEYINPUT115), .A3(new_n999), .A4(new_n1002), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n763), .A2(new_n995), .A3(new_n996), .A4(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n763), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n717), .B(KEYINPUT41), .Z(new_n1010));
  AOI21_X1  g0810(.A(new_n972), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n985), .A2(new_n1000), .ZN(new_n1012));
  XOR2_X1   g0812(.A(KEYINPUT110), .B(KEYINPUT42), .Z(new_n1013));
  XOR2_X1   g0813(.A(new_n1012), .B(new_n1013), .Z(new_n1014));
  OAI21_X1  g0814(.A(new_n645), .B1(new_n985), .B2(new_n549), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(new_n697), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n1014), .A2(new_n1016), .B1(KEYINPUT43), .B2(new_n944), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT111), .ZN(new_n1019));
  OR3_X1    g0819(.A1(new_n944), .A2(KEYINPUT108), .A3(KEYINPUT43), .ZN(new_n1020));
  OAI21_X1  g0820(.A(KEYINPUT108), .B1(new_n944), .B2(KEYINPUT43), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1019), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1020), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n994), .A2(new_n982), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1024), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n711), .A2(new_n985), .B1(new_n1026), .B2(new_n1022), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1018), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1017), .A2(new_n1027), .A3(new_n1025), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n970), .B1(new_n1011), .B2(new_n1031), .ZN(G387));
  OAI21_X1  g0832(.A(new_n818), .B1(new_n237), .B2(new_n309), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n260), .A2(new_n226), .A3(new_n719), .ZN(new_n1034));
  AOI211_X1 g0834(.A(G45), .B(new_n719), .C1(G68), .C2(G77), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n284), .A2(G50), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT50), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n1033), .A2(new_n1034), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n226), .A2(G107), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n824), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n767), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1040), .B1(new_n710), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n794), .A2(G322), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1043), .B1(new_n771), .B2(new_n773), .C1(new_n951), .C2(new_n788), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(G303), .B2(new_n842), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n1045), .B(KEYINPUT48), .Z(new_n1046));
  INV_X1    g0846(.A(G294), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1046), .B1(new_n780), .B2(new_n777), .C1(new_n1047), .C2(new_n791), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT49), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n260), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n785), .A2(G326), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n801), .A2(new_n533), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n260), .B1(new_n202), .B2(new_n788), .C1(new_n803), .C2(new_n848), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n577), .A2(new_n777), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n284), .A2(new_n773), .B1(new_n770), .B2(new_n806), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n1056), .B(new_n1057), .C1(G77), .C2(new_n792), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1058), .B(new_n955), .C1(new_n393), .C2(new_n784), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1054), .B1(new_n1055), .B2(new_n1059), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n827), .B(new_n1042), .C1(new_n1060), .C2(new_n814), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(new_n1007), .B2(new_n972), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n763), .A2(new_n1007), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n717), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n763), .B2(new_n1007), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1062), .B1(new_n1064), .B2(new_n1066), .ZN(G393));
  NAND3_X1  g0867(.A1(new_n995), .A2(new_n972), .A3(new_n996), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n985), .A2(new_n767), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n803), .A2(new_n951), .B1(new_n771), .B2(new_n788), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT52), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n785), .A2(G322), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n774), .A2(G303), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n1047), .A2(new_n770), .B1(new_n791), .B2(new_n780), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(new_n533), .B2(new_n778), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .A4(new_n1075), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n260), .B(new_n1076), .C1(G107), .C2(new_n801), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n255), .B1(new_n785), .B2(G143), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n792), .A2(new_n220), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n778), .A2(G77), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1078), .A2(new_n1079), .A3(new_n841), .A4(new_n1080), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n803), .A2(new_n393), .B1(new_n848), .B2(new_n788), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT51), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n284), .B2(new_n811), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n1081), .B(new_n1084), .C1(G50), .C2(new_n774), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n814), .B1(new_n1077), .B2(new_n1085), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n824), .B1(new_n210), .B2(new_n226), .C1(new_n947), .C2(new_n246), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1069), .A2(new_n816), .A3(new_n1086), .A4(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1068), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(KEYINPUT116), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT116), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1068), .A2(new_n1091), .A3(new_n1088), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n995), .A2(new_n996), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n717), .B1(new_n1063), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n1008), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1093), .A2(new_n1096), .ZN(G390));
  AND3_X1   g0897(.A1(new_n922), .A2(new_n688), .A3(new_n915), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n756), .A2(new_n758), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n506), .A2(new_n510), .A3(new_n512), .ZN(new_n1100));
  NOR4_X1   g0900(.A1(new_n1100), .A2(new_n601), .A3(new_n646), .A4(new_n701), .ZN(new_n1101));
  OAI211_X1 g0901(.A(KEYINPUT117), .B(G330), .C1(new_n1099), .C2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n834), .ZN(new_n1103));
  AOI21_X1  g0903(.A(KEYINPUT117), .B1(new_n874), .B2(G330), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n931), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n833), .A2(new_n382), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n732), .A2(new_n697), .A3(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n761), .A2(G330), .A3(new_n879), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1105), .A2(new_n933), .A3(new_n1107), .A4(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n761), .A2(G330), .A3(new_n834), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n931), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n879), .A2(new_n874), .A3(G330), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n932), .A2(new_n933), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1109), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1098), .A2(new_n1116), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n934), .A2(new_n929), .B1(new_n926), .B2(new_n927), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n931), .B1(new_n1107), .B2(new_n933), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n912), .B1(new_n440), .B2(new_n701), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1118), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1112), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1118), .B(new_n1108), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n1117), .A2(KEYINPUT118), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  AND2_X1   g0925(.A1(new_n1125), .A2(new_n1065), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1117), .A2(KEYINPUT118), .A3(new_n1065), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1127), .B1(new_n1128), .B2(new_n971), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n765), .B1(new_n926), .B2(new_n927), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n858), .A2(new_n284), .ZN(new_n1131));
  XOR2_X1   g0931(.A(KEYINPUT54), .B(G143), .Z(new_n1132));
  NAND2_X1  g0932(.A1(new_n842), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n792), .A2(G150), .ZN(new_n1134));
  OR2_X1    g0934(.A1(new_n1134), .A2(KEYINPUT53), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n774), .A2(G137), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n801), .A2(G50), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1133), .A2(new_n1135), .A3(new_n1136), .A4(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(KEYINPUT53), .B2(new_n1134), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(G125), .A2(new_n785), .B1(new_n778), .B2(G159), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n789), .A2(G132), .B1(new_n794), .B2(G128), .ZN(new_n1141));
  XOR2_X1   g0941(.A(new_n1141), .B(KEYINPUT119), .Z(new_n1142));
  NAND4_X1  g0942(.A1(new_n1139), .A2(new_n260), .A3(new_n1140), .A4(new_n1142), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n853), .B1(new_n604), .B2(new_n773), .C1(new_n1047), .C2(new_n784), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n255), .B1(new_n780), .B2(new_n803), .C1(new_n811), .C2(new_n210), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(G116), .B2(new_n789), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1146), .A2(new_n799), .A3(new_n1080), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1143), .B1(new_n1144), .B2(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(new_n1148), .B(KEYINPUT120), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n814), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1130), .A2(new_n816), .A3(new_n1131), .A4(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n1126), .A2(new_n1129), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(G378));
  NOR2_X1   g0954(.A1(new_n405), .A2(new_n883), .ZN(new_n1155));
  AND2_X1   g0955(.A1(new_n409), .A2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n409), .A2(new_n1155), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  OR3_X1    g0959(.A1(new_n1156), .A2(new_n1157), .A3(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1159), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n765), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(KEYINPUT122), .B(G124), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n785), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(new_n295), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n770), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(G137), .A2(new_n1168), .B1(new_n794), .B2(G125), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n789), .A2(G128), .B1(new_n778), .B2(G150), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n792), .A2(new_n1132), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n774), .A2(G132), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .A4(new_n1172), .ZN(new_n1173));
  AOI211_X1 g0973(.A(G33), .B(new_n1167), .C1(new_n1173), .C2(KEYINPUT59), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n1174), .B1(KEYINPUT59), .B2(new_n1173), .C1(new_n848), .C2(new_n782), .ZN(new_n1175));
  AOI21_X1  g0975(.A(G41), .B1(KEYINPUT3), .B2(G33), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1175), .B1(G50), .B2(new_n1176), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(G116), .A2(new_n794), .B1(new_n801), .B2(G58), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1178), .B1(new_n210), .B2(new_n773), .C1(new_n780), .C2(new_n784), .ZN(new_n1179));
  AOI211_X1 g0979(.A(G41), .B(new_n260), .C1(new_n792), .C2(G77), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n577), .B2(new_n770), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n788), .A2(new_n604), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT121), .ZN(new_n1183));
  NOR4_X1   g0983(.A1(new_n1179), .A2(new_n1181), .A3(new_n1183), .A4(new_n960), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1184), .B(KEYINPUT58), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n814), .B1(new_n1177), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n858), .A2(new_n202), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1164), .A2(new_n816), .A3(new_n1186), .A4(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n914), .A2(new_n1163), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1162), .B1(new_n919), .B2(G330), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n938), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n938), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n914), .A2(new_n1163), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n919), .A2(G330), .A3(new_n1162), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1192), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1189), .B1(new_n1197), .B2(new_n972), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1123), .A2(new_n1116), .A3(new_n1124), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n1196), .A2(new_n1192), .B1(new_n1199), .B2(new_n1098), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1065), .B1(new_n1200), .B2(KEYINPUT57), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1199), .A2(new_n1098), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1197), .A2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT57), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1198), .B1(new_n1201), .B2(new_n1205), .ZN(G375));
  OAI21_X1  g1006(.A(KEYINPUT123), .B1(new_n1098), .B2(new_n1116), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n922), .A2(new_n688), .A3(new_n915), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT123), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1208), .A2(new_n1209), .A3(new_n1115), .A4(new_n1109), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1207), .A2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1211), .A2(new_n1010), .A3(new_n1117), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n931), .A2(new_n765), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n774), .A2(new_n1132), .B1(new_n794), .B2(G132), .ZN(new_n1214));
  INV_X1    g1014(.A(G137), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1214), .B1(new_n1215), .B2(new_n788), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n260), .B1(new_n1216), .B2(KEYINPUT124), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(KEYINPUT124), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(G128), .A2(new_n785), .B1(new_n778), .B2(G50), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(G159), .A2(new_n792), .B1(new_n801), .B2(G58), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1217), .B(new_n1221), .C1(G150), .C2(new_n1168), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n533), .A2(new_n774), .B1(new_n792), .B2(G97), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n1223), .B1(new_n780), .B2(new_n788), .C1(new_n1047), .C2(new_n803), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1056), .B1(G77), .B2(new_n801), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1225), .B(new_n255), .C1(new_n604), .C2(new_n811), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n1224), .B(new_n1226), .C1(G303), .C2(new_n785), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n814), .B1(new_n1222), .B2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n858), .A2(new_n806), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1213), .A2(new_n816), .A3(new_n1228), .A4(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(new_n1116), .B2(new_n972), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1212), .A2(new_n1232), .ZN(G381));
  NAND2_X1  g1033(.A1(new_n1197), .A2(new_n972), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n1188), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n717), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1200), .A2(KEYINPUT57), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1235), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  NOR4_X1   g1038(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(G387), .A2(G390), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1238), .A2(new_n1239), .A3(new_n1153), .A4(new_n1240), .ZN(G407));
  NAND2_X1  g1041(.A1(new_n1238), .A2(new_n1153), .ZN(new_n1242));
  OAI211_X1 g1042(.A(G407), .B(G213), .C1(G343), .C2(new_n1242), .ZN(G409));
  NAND2_X1  g1043(.A1(G387), .A2(G390), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n1090), .A2(new_n1092), .B1(new_n1008), .B2(new_n1095), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1245), .B(new_n970), .C1(new_n1011), .C2(new_n1031), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1244), .A2(new_n1246), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(G393), .B(G396), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1247), .A2(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1244), .A2(new_n1246), .A3(new_n1248), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1253), .A2(new_n1237), .A3(new_n1065), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1153), .B1(new_n1254), .B2(new_n1198), .ZN(new_n1255));
  INV_X1    g1055(.A(G384), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1208), .A2(KEYINPUT60), .A3(new_n1115), .A4(new_n1109), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n1065), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1117), .A2(KEYINPUT60), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1258), .B1(new_n1211), .B2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1232), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1256), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n1207), .A2(new_n1210), .B1(new_n1117), .B2(KEYINPUT60), .ZN(new_n1263));
  OAI211_X1 g1063(.A(G384), .B(new_n1232), .C1(new_n1263), .C2(new_n1258), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1262), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1129), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1152), .B1(new_n1125), .B2(new_n1065), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1197), .A2(new_n1202), .A3(new_n1010), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1266), .A2(new_n1198), .A3(new_n1267), .A4(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(G343), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(G213), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1269), .A2(new_n1271), .ZN(new_n1272));
  NOR3_X1   g1072(.A1(new_n1255), .A2(new_n1265), .A3(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT62), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(G375), .A2(G378), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1265), .ZN(new_n1277));
  AND2_X1   g1077(.A1(new_n1269), .A2(new_n1271), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1276), .A2(new_n1277), .A3(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(KEYINPUT62), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT61), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1275), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1270), .A2(KEYINPUT125), .A3(G213), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1262), .A2(new_n1264), .A3(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1270), .A2(G213), .A3(G2897), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1285), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1262), .A2(new_n1264), .A3(new_n1287), .A4(new_n1283), .ZN(new_n1288));
  AOI22_X1  g1088(.A1(new_n1276), .A2(new_n1278), .B1(new_n1286), .B2(new_n1288), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1252), .B1(new_n1282), .B2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT63), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1286), .A2(new_n1288), .ZN(new_n1292));
  OAI211_X1 g1092(.A(new_n1271), .B(new_n1269), .C1(new_n1238), .C2(new_n1153), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1291), .B1(new_n1294), .B2(new_n1279), .ZN(new_n1295));
  AND3_X1   g1095(.A1(new_n1244), .A2(new_n1246), .A3(new_n1248), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1248), .B1(new_n1244), .B2(new_n1246), .ZN(new_n1297));
  NOR3_X1   g1097(.A1(new_n1296), .A2(new_n1297), .A3(KEYINPUT61), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1298), .B1(new_n1273), .B2(KEYINPUT63), .ZN(new_n1299));
  NOR3_X1   g1099(.A1(new_n1295), .A2(new_n1299), .A3(KEYINPUT126), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT126), .ZN(new_n1301));
  OAI21_X1  g1101(.A(KEYINPUT63), .B1(new_n1289), .B2(new_n1273), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1250), .A2(new_n1281), .A3(new_n1251), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1303), .B1(new_n1279), .B2(new_n1291), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1301), .B1(new_n1302), .B2(new_n1304), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1290), .B1(new_n1300), .B2(new_n1305), .ZN(G405));
  NAND2_X1  g1106(.A1(new_n1242), .A2(new_n1276), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1277), .A2(KEYINPUT127), .ZN(new_n1308));
  XNOR2_X1  g1108(.A(new_n1307), .B(new_n1308), .ZN(new_n1309));
  XNOR2_X1  g1109(.A(new_n1309), .B(new_n1252), .ZN(G402));
endmodule


