

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583;

  NOR2_X1 U324 ( .A1(n538), .A2(n514), .ZN(n465) );
  XNOR2_X1 U325 ( .A(n405), .B(n293), .ZN(n317) );
  XNOR2_X1 U326 ( .A(n384), .B(n383), .ZN(n391) );
  XNOR2_X1 U327 ( .A(n322), .B(n321), .ZN(n514) );
  XOR2_X1 U328 ( .A(KEYINPUT92), .B(KEYINPUT21), .Z(n292) );
  AND2_X1 U329 ( .A1(G226GAT), .A2(G233GAT), .ZN(n293) );
  XOR2_X1 U330 ( .A(n440), .B(n439), .Z(n294) );
  XNOR2_X1 U331 ( .A(KEYINPUT45), .B(KEYINPUT65), .ZN(n456) );
  XNOR2_X1 U332 ( .A(n457), .B(n456), .ZN(n459) );
  NOR2_X1 U333 ( .A1(n563), .A2(n454), .ZN(n455) );
  INV_X1 U334 ( .A(KEYINPUT102), .ZN(n371) );
  XNOR2_X1 U335 ( .A(n441), .B(n294), .ZN(n442) );
  XNOR2_X1 U336 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U337 ( .A(n372), .B(n371), .ZN(n478) );
  XNOR2_X1 U338 ( .A(n443), .B(n442), .ZN(n444) );
  OR2_X1 U339 ( .A1(n364), .A2(n512), .ZN(n343) );
  XNOR2_X1 U340 ( .A(n464), .B(KEYINPUT48), .ZN(n538) );
  XNOR2_X1 U341 ( .A(n343), .B(KEYINPUT99), .ZN(n540) );
  NOR2_X1 U342 ( .A1(n567), .A2(n566), .ZN(n581) );
  INV_X1 U343 ( .A(G169GAT), .ZN(n471) );
  XNOR2_X1 U344 ( .A(KEYINPUT41), .B(n575), .ZN(n545) );
  INV_X1 U345 ( .A(G43GAT), .ZN(n447) );
  XNOR2_X1 U346 ( .A(n315), .B(n321), .ZN(n524) );
  XNOR2_X1 U347 ( .A(n471), .B(KEYINPUT123), .ZN(n472) );
  XNOR2_X1 U348 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U349 ( .A(n473), .B(n472), .ZN(G1348GAT) );
  XNOR2_X1 U350 ( .A(n450), .B(n449), .ZN(G1330GAT) );
  XOR2_X1 U351 ( .A(KEYINPUT84), .B(KEYINPUT0), .Z(n296) );
  XNOR2_X1 U352 ( .A(G113GAT), .B(G134GAT), .ZN(n295) );
  XNOR2_X1 U353 ( .A(n296), .B(n295), .ZN(n329) );
  XOR2_X1 U354 ( .A(G15GAT), .B(G127GAT), .Z(n393) );
  XOR2_X1 U355 ( .A(n329), .B(n393), .Z(n298) );
  XNOR2_X1 U356 ( .A(G43GAT), .B(G99GAT), .ZN(n297) );
  XNOR2_X1 U357 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U358 ( .A(KEYINPUT20), .B(KEYINPUT85), .Z(n300) );
  NAND2_X1 U359 ( .A1(G227GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U360 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U361 ( .A(n302), .B(n301), .Z(n307) );
  XOR2_X1 U362 ( .A(KEYINPUT89), .B(KEYINPUT88), .Z(n304) );
  XNOR2_X1 U363 ( .A(G71GAT), .B(G120GAT), .ZN(n303) );
  XNOR2_X1 U364 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U365 ( .A(n305), .B(KEYINPUT90), .ZN(n306) );
  XNOR2_X1 U366 ( .A(n307), .B(n306), .ZN(n315) );
  XOR2_X1 U367 ( .A(KEYINPUT87), .B(KEYINPUT17), .Z(n309) );
  XNOR2_X1 U368 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n308) );
  XNOR2_X1 U369 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U370 ( .A(n310), .B(KEYINPUT86), .Z(n312) );
  XNOR2_X1 U371 ( .A(G190GAT), .B(G183GAT), .ZN(n311) );
  XNOR2_X1 U372 ( .A(n312), .B(n311), .ZN(n314) );
  XOR2_X1 U373 ( .A(G169GAT), .B(G176GAT), .Z(n313) );
  XNOR2_X1 U374 ( .A(n314), .B(n313), .ZN(n321) );
  XNOR2_X1 U375 ( .A(G197GAT), .B(G218GAT), .ZN(n316) );
  XNOR2_X1 U376 ( .A(n292), .B(n316), .ZN(n344) );
  XOR2_X1 U377 ( .A(G8GAT), .B(G211GAT), .Z(n405) );
  XNOR2_X1 U378 ( .A(n344), .B(n317), .ZN(n318) );
  XOR2_X1 U379 ( .A(n318), .B(G204GAT), .Z(n320) );
  XOR2_X1 U380 ( .A(G92GAT), .B(G64GAT), .Z(n431) );
  XNOR2_X1 U381 ( .A(G36GAT), .B(n431), .ZN(n319) );
  XNOR2_X1 U382 ( .A(n320), .B(n319), .ZN(n322) );
  XNOR2_X1 U383 ( .A(n514), .B(KEYINPUT98), .ZN(n323) );
  XNOR2_X1 U384 ( .A(n323), .B(KEYINPUT27), .ZN(n364) );
  XOR2_X1 U385 ( .A(KEYINPUT4), .B(KEYINPUT1), .Z(n325) );
  NAND2_X1 U386 ( .A1(G225GAT), .A2(G233GAT), .ZN(n324) );
  XNOR2_X1 U387 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U388 ( .A(n326), .B(KEYINPUT95), .Z(n331) );
  XOR2_X1 U389 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n328) );
  XNOR2_X1 U390 ( .A(G141GAT), .B(G162GAT), .ZN(n327) );
  XNOR2_X1 U391 ( .A(n328), .B(n327), .ZN(n355) );
  XNOR2_X1 U392 ( .A(n329), .B(n355), .ZN(n330) );
  XNOR2_X1 U393 ( .A(n331), .B(n330), .ZN(n342) );
  XOR2_X1 U394 ( .A(KEYINPUT6), .B(KEYINPUT5), .Z(n333) );
  XNOR2_X1 U395 ( .A(KEYINPUT94), .B(KEYINPUT96), .ZN(n332) );
  XNOR2_X1 U396 ( .A(n333), .B(n332), .ZN(n340) );
  XOR2_X1 U397 ( .A(G155GAT), .B(G57GAT), .Z(n335) );
  XNOR2_X1 U398 ( .A(G1GAT), .B(G127GAT), .ZN(n334) );
  XNOR2_X1 U399 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U400 ( .A(n336), .B(G85GAT), .Z(n338) );
  XOR2_X1 U401 ( .A(G120GAT), .B(G148GAT), .Z(n438) );
  XNOR2_X1 U402 ( .A(G29GAT), .B(n438), .ZN(n337) );
  XNOR2_X1 U403 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U404 ( .A(n340), .B(n339), .Z(n341) );
  XNOR2_X1 U405 ( .A(n342), .B(n341), .ZN(n368) );
  XNOR2_X1 U406 ( .A(KEYINPUT97), .B(n368), .ZN(n512) );
  XOR2_X1 U407 ( .A(KEYINPUT93), .B(n344), .Z(n346) );
  NAND2_X1 U408 ( .A1(G228GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U409 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U410 ( .A(G22GAT), .B(G155GAT), .Z(n392) );
  XOR2_X1 U411 ( .A(n347), .B(n392), .Z(n349) );
  XNOR2_X1 U412 ( .A(G50GAT), .B(G211GAT), .ZN(n348) );
  XNOR2_X1 U413 ( .A(n349), .B(n348), .ZN(n353) );
  XOR2_X1 U414 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n351) );
  XNOR2_X1 U415 ( .A(G148GAT), .B(KEYINPUT24), .ZN(n350) );
  XNOR2_X1 U416 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U417 ( .A(n353), .B(n352), .Z(n357) );
  XNOR2_X1 U418 ( .A(G204GAT), .B(G106GAT), .ZN(n354) );
  XNOR2_X1 U419 ( .A(n354), .B(G78GAT), .ZN(n429) );
  XNOR2_X1 U420 ( .A(n355), .B(n429), .ZN(n356) );
  XNOR2_X1 U421 ( .A(n357), .B(n356), .ZN(n468) );
  XOR2_X1 U422 ( .A(n468), .B(KEYINPUT28), .Z(n520) );
  NAND2_X1 U423 ( .A1(n540), .A2(n520), .ZN(n523) );
  XNOR2_X1 U424 ( .A(KEYINPUT91), .B(n524), .ZN(n358) );
  NOR2_X1 U425 ( .A1(n523), .A2(n358), .ZN(n370) );
  NOR2_X1 U426 ( .A1(n524), .A2(n514), .ZN(n359) );
  XOR2_X1 U427 ( .A(KEYINPUT101), .B(n359), .Z(n360) );
  NOR2_X1 U428 ( .A1(n468), .A2(n360), .ZN(n361) );
  XOR2_X1 U429 ( .A(KEYINPUT25), .B(n361), .Z(n366) );
  NAND2_X1 U430 ( .A1(n468), .A2(n524), .ZN(n362) );
  XNOR2_X1 U431 ( .A(n362), .B(KEYINPUT100), .ZN(n363) );
  XNOR2_X1 U432 ( .A(n363), .B(KEYINPUT26), .ZN(n566) );
  NOR2_X1 U433 ( .A1(n364), .A2(n566), .ZN(n365) );
  NOR2_X1 U434 ( .A1(n366), .A2(n365), .ZN(n367) );
  NOR2_X1 U435 ( .A1(n368), .A2(n367), .ZN(n369) );
  NOR2_X1 U436 ( .A1(n370), .A2(n369), .ZN(n372) );
  XOR2_X1 U437 ( .A(KEYINPUT66), .B(KEYINPUT10), .Z(n374) );
  XNOR2_X1 U438 ( .A(KEYINPUT11), .B(KEYINPUT76), .ZN(n373) );
  XNOR2_X1 U439 ( .A(n374), .B(n373), .ZN(n378) );
  XOR2_X1 U440 ( .A(G99GAT), .B(G85GAT), .Z(n432) );
  XNOR2_X1 U441 ( .A(G218GAT), .B(n432), .ZN(n376) );
  XOR2_X1 U442 ( .A(G106GAT), .B(KEYINPUT9), .Z(n375) );
  XNOR2_X1 U443 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U444 ( .A(n378), .B(n377), .ZN(n384) );
  XOR2_X1 U445 ( .A(G92GAT), .B(G162GAT), .Z(n380) );
  XNOR2_X1 U446 ( .A(G190GAT), .B(G134GAT), .ZN(n379) );
  XNOR2_X1 U447 ( .A(n380), .B(n379), .ZN(n382) );
  AND2_X1 U448 ( .A1(G232GAT), .A2(G233GAT), .ZN(n381) );
  XOR2_X1 U449 ( .A(G29GAT), .B(G36GAT), .Z(n386) );
  XNOR2_X1 U450 ( .A(G50GAT), .B(G43GAT), .ZN(n385) );
  XNOR2_X1 U451 ( .A(n386), .B(n385), .ZN(n390) );
  XOR2_X1 U452 ( .A(KEYINPUT68), .B(KEYINPUT8), .Z(n388) );
  XNOR2_X1 U453 ( .A(KEYINPUT67), .B(KEYINPUT7), .ZN(n387) );
  XNOR2_X1 U454 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U455 ( .A(n390), .B(n389), .ZN(n428) );
  XNOR2_X1 U456 ( .A(n391), .B(n428), .ZN(n563) );
  XNOR2_X1 U457 ( .A(KEYINPUT36), .B(n563), .ZN(n580) );
  NAND2_X1 U458 ( .A1(n478), .A2(n580), .ZN(n413) );
  XNOR2_X1 U459 ( .A(KEYINPUT81), .B(n392), .ZN(n395) );
  XNOR2_X1 U460 ( .A(n393), .B(G78GAT), .ZN(n394) );
  XNOR2_X1 U461 ( .A(n395), .B(n394), .ZN(n399) );
  XOR2_X1 U462 ( .A(KEYINPUT77), .B(KEYINPUT78), .Z(n397) );
  XNOR2_X1 U463 ( .A(KEYINPUT12), .B(KEYINPUT15), .ZN(n396) );
  XNOR2_X1 U464 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U465 ( .A(n399), .B(n398), .ZN(n401) );
  XNOR2_X1 U466 ( .A(G183GAT), .B(G64GAT), .ZN(n400) );
  XNOR2_X1 U467 ( .A(n401), .B(n400), .ZN(n404) );
  XOR2_X1 U468 ( .A(KEYINPUT13), .B(KEYINPUT71), .Z(n403) );
  XNOR2_X1 U469 ( .A(G71GAT), .B(G57GAT), .ZN(n402) );
  XNOR2_X1 U470 ( .A(n403), .B(n402), .ZN(n430) );
  XNOR2_X1 U471 ( .A(n404), .B(n430), .ZN(n407) );
  XOR2_X1 U472 ( .A(KEYINPUT69), .B(G1GAT), .Z(n417) );
  XOR2_X1 U473 ( .A(n417), .B(n405), .Z(n406) );
  XNOR2_X1 U474 ( .A(n407), .B(n406), .ZN(n412) );
  XOR2_X1 U475 ( .A(KEYINPUT14), .B(KEYINPUT80), .Z(n409) );
  NAND2_X1 U476 ( .A1(G231GAT), .A2(G233GAT), .ZN(n408) );
  XNOR2_X1 U477 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U478 ( .A(KEYINPUT79), .B(n410), .ZN(n411) );
  XNOR2_X1 U479 ( .A(n412), .B(n411), .ZN(n578) );
  NOR2_X1 U480 ( .A1(n413), .A2(n578), .ZN(n414) );
  XNOR2_X1 U481 ( .A(n414), .B(KEYINPUT37), .ZN(n511) );
  XOR2_X1 U482 ( .A(KEYINPUT70), .B(G141GAT), .Z(n416) );
  NAND2_X1 U483 ( .A1(G229GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U484 ( .A(n416), .B(n415), .ZN(n418) );
  XOR2_X1 U485 ( .A(n418), .B(n417), .Z(n426) );
  XOR2_X1 U486 ( .A(KEYINPUT30), .B(G8GAT), .Z(n420) );
  XNOR2_X1 U487 ( .A(G169GAT), .B(G197GAT), .ZN(n419) );
  XNOR2_X1 U488 ( .A(n420), .B(n419), .ZN(n424) );
  XOR2_X1 U489 ( .A(G22GAT), .B(G113GAT), .Z(n422) );
  XNOR2_X1 U490 ( .A(KEYINPUT29), .B(G15GAT), .ZN(n421) );
  XNOR2_X1 U491 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U492 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U493 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U494 ( .A(n428), .B(n427), .ZN(n568) );
  XNOR2_X1 U495 ( .A(n430), .B(n429), .ZN(n445) );
  XOR2_X1 U496 ( .A(n432), .B(n431), .Z(n434) );
  NAND2_X1 U497 ( .A1(G230GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U498 ( .A(n434), .B(n433), .ZN(n443) );
  XOR2_X1 U499 ( .A(KEYINPUT31), .B(KEYINPUT73), .Z(n436) );
  XNOR2_X1 U500 ( .A(G176GAT), .B(KEYINPUT32), .ZN(n435) );
  XNOR2_X1 U501 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U502 ( .A(n438), .B(n437), .ZN(n441) );
  XOR2_X1 U503 ( .A(KEYINPUT72), .B(KEYINPUT75), .Z(n440) );
  XNOR2_X1 U504 ( .A(KEYINPUT33), .B(KEYINPUT74), .ZN(n439) );
  XNOR2_X1 U505 ( .A(n445), .B(n444), .ZN(n458) );
  NAND2_X1 U506 ( .A1(n568), .A2(n458), .ZN(n479) );
  NOR2_X1 U507 ( .A1(n511), .A2(n479), .ZN(n446) );
  XOR2_X1 U508 ( .A(KEYINPUT38), .B(n446), .Z(n495) );
  NOR2_X1 U509 ( .A1(n524), .A2(n495), .ZN(n450) );
  XNOR2_X1 U510 ( .A(KEYINPUT108), .B(KEYINPUT40), .ZN(n448) );
  XOR2_X1 U511 ( .A(KEYINPUT46), .B(KEYINPUT117), .Z(n452) );
  INV_X1 U512 ( .A(n458), .ZN(n575) );
  INV_X1 U513 ( .A(n545), .ZN(n553) );
  NAND2_X1 U514 ( .A1(n568), .A2(n553), .ZN(n451) );
  XNOR2_X1 U515 ( .A(n452), .B(n451), .ZN(n453) );
  INV_X1 U516 ( .A(n578), .ZN(n548) );
  XNOR2_X1 U517 ( .A(KEYINPUT116), .B(n548), .ZN(n559) );
  NAND2_X1 U518 ( .A1(n453), .A2(n559), .ZN(n454) );
  XOR2_X1 U519 ( .A(n455), .B(KEYINPUT47), .Z(n463) );
  NAND2_X1 U520 ( .A1(n578), .A2(n580), .ZN(n457) );
  NAND2_X1 U521 ( .A1(n459), .A2(n458), .ZN(n460) );
  NOR2_X1 U522 ( .A1(n568), .A2(n460), .ZN(n461) );
  XNOR2_X1 U523 ( .A(KEYINPUT118), .B(n461), .ZN(n462) );
  NOR2_X1 U524 ( .A1(n463), .A2(n462), .ZN(n464) );
  XNOR2_X1 U525 ( .A(KEYINPUT54), .B(n465), .ZN(n466) );
  NAND2_X1 U526 ( .A1(n466), .A2(n512), .ZN(n467) );
  XNOR2_X1 U527 ( .A(n467), .B(KEYINPUT64), .ZN(n567) );
  NOR2_X1 U528 ( .A1(n567), .A2(n468), .ZN(n469) );
  XNOR2_X1 U529 ( .A(n469), .B(KEYINPUT55), .ZN(n470) );
  NOR2_X2 U530 ( .A1(n524), .A2(n470), .ZN(n562) );
  NAND2_X1 U531 ( .A1(n562), .A2(n568), .ZN(n473) );
  NOR2_X1 U532 ( .A1(n563), .A2(n548), .ZN(n475) );
  XNOR2_X1 U533 ( .A(KEYINPUT16), .B(KEYINPUT83), .ZN(n474) );
  XNOR2_X1 U534 ( .A(n475), .B(n474), .ZN(n476) );
  XOR2_X1 U535 ( .A(KEYINPUT82), .B(n476), .Z(n477) );
  NAND2_X1 U536 ( .A1(n478), .A2(n477), .ZN(n497) );
  NOR2_X1 U537 ( .A1(n497), .A2(n479), .ZN(n480) );
  XNOR2_X1 U538 ( .A(n480), .B(KEYINPUT103), .ZN(n487) );
  NOR2_X1 U539 ( .A1(n512), .A2(n487), .ZN(n481) );
  XOR2_X1 U540 ( .A(KEYINPUT34), .B(n481), .Z(n482) );
  XNOR2_X1 U541 ( .A(G1GAT), .B(n482), .ZN(G1324GAT) );
  NOR2_X1 U542 ( .A1(n514), .A2(n487), .ZN(n483) );
  XOR2_X1 U543 ( .A(G8GAT), .B(n483), .Z(G1325GAT) );
  NOR2_X1 U544 ( .A1(n524), .A2(n487), .ZN(n485) );
  XNOR2_X1 U545 ( .A(KEYINPUT104), .B(KEYINPUT35), .ZN(n484) );
  XNOR2_X1 U546 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U547 ( .A(G15GAT), .B(n486), .ZN(G1326GAT) );
  NOR2_X1 U548 ( .A1(n520), .A2(n487), .ZN(n489) );
  XNOR2_X1 U549 ( .A(G22GAT), .B(KEYINPUT105), .ZN(n488) );
  XNOR2_X1 U550 ( .A(n489), .B(n488), .ZN(G1327GAT) );
  NOR2_X1 U551 ( .A1(n495), .A2(n512), .ZN(n493) );
  XOR2_X1 U552 ( .A(KEYINPUT106), .B(KEYINPUT39), .Z(n491) );
  XNOR2_X1 U553 ( .A(G29GAT), .B(KEYINPUT107), .ZN(n490) );
  XNOR2_X1 U554 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U555 ( .A(n493), .B(n492), .ZN(G1328GAT) );
  NOR2_X1 U556 ( .A1(n514), .A2(n495), .ZN(n494) );
  XOR2_X1 U557 ( .A(G36GAT), .B(n494), .Z(G1329GAT) );
  NOR2_X1 U558 ( .A1(n520), .A2(n495), .ZN(n496) );
  XOR2_X1 U559 ( .A(G50GAT), .B(n496), .Z(G1331GAT) );
  INV_X1 U560 ( .A(n568), .ZN(n541) );
  NAND2_X1 U561 ( .A1(n541), .A2(n553), .ZN(n510) );
  NOR2_X1 U562 ( .A1(n510), .A2(n497), .ZN(n498) );
  XNOR2_X1 U563 ( .A(n498), .B(KEYINPUT109), .ZN(n505) );
  NOR2_X1 U564 ( .A1(n512), .A2(n505), .ZN(n499) );
  XOR2_X1 U565 ( .A(KEYINPUT42), .B(n499), .Z(n500) );
  XNOR2_X1 U566 ( .A(G57GAT), .B(n500), .ZN(G1332GAT) );
  NOR2_X1 U567 ( .A1(n514), .A2(n505), .ZN(n501) );
  XOR2_X1 U568 ( .A(KEYINPUT110), .B(n501), .Z(n502) );
  XNOR2_X1 U569 ( .A(G64GAT), .B(n502), .ZN(G1333GAT) );
  NOR2_X1 U570 ( .A1(n524), .A2(n505), .ZN(n504) );
  XNOR2_X1 U571 ( .A(G71GAT), .B(KEYINPUT111), .ZN(n503) );
  XNOR2_X1 U572 ( .A(n504), .B(n503), .ZN(G1334GAT) );
  NOR2_X1 U573 ( .A1(n505), .A2(n520), .ZN(n509) );
  XOR2_X1 U574 ( .A(KEYINPUT112), .B(KEYINPUT43), .Z(n507) );
  XNOR2_X1 U575 ( .A(G78GAT), .B(KEYINPUT113), .ZN(n506) );
  XNOR2_X1 U576 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U577 ( .A(n509), .B(n508), .ZN(G1335GAT) );
  OR2_X1 U578 ( .A1(n511), .A2(n510), .ZN(n519) );
  NOR2_X1 U579 ( .A1(n512), .A2(n519), .ZN(n513) );
  XOR2_X1 U580 ( .A(G85GAT), .B(n513), .Z(G1336GAT) );
  NOR2_X1 U581 ( .A1(n514), .A2(n519), .ZN(n515) );
  XOR2_X1 U582 ( .A(G92GAT), .B(n515), .Z(G1337GAT) );
  NOR2_X1 U583 ( .A1(n524), .A2(n519), .ZN(n517) );
  XNOR2_X1 U584 ( .A(KEYINPUT114), .B(KEYINPUT115), .ZN(n516) );
  XNOR2_X1 U585 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U586 ( .A(G99GAT), .B(n518), .ZN(G1338GAT) );
  NOR2_X1 U587 ( .A1(n520), .A2(n519), .ZN(n521) );
  XOR2_X1 U588 ( .A(KEYINPUT44), .B(n521), .Z(n522) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(n522), .ZN(G1339GAT) );
  NOR2_X1 U590 ( .A1(n538), .A2(n523), .ZN(n526) );
  INV_X1 U591 ( .A(n524), .ZN(n525) );
  NAND2_X1 U592 ( .A1(n526), .A2(n525), .ZN(n535) );
  NOR2_X1 U593 ( .A1(n541), .A2(n535), .ZN(n528) );
  XNOR2_X1 U594 ( .A(G113GAT), .B(KEYINPUT119), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n528), .B(n527), .ZN(G1340GAT) );
  NOR2_X1 U596 ( .A1(n545), .A2(n535), .ZN(n530) );
  XNOR2_X1 U597 ( .A(KEYINPUT49), .B(KEYINPUT120), .ZN(n529) );
  XNOR2_X1 U598 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U599 ( .A(G120GAT), .B(n531), .ZN(G1341GAT) );
  NOR2_X1 U600 ( .A1(n559), .A2(n535), .ZN(n533) );
  XNOR2_X1 U601 ( .A(KEYINPUT50), .B(KEYINPUT121), .ZN(n532) );
  XNOR2_X1 U602 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U603 ( .A(G127GAT), .B(n534), .ZN(G1342GAT) );
  INV_X1 U604 ( .A(n563), .ZN(n551) );
  NOR2_X1 U605 ( .A1(n551), .A2(n535), .ZN(n537) );
  XNOR2_X1 U606 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n536) );
  XNOR2_X1 U607 ( .A(n537), .B(n536), .ZN(G1343GAT) );
  NOR2_X1 U608 ( .A1(n538), .A2(n566), .ZN(n539) );
  NAND2_X1 U609 ( .A1(n540), .A2(n539), .ZN(n550) );
  NOR2_X1 U610 ( .A1(n541), .A2(n550), .ZN(n542) );
  XOR2_X1 U611 ( .A(G141GAT), .B(n542), .Z(G1344GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT122), .B(KEYINPUT52), .Z(n544) );
  XNOR2_X1 U613 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n543) );
  XNOR2_X1 U614 ( .A(n544), .B(n543), .ZN(n547) );
  NOR2_X1 U615 ( .A1(n545), .A2(n550), .ZN(n546) );
  XOR2_X1 U616 ( .A(n547), .B(n546), .Z(G1345GAT) );
  NOR2_X1 U617 ( .A1(n548), .A2(n550), .ZN(n549) );
  XOR2_X1 U618 ( .A(G155GAT), .B(n549), .Z(G1346GAT) );
  NOR2_X1 U619 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U620 ( .A(G162GAT), .B(n552), .Z(G1347GAT) );
  XNOR2_X1 U621 ( .A(G176GAT), .B(KEYINPUT124), .ZN(n557) );
  XOR2_X1 U622 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n555) );
  NAND2_X1 U623 ( .A1(n562), .A2(n553), .ZN(n554) );
  XNOR2_X1 U624 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U625 ( .A(n557), .B(n556), .ZN(G1349GAT) );
  INV_X1 U626 ( .A(n562), .ZN(n558) );
  NOR2_X1 U627 ( .A1(n559), .A2(n558), .ZN(n561) );
  XNOR2_X1 U628 ( .A(G183GAT), .B(KEYINPUT125), .ZN(n560) );
  XNOR2_X1 U629 ( .A(n561), .B(n560), .ZN(G1350GAT) );
  NAND2_X1 U630 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n564), .B(KEYINPUT58), .ZN(n565) );
  XNOR2_X1 U632 ( .A(G190GAT), .B(n565), .ZN(G1351GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT127), .B(KEYINPUT60), .Z(n570) );
  NAND2_X1 U634 ( .A1(n581), .A2(n568), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n571), .B(KEYINPUT59), .ZN(n572) );
  INV_X1 U637 ( .A(n572), .ZN(n574) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  XOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT61), .Z(n577) );
  NAND2_X1 U641 ( .A1(n581), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  NAND2_X1 U643 ( .A1(n581), .A2(n578), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n579), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U646 ( .A(n582), .B(KEYINPUT62), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

