

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812;

  AND2_X1 U370 ( .A1(n408), .A2(n494), .ZN(n349) );
  INV_X2 U371 ( .A(G953), .ZN(n795) );
  XNOR2_X2 U372 ( .A(n671), .B(KEYINPUT59), .ZN(n672) );
  XNOR2_X2 U373 ( .A(KEYINPUT76), .B(KEYINPUT22), .ZN(n634) );
  XNOR2_X2 U374 ( .A(n591), .B(n590), .ZN(n810) );
  AND2_X2 U375 ( .A1(n645), .A2(KEYINPUT106), .ZN(n422) );
  OR2_X2 U376 ( .A1(n700), .A2(G902), .ZN(n539) );
  NAND2_X2 U377 ( .A1(n459), .A2(n406), .ZN(n460) );
  XNOR2_X2 U378 ( .A(n460), .B(n498), .ZN(n811) );
  NOR2_X1 U379 ( .A1(n651), .A2(n592), .ZN(n589) );
  BUF_X1 U380 ( .A(G146), .Z(n355) );
  OR2_X1 U381 ( .A1(n785), .A2(n351), .ZN(n346) );
  AND2_X2 U382 ( .A1(n496), .A2(n492), .ZN(n459) );
  AND2_X2 U383 ( .A1(n398), .A2(n467), .ZN(n399) );
  OR2_X2 U384 ( .A1(n722), .A2(n425), .ZN(n467) );
  XNOR2_X2 U385 ( .A(n452), .B(n624), .ZN(n768) );
  NOR2_X2 U386 ( .A1(n811), .A2(n810), .ZN(n445) );
  XNOR2_X2 U387 ( .A(n350), .B(n499), .ZN(n417) );
  INV_X1 U388 ( .A(n786), .ZN(n789) );
  XNOR2_X1 U389 ( .A(KEYINPUT68), .B(G101), .ZN(n545) );
  NOR2_X1 U390 ( .A1(n787), .A2(n753), .ZN(n607) );
  XNOR2_X1 U391 ( .A(n461), .B(n524), .ZN(n738) );
  INV_X1 U392 ( .A(KEYINPUT47), .ZN(n352) );
  INV_X1 U393 ( .A(KEYINPUT28), .ZN(n354) );
  NOR2_X1 U394 ( .A1(n346), .A2(n808), .ZN(n444) );
  AND2_X1 U395 ( .A1(n644), .A2(n383), .ZN(n359) );
  XNOR2_X1 U396 ( .A(n437), .B(n632), .ZN(n686) );
  AND2_X1 U397 ( .A1(n432), .A2(n394), .ZN(n430) );
  XNOR2_X1 U398 ( .A(n418), .B(KEYINPUT115), .ZN(n808) );
  BUF_X1 U399 ( .A(n643), .Z(n382) );
  AND2_X1 U400 ( .A1(n449), .A2(n451), .ZN(n448) );
  XNOR2_X1 U401 ( .A(n722), .B(n721), .ZN(n723) );
  INV_X1 U402 ( .A(n738), .ZN(n347) );
  BUF_X2 U403 ( .A(n720), .Z(n722) );
  INV_X1 U404 ( .A(n739), .ZN(n348) );
  INV_X1 U405 ( .A(n355), .ZN(n487) );
  NAND2_X1 U406 ( .A1(n349), .A2(n409), .ZN(n406) );
  NAND2_X1 U407 ( .A1(n443), .A2(n444), .ZN(n350) );
  AND2_X1 U408 ( .A1(n738), .A2(n348), .ZN(n588) );
  XNOR2_X1 U409 ( .A(n607), .B(n352), .ZN(n351) );
  OR2_X1 U410 ( .A1(n353), .A2(n597), .ZN(n604) );
  XNOR2_X1 U411 ( .A(n589), .B(n354), .ZN(n353) );
  NAND2_X1 U412 ( .A1(n347), .A2(n348), .ZN(n735) );
  NAND2_X1 U413 ( .A1(n399), .A2(n356), .ZN(n603) );
  NAND2_X1 U414 ( .A1(n358), .A2(n357), .ZN(n356) );
  INV_X1 U415 ( .A(n400), .ZN(n357) );
  INV_X1 U416 ( .A(n468), .ZN(n358) );
  NOR2_X1 U417 ( .A1(n478), .A2(n757), .ZN(n477) );
  XNOR2_X1 U418 ( .A(n593), .B(n559), .ZN(n752) );
  INV_X1 U419 ( .A(KEYINPUT89), .ZN(n647) );
  XNOR2_X1 U420 ( .A(KEYINPUT83), .B(KEYINPUT17), .ZN(n547) );
  NOR2_X1 U421 ( .A1(n371), .A2(KEYINPUT105), .ZN(n450) );
  INV_X1 U422 ( .A(KEYINPUT44), .ZN(n403) );
  INV_X1 U423 ( .A(KEYINPUT90), .ZN(n424) );
  INV_X1 U424 ( .A(G137), .ZN(n504) );
  XNOR2_X1 U425 ( .A(n362), .B(n521), .ZN(n688) );
  XNOR2_X1 U426 ( .A(G134), .B(G122), .ZN(n573) );
  XOR2_X1 U427 ( .A(G131), .B(KEYINPUT71), .Z(n560) );
  XOR2_X1 U428 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n562) );
  XOR2_X1 U429 ( .A(G122), .B(G104), .Z(n565) );
  XNOR2_X1 U430 ( .A(G113), .B(G143), .ZN(n567) );
  XNOR2_X1 U431 ( .A(n688), .B(n487), .ZN(n563) );
  XNOR2_X1 U432 ( .A(n667), .B(KEYINPUT67), .ZN(n668) );
  NAND2_X1 U433 ( .A1(n421), .A2(n364), .ZN(n396) );
  NOR2_X1 U434 ( .A1(n423), .A2(n422), .ZN(n421) );
  NAND2_X1 U435 ( .A1(n592), .A2(KEYINPUT106), .ZN(n454) );
  OR2_X1 U436 ( .A1(n480), .A2(KEYINPUT92), .ZN(n425) );
  XNOR2_X1 U437 ( .A(G119), .B(G116), .ZN(n473) );
  XNOR2_X1 U438 ( .A(n586), .B(KEYINPUT41), .ZN(n767) );
  NOR2_X1 U439 ( .A1(n493), .A2(n786), .ZN(n492) );
  AND2_X1 U440 ( .A1(n540), .A2(n411), .ZN(n410) );
  NAND2_X1 U441 ( .A1(n413), .A2(n412), .ZN(n411) );
  XNOR2_X1 U442 ( .A(n466), .B(n464), .ZN(n606) );
  XNOR2_X1 U443 ( .A(n571), .B(n465), .ZN(n464) );
  NOR2_X1 U444 ( .A1(n671), .A2(G902), .ZN(n466) );
  INV_X1 U445 ( .A(G475), .ZN(n465) );
  INV_X1 U446 ( .A(n382), .ZN(n427) );
  NOR2_X1 U447 ( .A1(n646), .A2(n647), .ZN(n436) );
  NAND2_X1 U448 ( .A1(n427), .A2(n426), .ZN(n432) );
  AND2_X1 U449 ( .A1(n436), .A2(KEYINPUT103), .ZN(n426) );
  INV_X1 U450 ( .A(KEYINPUT103), .ZN(n429) );
  XNOR2_X1 U451 ( .A(KEYINPUT15), .B(G902), .ZN(n662) );
  XNOR2_X1 U452 ( .A(KEYINPUT18), .B(G125), .ZN(n548) );
  NAND2_X1 U453 ( .A1(n448), .A2(n446), .ZN(n453) );
  NAND2_X1 U454 ( .A1(n447), .A2(n450), .ZN(n446) );
  NAND2_X1 U455 ( .A1(n371), .A2(KEYINPUT105), .ZN(n451) );
  NAND2_X1 U456 ( .A1(n481), .A2(n662), .ZN(n480) );
  INV_X1 U457 ( .A(n558), .ZN(n481) );
  INV_X1 U458 ( .A(G902), .ZN(n582) );
  XNOR2_X1 U459 ( .A(n462), .B(KEYINPUT79), .ZN(n564) );
  NAND2_X1 U460 ( .A1(n795), .A2(n463), .ZN(n462) );
  NAND2_X1 U461 ( .A1(n359), .A2(n403), .ZN(n402) );
  INV_X1 U462 ( .A(n587), .ZN(n413) );
  INV_X1 U463 ( .A(KEYINPUT81), .ZN(n412) );
  XNOR2_X1 U464 ( .A(n393), .B(n392), .ZN(n540) );
  INV_X1 U465 ( .A(KEYINPUT30), .ZN(n392) );
  INV_X1 U466 ( .A(KEYINPUT94), .ZN(n405) );
  XNOR2_X1 U467 ( .A(n441), .B(n501), .ZN(n440) );
  XNOR2_X1 U468 ( .A(G134), .B(G131), .ZN(n501) );
  XNOR2_X1 U469 ( .A(n504), .B(KEYINPUT71), .ZN(n441) );
  INV_X1 U470 ( .A(G104), .ZN(n506) );
  XNOR2_X1 U471 ( .A(G110), .B(G107), .ZN(n507) );
  INV_X1 U472 ( .A(KEYINPUT8), .ZN(n519) );
  XNOR2_X1 U473 ( .A(G116), .B(G107), .ZN(n572) );
  XNOR2_X1 U474 ( .A(n570), .B(n569), .ZN(n671) );
  NAND2_X1 U475 ( .A1(G234), .A2(G237), .ZN(n529) );
  XNOR2_X1 U476 ( .A(n396), .B(KEYINPUT113), .ZN(n500) );
  BUF_X1 U477 ( .A(n347), .Z(n395) );
  INV_X1 U478 ( .A(KEYINPUT97), .ZN(n527) );
  XNOR2_X1 U479 ( .A(KEYINPUT78), .B(KEYINPUT16), .ZN(n542) );
  XNOR2_X1 U480 ( .A(G122), .B(KEYINPUT77), .ZN(n541) );
  OR2_X1 U481 ( .A1(n616), .A2(n780), .ZN(n794) );
  INV_X1 U482 ( .A(KEYINPUT40), .ZN(n498) );
  NAND2_X1 U483 ( .A1(n427), .A2(n436), .ZN(n435) );
  AND2_X1 U484 ( .A1(n433), .A2(n365), .ZN(n360) );
  AND2_X1 U485 ( .A1(n434), .A2(n395), .ZN(n361) );
  XOR2_X1 U486 ( .A(KEYINPUT70), .B(KEYINPUT10), .Z(n362) );
  AND2_X1 U487 ( .A1(n698), .A2(n794), .ZN(n363) );
  AND2_X1 U488 ( .A1(n789), .A2(n454), .ZN(n364) );
  AND2_X1 U489 ( .A1(n361), .A2(n429), .ZN(n365) );
  INV_X1 U490 ( .A(G237), .ZN(n463) );
  AND2_X1 U491 ( .A1(n479), .A2(n482), .ZN(n366) );
  AND2_X1 U492 ( .A1(n496), .A2(n495), .ZN(n367) );
  XNOR2_X1 U493 ( .A(KEYINPUT75), .B(KEYINPUT34), .ZN(n368) );
  INV_X1 U494 ( .A(KEYINPUT106), .ZN(n457) );
  XOR2_X1 U495 ( .A(KEYINPUT65), .B(KEYINPUT45), .Z(n369) );
  OR2_X1 U496 ( .A1(n400), .A2(n468), .ZN(n370) );
  OR2_X1 U497 ( .A1(n738), .A2(n739), .ZN(n371) );
  AND2_X1 U498 ( .A1(n390), .A2(n476), .ZN(n372) );
  NAND2_X1 U499 ( .A1(n483), .A2(n477), .ZN(n373) );
  NAND2_X1 U500 ( .A1(n483), .A2(n477), .ZN(n468) );
  BUF_X1 U501 ( .A(n577), .Z(n374) );
  BUF_X1 U502 ( .A(n552), .Z(n375) );
  NAND2_X1 U503 ( .A1(n720), .A2(n558), .ZN(n483) );
  XNOR2_X1 U504 ( .A(n458), .B(KEYINPUT110), .ZN(n376) );
  XNOR2_X1 U505 ( .A(n458), .B(KEYINPUT110), .ZN(n416) );
  INV_X1 U506 ( .A(n730), .ZN(n485) );
  NAND2_X1 U507 ( .A1(n389), .A2(n388), .ZN(n387) );
  BUF_X1 U508 ( .A(n544), .Z(n377) );
  OR2_X2 U509 ( .A1(n376), .A2(KEYINPUT81), .ZN(n408) );
  BUF_X1 U510 ( .A(n768), .Z(n438) );
  NOR2_X1 U511 ( .A1(n768), .A2(n368), .ZN(n389) );
  BUF_X1 U512 ( .A(n736), .Z(n439) );
  XNOR2_X2 U513 ( .A(n803), .B(n551), .ZN(n470) );
  NAND2_X1 U514 ( .A1(n409), .A2(n408), .ZN(n378) );
  NAND2_X1 U515 ( .A1(n409), .A2(n408), .ZN(n599) );
  XNOR2_X1 U516 ( .A(n488), .B(n563), .ZN(n705) );
  XNOR2_X1 U517 ( .A(n490), .B(n489), .ZN(n488) );
  BUF_X1 U518 ( .A(n385), .Z(n710) );
  XNOR2_X1 U519 ( .A(n597), .B(n596), .ZN(n736) );
  XNOR2_X1 U520 ( .A(n689), .B(n545), .ZN(n379) );
  XNOR2_X1 U521 ( .A(n689), .B(n545), .ZN(n407) );
  NAND2_X1 U522 ( .A1(n399), .A2(n370), .ZN(n380) );
  XNOR2_X1 U523 ( .A(n603), .B(n602), .ZN(n629) );
  AND2_X1 U524 ( .A1(n759), .A2(n609), .ZN(n586) );
  XOR2_X1 U525 ( .A(n700), .B(KEYINPUT62), .Z(n701) );
  NAND2_X1 U526 ( .A1(n745), .A2(n609), .ZN(n393) );
  BUF_X1 U527 ( .A(n391), .Z(n381) );
  AND2_X2 U528 ( .A1(n486), .A2(n391), .ZN(n661) );
  BUF_X1 U529 ( .A(n686), .Z(n383) );
  INV_X1 U530 ( .A(n388), .ZN(n384) );
  NOR2_X1 U531 ( .A1(n729), .A2(n670), .ZN(n385) );
  BUF_X1 U532 ( .A(n652), .Z(n386) );
  XNOR2_X1 U533 ( .A(n652), .B(n405), .ZN(n649) );
  NOR2_X1 U534 ( .A1(n729), .A2(n670), .ZN(n719) );
  NAND2_X1 U535 ( .A1(n659), .A2(KEYINPUT44), .ZN(n658) );
  NAND2_X1 U536 ( .A1(n644), .A2(n686), .ZN(n659) );
  NAND2_X1 U537 ( .A1(n372), .A2(n387), .ZN(n475) );
  INV_X1 U538 ( .A(n649), .ZN(n388) );
  NAND2_X1 U539 ( .A1(n649), .A2(n368), .ZN(n390) );
  NAND2_X1 U540 ( .A1(n652), .A2(n633), .ZN(n635) );
  XNOR2_X2 U541 ( .A(n469), .B(KEYINPUT0), .ZN(n652) );
  NAND2_X1 U542 ( .A1(n663), .A2(n391), .ZN(n665) );
  AND2_X1 U543 ( .A1(n381), .A2(n485), .ZN(n731) );
  NAND2_X1 U544 ( .A1(n381), .A2(n795), .ZN(n799) );
  XNOR2_X2 U545 ( .A(n401), .B(n369), .ZN(n391) );
  NAND2_X2 U546 ( .A1(n417), .A2(n363), .ZN(n687) );
  XNOR2_X2 U547 ( .A(n528), .B(n527), .ZN(n458) );
  XNOR2_X1 U548 ( .A(n407), .B(n510), .ZN(n711) );
  NAND2_X1 U549 ( .A1(n431), .A2(KEYINPUT103), .ZN(n394) );
  NOR2_X1 U550 ( .A1(n699), .A2(n656), .ZN(n657) );
  NAND2_X1 U551 ( .A1(n430), .A2(n428), .ZN(n699) );
  NAND2_X1 U552 ( .A1(n658), .A2(n657), .ZN(n404) );
  XNOR2_X1 U553 ( .A(n420), .B(n595), .ZN(n419) );
  NAND2_X1 U554 ( .A1(n419), .A2(n447), .ZN(n418) );
  NAND2_X1 U555 ( .A1(n456), .A2(n457), .ZN(n455) );
  INV_X1 U556 ( .A(n396), .ZN(n610) );
  NAND2_X1 U557 ( .A1(n397), .A2(n402), .ZN(n401) );
  XNOR2_X1 U558 ( .A(n404), .B(n424), .ZN(n397) );
  NAND2_X1 U559 ( .A1(n373), .A2(n484), .ZN(n398) );
  NAND2_X1 U560 ( .A1(n479), .A2(KEYINPUT92), .ZN(n400) );
  NAND2_X1 U561 ( .A1(n367), .A2(n406), .ZN(n616) );
  XNOR2_X1 U562 ( .A(n379), .B(n538), .ZN(n700) );
  AND2_X2 U563 ( .A1(n414), .A2(n410), .ZN(n409) );
  NAND2_X1 U564 ( .A1(n416), .A2(n415), .ZN(n414) );
  AND2_X1 U565 ( .A1(n587), .A2(KEYINPUT81), .ZN(n415) );
  NAND2_X1 U566 ( .A1(n417), .A2(n698), .ZN(n621) );
  NAND2_X1 U567 ( .A1(n500), .A2(n380), .ZN(n420) );
  NOR2_X1 U568 ( .A1(n645), .A2(n455), .ZN(n423) );
  XNOR2_X2 U569 ( .A(n745), .B(KEYINPUT6), .ZN(n645) );
  XNOR2_X2 U570 ( .A(n552), .B(n440), .ZN(n689) );
  OR2_X2 U571 ( .A1(n720), .A2(n480), .ZN(n479) );
  XNOR2_X2 U572 ( .A(n470), .B(n554), .ZN(n720) );
  NAND2_X1 U573 ( .A1(n435), .A2(n360), .ZN(n428) );
  NAND2_X1 U574 ( .A1(n433), .A2(n361), .ZN(n431) );
  NAND2_X1 U575 ( .A1(n643), .A2(n647), .ZN(n433) );
  NAND2_X1 U576 ( .A1(n646), .A2(n647), .ZN(n434) );
  XNOR2_X1 U577 ( .A(n665), .B(n664), .ZN(n669) );
  NOR2_X2 U578 ( .A1(n629), .A2(n628), .ZN(n469) );
  NAND2_X1 U579 ( .A1(n475), .A2(n631), .ZN(n437) );
  NOR2_X1 U580 ( .A1(n643), .A2(n638), .ZN(n640) );
  XNOR2_X2 U581 ( .A(n635), .B(n634), .ZN(n643) );
  XNOR2_X1 U582 ( .A(n445), .B(KEYINPUT46), .ZN(n443) );
  XNOR2_X2 U583 ( .A(n577), .B(n442), .ZN(n552) );
  XNOR2_X2 U584 ( .A(n505), .B(KEYINPUT69), .ZN(n442) );
  XNOR2_X2 U585 ( .A(n471), .B(G143), .ZN(n577) );
  INV_X1 U586 ( .A(n736), .ZN(n447) );
  NAND2_X1 U587 ( .A1(n736), .A2(KEYINPUT105), .ZN(n449) );
  OR2_X1 U588 ( .A1(n439), .A2(n371), .ZN(n650) );
  NAND2_X1 U589 ( .A1(n453), .A2(n472), .ZN(n452) );
  INV_X1 U590 ( .A(n592), .ZN(n456) );
  NAND2_X1 U591 ( .A1(n651), .A2(n458), .ZN(n648) );
  NAND2_X1 U592 ( .A1(n582), .A2(n705), .ZN(n461) );
  XNOR2_X2 U593 ( .A(G128), .B(KEYINPUT85), .ZN(n471) );
  INV_X1 U594 ( .A(n645), .ZN(n472) );
  XNOR2_X2 U595 ( .A(KEYINPUT4), .B(G146), .ZN(n505) );
  XNOR2_X2 U596 ( .A(n474), .B(n473), .ZN(n544) );
  XNOR2_X2 U597 ( .A(n536), .B(KEYINPUT3), .ZN(n474) );
  NAND2_X1 U598 ( .A1(n768), .A2(n368), .ZN(n476) );
  NAND2_X1 U599 ( .A1(n366), .A2(n483), .ZN(n593) );
  INV_X1 U600 ( .A(n482), .ZN(n478) );
  NAND2_X1 U601 ( .A1(n558), .A2(n666), .ZN(n482) );
  INV_X1 U602 ( .A(KEYINPUT92), .ZN(n484) );
  INV_X1 U603 ( .A(n660), .ZN(n486) );
  XNOR2_X1 U604 ( .A(n518), .B(n517), .ZN(n489) );
  NAND2_X1 U605 ( .A1(n579), .A2(G221), .ZN(n490) );
  INV_X2 U606 ( .A(KEYINPUT64), .ZN(n491) );
  XNOR2_X2 U607 ( .A(n491), .B(G953), .ZN(n690) );
  INV_X1 U608 ( .A(n495), .ZN(n493) );
  NOR2_X1 U609 ( .A1(n752), .A2(n497), .ZN(n494) );
  NAND2_X1 U610 ( .A1(n752), .A2(n497), .ZN(n495) );
  NAND2_X1 U611 ( .A1(n599), .A2(n497), .ZN(n496) );
  INV_X1 U612 ( .A(KEYINPUT39), .ZN(n497) );
  INV_X1 U613 ( .A(KEYINPUT48), .ZN(n499) );
  XNOR2_X2 U614 ( .A(n661), .B(KEYINPUT80), .ZN(n729) );
  NOR2_X2 U615 ( .A1(n597), .A2(n735), .ZN(n528) );
  XNOR2_X1 U616 ( .A(KEYINPUT96), .B(KEYINPUT25), .ZN(n502) );
  XOR2_X1 U617 ( .A(n562), .B(n561), .Z(n503) );
  XNOR2_X1 U618 ( .A(n516), .B(n515), .ZN(n517) );
  INV_X1 U619 ( .A(KEYINPUT88), .ZN(n664) );
  XNOR2_X1 U620 ( .A(n563), .B(n503), .ZN(n570) );
  XNOR2_X1 U621 ( .A(n594), .B(KEYINPUT91), .ZN(n595) );
  BUF_X1 U622 ( .A(n687), .Z(n730) );
  BUF_X1 U623 ( .A(n711), .Z(n714) );
  INV_X1 U624 ( .A(n679), .ZN(n680) );
  XNOR2_X1 U625 ( .A(n681), .B(n680), .ZN(n682) );
  XNOR2_X1 U626 ( .A(n507), .B(n506), .ZN(n801) );
  XNOR2_X1 U627 ( .A(n801), .B(KEYINPUT74), .ZN(n553) );
  NAND2_X1 U628 ( .A1(n690), .A2(G227), .ZN(n508) );
  XNOR2_X1 U629 ( .A(n508), .B(G140), .ZN(n509) );
  XNOR2_X1 U630 ( .A(n553), .B(n509), .ZN(n510) );
  OR2_X2 U631 ( .A1(n711), .A2(G902), .ZN(n512) );
  XOR2_X1 U632 ( .A(KEYINPUT72), .B(G469), .Z(n511) );
  XNOR2_X2 U633 ( .A(n512), .B(n511), .ZN(n597) );
  XOR2_X1 U634 ( .A(KEYINPUT23), .B(KEYINPUT95), .Z(n514) );
  XNOR2_X1 U635 ( .A(G119), .B(G137), .ZN(n513) );
  XNOR2_X1 U636 ( .A(n514), .B(n513), .ZN(n518) );
  XNOR2_X1 U637 ( .A(G128), .B(G110), .ZN(n516) );
  INV_X1 U638 ( .A(KEYINPUT24), .ZN(n515) );
  NAND2_X1 U639 ( .A1(n690), .A2(G234), .ZN(n520) );
  XNOR2_X1 U640 ( .A(n520), .B(n519), .ZN(n579) );
  XNOR2_X1 U641 ( .A(G125), .B(G140), .ZN(n521) );
  NAND2_X1 U642 ( .A1(n662), .A2(G234), .ZN(n522) );
  XNOR2_X1 U643 ( .A(n522), .B(KEYINPUT20), .ZN(n525) );
  NAND2_X1 U644 ( .A1(G217), .A2(n525), .ZN(n523) );
  XNOR2_X1 U645 ( .A(n523), .B(n502), .ZN(n524) );
  NAND2_X1 U646 ( .A1(n525), .A2(G221), .ZN(n526) );
  XNOR2_X1 U647 ( .A(n526), .B(KEYINPUT21), .ZN(n739) );
  XNOR2_X1 U648 ( .A(KEYINPUT14), .B(n529), .ZN(n734) );
  INV_X1 U649 ( .A(n690), .ZN(n675) );
  NOR2_X1 U650 ( .A1(n582), .A2(G900), .ZN(n530) );
  NAND2_X1 U651 ( .A1(n675), .A2(n530), .ZN(n531) );
  NAND2_X1 U652 ( .A1(G952), .A2(n795), .ZN(n625) );
  NAND2_X1 U653 ( .A1(n531), .A2(n625), .ZN(n532) );
  NAND2_X1 U654 ( .A1(n734), .A2(n532), .ZN(n533) );
  XOR2_X1 U655 ( .A(KEYINPUT86), .B(n533), .Z(n587) );
  NAND2_X1 U656 ( .A1(n564), .A2(G210), .ZN(n535) );
  XOR2_X1 U657 ( .A(KEYINPUT98), .B(KEYINPUT5), .Z(n534) );
  XNOR2_X1 U658 ( .A(n535), .B(n534), .ZN(n537) );
  XNOR2_X2 U659 ( .A(G113), .B(KEYINPUT73), .ZN(n536) );
  XNOR2_X1 U660 ( .A(n377), .B(n537), .ZN(n538) );
  XNOR2_X2 U661 ( .A(n539), .B(G472), .ZN(n745) );
  NAND2_X1 U662 ( .A1(n582), .A2(n463), .ZN(n555) );
  NAND2_X1 U663 ( .A1(n555), .A2(G214), .ZN(n609) );
  XNOR2_X1 U664 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X2 U665 ( .A(n544), .B(n543), .ZN(n803) );
  NAND2_X1 U666 ( .A1(n690), .A2(G224), .ZN(n546) );
  XNOR2_X1 U667 ( .A(n546), .B(n545), .ZN(n550) );
  XNOR2_X1 U668 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U669 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U670 ( .A(n375), .B(n553), .ZN(n554) );
  INV_X1 U671 ( .A(n662), .ZN(n666) );
  NAND2_X1 U672 ( .A1(n555), .A2(G210), .ZN(n557) );
  INV_X1 U673 ( .A(KEYINPUT93), .ZN(n556) );
  XNOR2_X1 U674 ( .A(n557), .B(n556), .ZN(n558) );
  INV_X1 U675 ( .A(KEYINPUT38), .ZN(n559) );
  XNOR2_X1 U676 ( .A(n560), .B(KEYINPUT100), .ZN(n561) );
  NAND2_X1 U677 ( .A1(G214), .A2(n564), .ZN(n566) );
  XNOR2_X1 U678 ( .A(n566), .B(n565), .ZN(n568) );
  XNOR2_X1 U679 ( .A(n568), .B(n567), .ZN(n569) );
  INV_X1 U680 ( .A(KEYINPUT13), .ZN(n571) );
  XNOR2_X1 U681 ( .A(n572), .B(KEYINPUT7), .ZN(n576) );
  XOR2_X1 U682 ( .A(KEYINPUT9), .B(KEYINPUT101), .Z(n574) );
  XNOR2_X1 U683 ( .A(n574), .B(n573), .ZN(n575) );
  XOR2_X1 U684 ( .A(n576), .B(n575), .Z(n578) );
  XNOR2_X1 U685 ( .A(n374), .B(n578), .ZN(n581) );
  AND2_X1 U686 ( .A1(n579), .A2(G217), .ZN(n580) );
  XNOR2_X1 U687 ( .A(n581), .B(n580), .ZN(n679) );
  NAND2_X1 U688 ( .A1(n679), .A2(n582), .ZN(n583) );
  XNOR2_X1 U689 ( .A(n583), .B(G478), .ZN(n598) );
  INV_X1 U690 ( .A(n598), .ZN(n605) );
  NAND2_X1 U691 ( .A1(n606), .A2(n605), .ZN(n786) );
  NOR2_X1 U692 ( .A1(n606), .A2(n598), .ZN(n585) );
  INV_X1 U693 ( .A(KEYINPUT102), .ZN(n584) );
  XNOR2_X1 U694 ( .A(n585), .B(n584), .ZN(n751) );
  NOR2_X1 U695 ( .A1(n751), .A2(n752), .ZN(n759) );
  INV_X1 U696 ( .A(n745), .ZN(n651) );
  NAND2_X1 U697 ( .A1(n588), .A2(n587), .ZN(n592) );
  NOR2_X1 U698 ( .A1(n767), .A2(n604), .ZN(n591) );
  XNOR2_X1 U699 ( .A(KEYINPUT112), .B(KEYINPUT42), .ZN(n590) );
  INV_X1 U700 ( .A(n609), .ZN(n757) );
  XNOR2_X1 U701 ( .A(KEYINPUT114), .B(KEYINPUT36), .ZN(n594) );
  XNOR2_X1 U702 ( .A(KEYINPUT66), .B(KEYINPUT1), .ZN(n596) );
  NAND2_X1 U703 ( .A1(n606), .A2(n598), .ZN(n630) );
  NOR2_X1 U704 ( .A1(n378), .A2(n593), .ZN(n600) );
  XNOR2_X1 U705 ( .A(n600), .B(KEYINPUT111), .ZN(n601) );
  NOR2_X1 U706 ( .A1(n630), .A2(n601), .ZN(n785) );
  XNOR2_X1 U707 ( .A(KEYINPUT82), .B(KEYINPUT19), .ZN(n602) );
  OR2_X1 U708 ( .A1(n604), .A2(n629), .ZN(n787) );
  NOR2_X1 U709 ( .A1(n606), .A2(n605), .ZN(n791) );
  NOR2_X1 U710 ( .A1(n791), .A2(n789), .ZN(n753) );
  XNOR2_X1 U711 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n608) );
  XNOR2_X1 U712 ( .A(n608), .B(KEYINPUT43), .ZN(n614) );
  NAND2_X1 U713 ( .A1(n610), .A2(n609), .ZN(n611) );
  XOR2_X1 U714 ( .A(KEYINPUT107), .B(n611), .Z(n612) );
  NOR2_X1 U715 ( .A1(n447), .A2(n612), .ZN(n613) );
  XNOR2_X1 U716 ( .A(n614), .B(n613), .ZN(n615) );
  NAND2_X1 U717 ( .A1(n615), .A2(n593), .ZN(n698) );
  INV_X1 U718 ( .A(n791), .ZN(n780) );
  INV_X1 U719 ( .A(KEYINPUT87), .ZN(n617) );
  NAND2_X1 U720 ( .A1(n617), .A2(KEYINPUT2), .ZN(n618) );
  NOR2_X1 U721 ( .A1(n687), .A2(n618), .ZN(n623) );
  NAND2_X1 U722 ( .A1(n794), .A2(KEYINPUT2), .ZN(n619) );
  NAND2_X1 U723 ( .A1(n619), .A2(KEYINPUT87), .ZN(n620) );
  NOR2_X1 U724 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U725 ( .A1(n623), .A2(n622), .ZN(n660) );
  INV_X1 U726 ( .A(KEYINPUT33), .ZN(n624) );
  NOR2_X1 U727 ( .A1(G898), .A2(n795), .ZN(n805) );
  NAND2_X1 U728 ( .A1(n805), .A2(G902), .ZN(n626) );
  NAND2_X1 U729 ( .A1(n626), .A2(n625), .ZN(n627) );
  NAND2_X1 U730 ( .A1(n627), .A2(n734), .ZN(n628) );
  INV_X1 U731 ( .A(n630), .ZN(n631) );
  INV_X1 U732 ( .A(KEYINPUT35), .ZN(n632) );
  NOR2_X1 U733 ( .A1(n751), .A2(n739), .ZN(n633) );
  NOR2_X1 U734 ( .A1(n439), .A2(n395), .ZN(n636) );
  XNOR2_X1 U735 ( .A(n636), .B(KEYINPUT104), .ZN(n637) );
  NAND2_X1 U736 ( .A1(n637), .A2(n645), .ZN(n638) );
  XNOR2_X1 U737 ( .A(KEYINPUT84), .B(KEYINPUT32), .ZN(n639) );
  XNOR2_X1 U738 ( .A(n640), .B(n639), .ZN(n685) );
  NOR2_X1 U739 ( .A1(n745), .A2(n395), .ZN(n641) );
  NAND2_X1 U740 ( .A1(n439), .A2(n641), .ZN(n642) );
  NOR2_X1 U741 ( .A1(n382), .A2(n642), .ZN(n683) );
  NOR2_X1 U742 ( .A1(n685), .A2(n683), .ZN(n644) );
  NAND2_X1 U743 ( .A1(n645), .A2(n439), .ZN(n646) );
  NOR2_X1 U744 ( .A1(n384), .A2(n648), .ZN(n776) );
  NOR2_X1 U745 ( .A1(n651), .A2(n650), .ZN(n747) );
  NAND2_X1 U746 ( .A1(n386), .A2(n747), .ZN(n654) );
  XOR2_X1 U747 ( .A(KEYINPUT99), .B(KEYINPUT31), .Z(n653) );
  XNOR2_X1 U748 ( .A(n654), .B(n653), .ZN(n792) );
  NOR2_X1 U749 ( .A1(n776), .A2(n792), .ZN(n655) );
  NOR2_X1 U750 ( .A1(n655), .A2(n753), .ZN(n656) );
  NOR2_X1 U751 ( .A1(n687), .A2(n662), .ZN(n663) );
  NAND2_X1 U752 ( .A1(n666), .A2(KEYINPUT2), .ZN(n667) );
  NOR2_X1 U753 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U754 ( .A1(n719), .A2(G475), .ZN(n673) );
  XNOR2_X1 U755 ( .A(n673), .B(n672), .ZN(n676) );
  INV_X1 U756 ( .A(G952), .ZN(n674) );
  NAND2_X1 U757 ( .A1(n675), .A2(n674), .ZN(n725) );
  NAND2_X1 U758 ( .A1(n676), .A2(n725), .ZN(n678) );
  INV_X1 U759 ( .A(KEYINPUT60), .ZN(n677) );
  XNOR2_X1 U760 ( .A(n678), .B(n677), .ZN(G60) );
  NAND2_X1 U761 ( .A1(n710), .A2(G478), .ZN(n681) );
  INV_X1 U762 ( .A(n725), .ZN(n717) );
  NOR2_X1 U763 ( .A1(n682), .A2(n717), .ZN(G63) );
  XOR2_X1 U764 ( .A(G110), .B(n683), .Z(G12) );
  NAND2_X1 U765 ( .A1(n776), .A2(n789), .ZN(n684) );
  XNOR2_X1 U766 ( .A(n684), .B(G104), .ZN(G6) );
  XOR2_X1 U767 ( .A(n685), .B(G119), .Z(G21) );
  XNOR2_X1 U768 ( .A(n383), .B(G122), .ZN(G24) );
  XNOR2_X1 U769 ( .A(n689), .B(n688), .ZN(n692) );
  XNOR2_X1 U770 ( .A(n730), .B(n692), .ZN(n691) );
  NAND2_X1 U771 ( .A1(n691), .A2(n690), .ZN(n697) );
  XNOR2_X1 U772 ( .A(G227), .B(n692), .ZN(n693) );
  NAND2_X1 U773 ( .A1(n693), .A2(G900), .ZN(n694) );
  XOR2_X1 U774 ( .A(KEYINPUT127), .B(n694), .Z(n695) );
  NAND2_X1 U775 ( .A1(n695), .A2(G953), .ZN(n696) );
  NAND2_X1 U776 ( .A1(n697), .A2(n696), .ZN(G72) );
  XNOR2_X1 U777 ( .A(n698), .B(G140), .ZN(G42) );
  XOR2_X1 U778 ( .A(n699), .B(G101), .Z(G3) );
  NAND2_X1 U779 ( .A1(n385), .A2(G472), .ZN(n702) );
  XNOR2_X1 U780 ( .A(n702), .B(n701), .ZN(n703) );
  NAND2_X1 U781 ( .A1(n703), .A2(n725), .ZN(n704) );
  XNOR2_X1 U782 ( .A(n704), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U783 ( .A1(n710), .A2(G217), .ZN(n708) );
  XNOR2_X1 U784 ( .A(KEYINPUT124), .B(KEYINPUT125), .ZN(n706) );
  XNOR2_X1 U785 ( .A(n705), .B(n706), .ZN(n707) );
  XNOR2_X1 U786 ( .A(n708), .B(n707), .ZN(n709) );
  NOR2_X1 U787 ( .A1(n709), .A2(n717), .ZN(G66) );
  NAND2_X1 U788 ( .A1(n710), .A2(G469), .ZN(n716) );
  XNOR2_X1 U789 ( .A(KEYINPUT123), .B(KEYINPUT57), .ZN(n712) );
  XNOR2_X1 U790 ( .A(n712), .B(KEYINPUT58), .ZN(n713) );
  XNOR2_X1 U791 ( .A(n714), .B(n713), .ZN(n715) );
  XNOR2_X1 U792 ( .A(n716), .B(n715), .ZN(n718) );
  NOR2_X1 U793 ( .A1(n718), .A2(n717), .ZN(G54) );
  NAND2_X1 U794 ( .A1(n719), .A2(G210), .ZN(n724) );
  XNOR2_X1 U795 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n721) );
  XNOR2_X1 U796 ( .A(n724), .B(n723), .ZN(n726) );
  NAND2_X1 U797 ( .A1(n726), .A2(n725), .ZN(n728) );
  XOR2_X1 U798 ( .A(KEYINPUT122), .B(KEYINPUT56), .Z(n727) );
  XNOR2_X1 U799 ( .A(n728), .B(n727), .ZN(G51) );
  BUF_X1 U800 ( .A(n729), .Z(n733) );
  NOR2_X1 U801 ( .A1(n731), .A2(KEYINPUT2), .ZN(n732) );
  NOR2_X1 U802 ( .A1(n733), .A2(n732), .ZN(n773) );
  NAND2_X1 U803 ( .A1(G952), .A2(n734), .ZN(n765) );
  NAND2_X1 U804 ( .A1(n439), .A2(n371), .ZN(n737) );
  XNOR2_X1 U805 ( .A(KEYINPUT50), .B(n737), .ZN(n743) );
  XOR2_X1 U806 ( .A(KEYINPUT118), .B(KEYINPUT49), .Z(n741) );
  NAND2_X1 U807 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U808 ( .A(n741), .B(n740), .ZN(n742) );
  NAND2_X1 U809 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U810 ( .A1(n745), .A2(n744), .ZN(n746) );
  NOR2_X1 U811 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U812 ( .A(n748), .B(KEYINPUT119), .ZN(n749) );
  XNOR2_X1 U813 ( .A(KEYINPUT51), .B(n749), .ZN(n750) );
  NOR2_X1 U814 ( .A1(n767), .A2(n750), .ZN(n762) );
  INV_X1 U815 ( .A(n751), .ZN(n755) );
  NOR2_X1 U816 ( .A1(n753), .A2(n752), .ZN(n754) );
  NOR2_X1 U817 ( .A1(n755), .A2(n754), .ZN(n756) );
  NOR2_X1 U818 ( .A1(n757), .A2(n756), .ZN(n758) );
  NOR2_X1 U819 ( .A1(n759), .A2(n758), .ZN(n760) );
  NOR2_X1 U820 ( .A1(n438), .A2(n760), .ZN(n761) );
  NOR2_X1 U821 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U822 ( .A(n763), .B(KEYINPUT52), .ZN(n764) );
  NOR2_X1 U823 ( .A1(n765), .A2(n764), .ZN(n766) );
  XOR2_X1 U824 ( .A(KEYINPUT120), .B(n766), .Z(n771) );
  NOR2_X1 U825 ( .A1(n438), .A2(n767), .ZN(n769) );
  NOR2_X1 U826 ( .A1(n769), .A2(G953), .ZN(n770) );
  NAND2_X1 U827 ( .A1(n771), .A2(n770), .ZN(n772) );
  NOR2_X1 U828 ( .A1(n773), .A2(n772), .ZN(n775) );
  XOR2_X1 U829 ( .A(KEYINPUT121), .B(KEYINPUT53), .Z(n774) );
  XNOR2_X1 U830 ( .A(n775), .B(n774), .ZN(G75) );
  NAND2_X1 U831 ( .A1(n776), .A2(n791), .ZN(n778) );
  XOR2_X1 U832 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n777) );
  XNOR2_X1 U833 ( .A(n778), .B(n777), .ZN(n779) );
  XNOR2_X1 U834 ( .A(G107), .B(n779), .ZN(G9) );
  NOR2_X1 U835 ( .A1(n787), .A2(n780), .ZN(n784) );
  XOR2_X1 U836 ( .A(KEYINPUT116), .B(KEYINPUT29), .Z(n782) );
  XNOR2_X1 U837 ( .A(G128), .B(KEYINPUT117), .ZN(n781) );
  XNOR2_X1 U838 ( .A(n782), .B(n781), .ZN(n783) );
  XNOR2_X1 U839 ( .A(n784), .B(n783), .ZN(G30) );
  XOR2_X1 U840 ( .A(G143), .B(n785), .Z(G45) );
  NOR2_X1 U841 ( .A1(n787), .A2(n786), .ZN(n788) );
  XOR2_X1 U842 ( .A(n355), .B(n788), .Z(G48) );
  NAND2_X1 U843 ( .A1(n792), .A2(n789), .ZN(n790) );
  XNOR2_X1 U844 ( .A(n790), .B(G113), .ZN(G15) );
  NAND2_X1 U845 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U846 ( .A(n793), .B(G116), .ZN(G18) );
  XNOR2_X1 U847 ( .A(G134), .B(n794), .ZN(G36) );
  NAND2_X1 U848 ( .A1(G953), .A2(G224), .ZN(n796) );
  XNOR2_X1 U849 ( .A(KEYINPUT61), .B(n796), .ZN(n797) );
  NAND2_X1 U850 ( .A1(n797), .A2(G898), .ZN(n798) );
  NAND2_X1 U851 ( .A1(n799), .A2(n798), .ZN(n807) );
  XOR2_X1 U852 ( .A(G101), .B(KEYINPUT126), .Z(n800) );
  XNOR2_X1 U853 ( .A(n801), .B(n800), .ZN(n802) );
  XNOR2_X1 U854 ( .A(n803), .B(n802), .ZN(n804) );
  NOR2_X1 U855 ( .A1(n805), .A2(n804), .ZN(n806) );
  XNOR2_X1 U856 ( .A(n807), .B(n806), .ZN(G69) );
  XNOR2_X1 U857 ( .A(n808), .B(G125), .ZN(n809) );
  XNOR2_X1 U858 ( .A(n809), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U859 ( .A(n810), .B(G137), .Z(G39) );
  BUF_X1 U860 ( .A(n811), .Z(n812) );
  XOR2_X1 U861 ( .A(G131), .B(n812), .Z(G33) );
endmodule

