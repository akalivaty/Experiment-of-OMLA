//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 1 1 1 1 1 1 1 1 1 0 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1 0 1 0 0 0 0 0 1 0 1 0 1 1 1 1 1 1 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:33 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n604,
    new_n606, new_n607, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT65), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n451), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n451), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT66), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n460), .A2(G2105), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT70), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT67), .B(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(new_n463), .A2(G137), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(new_n460), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI22_X1  g043(.A1(G101), .A2(new_n462), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n470));
  AND2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  OAI21_X1  g047(.A(KEYINPUT68), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n466), .A2(new_n474), .A3(new_n467), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n473), .A2(new_n475), .A3(G125), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n463), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n470), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AOI211_X1 g055(.A(KEYINPUT69), .B(new_n463), .C1(new_n476), .C2(new_n477), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n469), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G160));
  OAI221_X1 g058(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n463), .C2(G112), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n484), .B(KEYINPUT71), .ZN(new_n485));
  INV_X1    g060(.A(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n468), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n489));
  AOI22_X1  g064(.A1(new_n488), .A2(G136), .B1(new_n489), .B2(G124), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n485), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n491), .B(KEYINPUT72), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  NAND3_X1  g068(.A1(new_n468), .A2(G126), .A3(G2105), .ZN(new_n494));
  OR2_X1    g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n495), .B(G2104), .C1(G114), .C2(new_n486), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n486), .A2(KEYINPUT67), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT67), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G2105), .ZN(new_n500));
  AND3_X1   g075(.A1(new_n498), .A2(new_n500), .A3(G138), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n501), .A2(new_n502), .A3(new_n473), .A4(new_n475), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT73), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n468), .A2(new_n463), .A3(G138), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n503), .A2(new_n504), .B1(KEYINPUT4), .B2(new_n505), .ZN(new_n506));
  AND4_X1   g081(.A1(new_n502), .A2(new_n498), .A3(new_n500), .A4(G138), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n507), .A2(KEYINPUT73), .A3(new_n473), .A4(new_n475), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n497), .B1(new_n506), .B2(new_n508), .ZN(G164));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT75), .A2(G543), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g088(.A1(KEYINPUT75), .A2(KEYINPUT5), .A3(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g090(.A(KEYINPUT76), .B1(new_n515), .B2(G62), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n516), .B1(G75), .B2(G543), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n515), .A2(KEYINPUT76), .A3(G62), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n510), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT6), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT74), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n520), .B1(new_n521), .B2(new_n510), .ZN(new_n522));
  NAND3_X1  g097(.A1(KEYINPUT74), .A2(KEYINPUT6), .A3(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n524), .A2(G50), .A3(G543), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n515), .ZN(new_n526));
  INV_X1    g101(.A(G88), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n519), .A2(new_n528), .ZN(G166));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  INV_X1    g106(.A(G89), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n531), .B1(new_n526), .B2(new_n532), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT78), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT77), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n524), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n522), .A2(KEYINPUT77), .A3(new_n523), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n536), .A2(G543), .A3(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  AND2_X1   g114(.A1(G63), .A2(G651), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n539), .A2(G51), .B1(new_n515), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n534), .A2(new_n541), .ZN(G286));
  INV_X1    g117(.A(G286), .ZN(G168));
  NAND2_X1  g118(.A1(new_n539), .A2(G52), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(new_n510), .ZN(new_n546));
  INV_X1    g121(.A(new_n526), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G90), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n544), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(G171));
  NAND2_X1  g125(.A1(new_n539), .A2(G43), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n515), .A2(G56), .ZN(new_n552));
  NAND2_X1  g127(.A1(G68), .A2(G543), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n510), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n554), .B1(G81), .B2(new_n547), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  AOI22_X1  g137(.A1(new_n515), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n563));
  OR3_X1    g138(.A1(new_n563), .A2(KEYINPUT79), .A3(new_n510), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT79), .B1(new_n563), .B2(new_n510), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n564), .A2(new_n565), .B1(G91), .B2(new_n547), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n536), .A2(G53), .A3(G543), .A4(new_n537), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT9), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n566), .A2(new_n568), .ZN(G299));
  XOR2_X1   g144(.A(new_n549), .B(KEYINPUT80), .Z(G301));
  INV_X1    g145(.A(G166), .ZN(G303));
  NAND2_X1  g146(.A1(new_n539), .A2(G49), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n547), .A2(G87), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(G288));
  NAND2_X1  g150(.A1(G73), .A2(G543), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT81), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n515), .A2(G61), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n510), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n524), .A2(G86), .A3(new_n515), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n524), .A2(G48), .A3(G543), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(G305));
  NAND2_X1  g160(.A1(new_n547), .A2(G85), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G47), .ZN(new_n588));
  OAI221_X1 g163(.A(new_n586), .B1(new_n510), .B2(new_n587), .C1(new_n588), .C2(new_n538), .ZN(G290));
  INV_X1    g164(.A(G868), .ZN(new_n590));
  NOR2_X1   g165(.A1(G301), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(G54), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n515), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n593));
  OAI22_X1  g168(.A1(new_n538), .A2(new_n592), .B1(new_n510), .B2(new_n593), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT82), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n547), .A2(G92), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n596), .B(KEYINPUT10), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n591), .B1(new_n590), .B2(new_n598), .ZN(G284));
  AOI21_X1  g174(.A(new_n591), .B1(new_n590), .B2(new_n598), .ZN(G321));
  NAND2_X1  g175(.A1(G299), .A2(new_n590), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(G168), .B2(new_n590), .ZN(G297));
  OAI21_X1  g177(.A(new_n601), .B1(G168), .B2(new_n590), .ZN(G280));
  INV_X1    g178(.A(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n598), .B1(new_n604), .B2(G860), .ZN(G148));
  NAND2_X1  g180(.A1(new_n598), .A2(new_n604), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(G868), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(G868), .B2(new_n557), .ZN(G323));
  XNOR2_X1  g183(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g184(.A1(new_n462), .A2(new_n473), .A3(new_n475), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT12), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT13), .ZN(new_n612));
  INV_X1    g187(.A(G2100), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(KEYINPUT83), .Z(new_n615));
  NAND2_X1  g190(.A1(new_n489), .A2(G123), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT84), .ZN(new_n617));
  OR2_X1    g192(.A1(new_n463), .A2(G111), .ZN(new_n618));
  OAI21_X1  g193(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n619));
  INV_X1    g194(.A(new_n619), .ZN(new_n620));
  AOI22_X1  g195(.A1(G135), .A2(new_n488), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2096), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n623), .B1(new_n612), .B2(new_n613), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n615), .A2(new_n624), .ZN(G156));
  INV_X1    g200(.A(KEYINPUT14), .ZN(new_n626));
  XNOR2_X1  g201(.A(G2427), .B(G2438), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2430), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT15), .B(G2435), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n626), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(new_n629), .B2(new_n628), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2451), .B(G2454), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT16), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT85), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n631), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2443), .B(G2446), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT86), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n635), .B(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G1341), .B(G1348), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  AND3_X1   g217(.A1(new_n641), .A2(new_n642), .A3(G14), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT87), .ZN(G401));
  INV_X1    g219(.A(KEYINPUT18), .ZN(new_n645));
  XOR2_X1   g220(.A(G2084), .B(G2090), .Z(new_n646));
  XNOR2_X1  g221(.A(G2067), .B(G2678), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(KEYINPUT17), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n646), .A2(new_n647), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n645), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(new_n613), .ZN(new_n652));
  XOR2_X1   g227(.A(G2072), .B(G2078), .Z(new_n653));
  AOI21_X1  g228(.A(new_n653), .B1(new_n648), .B2(KEYINPUT18), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(G2096), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n652), .B(new_n655), .ZN(G227));
  XNOR2_X1  g231(.A(G1961), .B(G1966), .ZN(new_n657));
  INV_X1    g232(.A(KEYINPUT89), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G1956), .B(G2474), .Z(new_n660));
  OR2_X1    g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1971), .B(G1976), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n661), .A2(new_n662), .A3(new_n665), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n662), .A2(new_n665), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT91), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT90), .B(KEYINPUT20), .ZN(new_n669));
  AND2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n668), .A2(new_n669), .ZN(new_n671));
  OAI221_X1 g246(.A(new_n666), .B1(new_n665), .B2(new_n661), .C1(new_n670), .C2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G1991), .B(G1996), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1981), .B(G1986), .ZN(new_n677));
  AND2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n676), .A2(new_n677), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(G229));
  INV_X1    g255(.A(G16), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(G20), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT23), .Z(new_n683));
  AOI21_X1  g258(.A(new_n683), .B1(G299), .B2(G16), .ZN(new_n684));
  INV_X1    g259(.A(G1956), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(G29), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(G35), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n688), .B(KEYINPUT99), .Z(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(G162), .B2(new_n687), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT29), .Z(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n686), .B1(new_n692), .B2(G2090), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT100), .Z(new_n694));
  NOR2_X1   g269(.A1(G6), .A2(G16), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(new_n584), .B2(G16), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT92), .Z(new_n697));
  XOR2_X1   g272(.A(KEYINPUT32), .B(G1981), .Z(new_n698));
  NAND2_X1  g273(.A1(G166), .A2(G16), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G16), .B2(G22), .ZN(new_n700));
  INV_X1    g275(.A(G1971), .ZN(new_n701));
  AOI22_X1  g276(.A1(new_n697), .A2(new_n698), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(new_n701), .B2(new_n700), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n681), .A2(G23), .ZN(new_n704));
  AND3_X1   g279(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n704), .B1(new_n705), .B2(new_n681), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT33), .B(G1976), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(new_n698), .B2(new_n697), .ZN(new_n709));
  OR3_X1    g284(.A1(new_n703), .A2(new_n709), .A3(KEYINPUT34), .ZN(new_n710));
  OAI21_X1  g285(.A(KEYINPUT34), .B1(new_n703), .B2(new_n709), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n681), .A2(G24), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(G290), .B2(G16), .ZN(new_n713));
  INV_X1    g288(.A(G1986), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n687), .A2(G25), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n488), .A2(G131), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n489), .A2(G119), .ZN(new_n718));
  OAI221_X1 g293(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n463), .C2(G107), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n716), .B1(new_n721), .B2(new_n687), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT35), .B(G1991), .Z(new_n723));
  XOR2_X1   g298(.A(new_n722), .B(new_n723), .Z(new_n724));
  INV_X1    g299(.A(new_n713), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n724), .B1(G1986), .B2(new_n725), .ZN(new_n726));
  NAND4_X1  g301(.A1(new_n710), .A2(new_n711), .A3(new_n715), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT36), .ZN(new_n728));
  INV_X1    g303(.A(G2090), .ZN(new_n729));
  INV_X1    g304(.A(G1348), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n598), .A2(G16), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G4), .B2(G16), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n691), .A2(new_n729), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(new_n730), .B2(new_n732), .ZN(new_n734));
  NOR2_X1   g309(.A1(G5), .A2(G16), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G171), .B2(G16), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G1961), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT30), .B(G28), .ZN(new_n738));
  OR2_X1    g313(.A1(KEYINPUT31), .A2(G11), .ZN(new_n739));
  NAND2_X1  g314(.A1(KEYINPUT31), .A2(G11), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n738), .A2(new_n687), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n617), .A2(G29), .A3(new_n621), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n741), .B1(new_n742), .B2(KEYINPUT98), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(KEYINPUT98), .B2(new_n742), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT93), .B(KEYINPUT28), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n687), .A2(G26), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n488), .A2(G140), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n489), .A2(G128), .ZN(new_n749));
  OAI221_X1 g324(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n463), .C2(G116), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n747), .B1(new_n751), .B2(G29), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(G2067), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n744), .A2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(G1966), .ZN(new_n755));
  NOR2_X1   g330(.A1(G168), .A2(new_n681), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n681), .B2(G21), .ZN(new_n757));
  AOI211_X1 g332(.A(new_n737), .B(new_n754), .C1(new_n755), .C2(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(G27), .A2(G29), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G164), .B2(G29), .ZN(new_n760));
  INV_X1    g335(.A(G2078), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n681), .A2(G19), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(new_n557), .B2(new_n681), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(G1341), .Z(new_n765));
  NAND2_X1  g340(.A1(new_n687), .A2(G32), .ZN(new_n766));
  AOI22_X1  g341(.A1(G141), .A2(new_n488), .B1(new_n462), .B2(G105), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n489), .A2(G129), .ZN(new_n768));
  NAND3_X1  g343(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT26), .Z(new_n770));
  NAND3_X1  g345(.A1(new_n767), .A2(new_n768), .A3(new_n770), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT96), .Z(new_n772));
  OAI21_X1  g347(.A(new_n766), .B1(new_n772), .B2(new_n687), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT27), .B(G1996), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n758), .A2(new_n762), .A3(new_n765), .A4(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n757), .A2(new_n755), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT97), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT24), .ZN(new_n779));
  INV_X1    g354(.A(G34), .ZN(new_n780));
  AOI21_X1  g355(.A(G29), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n779), .B2(new_n780), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G160), .B2(new_n687), .ZN(new_n783));
  INV_X1    g358(.A(G2084), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n778), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(G29), .A2(G33), .ZN(new_n787));
  NAND2_X1  g362(.A1(G115), .A2(G2104), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n473), .A2(new_n475), .ZN(new_n789));
  INV_X1    g364(.A(G127), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT94), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n463), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n792), .B2(new_n791), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT25), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G139), .B2(new_n488), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT95), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n787), .B1(new_n799), .B2(G29), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G2072), .ZN(new_n801));
  NOR4_X1   g376(.A1(new_n734), .A2(new_n776), .A3(new_n786), .A4(new_n801), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n694), .A2(new_n728), .A3(new_n802), .ZN(G150));
  INV_X1    g378(.A(G150), .ZN(G311));
  NAND2_X1  g379(.A1(new_n598), .A2(G559), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT38), .Z(new_n806));
  NAND2_X1  g381(.A1(new_n547), .A2(G93), .ZN(new_n807));
  AOI22_X1  g382(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n808));
  INV_X1    g383(.A(G55), .ZN(new_n809));
  OAI221_X1 g384(.A(new_n807), .B1(new_n510), .B2(new_n808), .C1(new_n809), .C2(new_n538), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n556), .B(new_n810), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n806), .B(new_n811), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n812), .A2(KEYINPUT39), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n812), .A2(KEYINPUT39), .ZN(new_n814));
  NOR3_X1   g389(.A1(new_n813), .A2(new_n814), .A3(G860), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n810), .A2(G860), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT37), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n815), .A2(new_n817), .ZN(G145));
  XOR2_X1   g393(.A(new_n720), .B(KEYINPUT102), .Z(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(new_n611), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n488), .A2(G142), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n489), .A2(G130), .ZN(new_n822));
  OAI221_X1 g397(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n463), .C2(G118), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n820), .B(new_n824), .Z(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT103), .Z(new_n826));
  INV_X1    g401(.A(new_n772), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT101), .ZN(new_n828));
  AND2_X1   g403(.A1(new_n799), .A2(new_n828), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n829), .A2(new_n751), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n751), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n827), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n830), .A2(new_n827), .A3(new_n831), .ZN(new_n834));
  AOI21_X1  g409(.A(G164), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n834), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n498), .A2(new_n500), .A3(new_n502), .A4(G138), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n504), .B1(new_n789), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n505), .A2(KEYINPUT4), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n838), .A2(new_n508), .A3(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n497), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NOR3_X1   g417(.A1(new_n836), .A2(new_n832), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n826), .B1(new_n835), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n842), .B1(new_n836), .B2(new_n832), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n833), .A2(new_n834), .A3(G164), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n825), .B(KEYINPUT103), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n844), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n492), .B(G160), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n622), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(G37), .B1(new_n849), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n825), .B1(new_n835), .B2(new_n843), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n854), .A2(new_n848), .A3(new_n851), .ZN(new_n855));
  AOI21_X1  g430(.A(KEYINPUT40), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n848), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n847), .B1(new_n845), .B2(new_n846), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n852), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(G37), .ZN(new_n860));
  AND4_X1   g435(.A1(KEYINPUT40), .A2(new_n859), .A3(new_n860), .A4(new_n855), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n856), .A2(new_n861), .ZN(G395));
  XNOR2_X1  g437(.A(G288), .B(KEYINPUT104), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n584), .ZN(new_n864));
  XNOR2_X1  g439(.A(G166), .B(G290), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT42), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n598), .B(G299), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n868), .A2(KEYINPUT41), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(KEYINPUT41), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n811), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n606), .B(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n874), .B1(new_n868), .B2(new_n873), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n867), .B(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(G868), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n810), .A2(new_n590), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(G331));
  INV_X1    g454(.A(KEYINPUT105), .ZN(new_n880));
  XNOR2_X1  g455(.A(G331), .B(new_n880), .ZN(G295));
  INV_X1    g456(.A(KEYINPUT44), .ZN(new_n882));
  NOR2_X1   g457(.A1(G168), .A2(G171), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n884), .B1(G301), .B2(G286), .ZN(new_n885));
  AND2_X1   g460(.A1(new_n885), .A2(new_n872), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n885), .A2(new_n872), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n888), .A2(new_n869), .A3(new_n870), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n868), .B1(new_n886), .B2(new_n887), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n866), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OR3_X1    g466(.A1(new_n891), .A2(KEYINPUT106), .A3(G37), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n889), .A2(new_n890), .ZN(new_n893));
  AOI21_X1  g468(.A(KEYINPUT43), .B1(new_n893), .B2(new_n866), .ZN(new_n894));
  OAI21_X1  g469(.A(KEYINPUT106), .B1(new_n891), .B2(G37), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n892), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n891), .A2(G37), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n893), .A2(new_n866), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(KEYINPUT43), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n882), .B1(new_n896), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n892), .A2(new_n895), .A3(new_n898), .ZN(new_n902));
  AOI22_X1  g477(.A1(new_n902), .A2(KEYINPUT43), .B1(new_n897), .B2(new_n894), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n901), .B1(new_n903), .B2(new_n882), .ZN(G397));
  INV_X1    g479(.A(KEYINPUT45), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n905), .B1(G164), .B2(G1384), .ZN(new_n906));
  OAI211_X1 g481(.A(G40), .B(new_n469), .C1(new_n480), .C2(new_n481), .ZN(new_n907));
  OR3_X1    g482(.A1(new_n906), .A2(KEYINPUT107), .A3(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(KEYINPUT107), .B1(new_n906), .B2(new_n907), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OR2_X1    g485(.A1(new_n910), .A2(G1996), .ZN(new_n911));
  OR2_X1    g486(.A1(new_n911), .A2(new_n827), .ZN(new_n912));
  INV_X1    g487(.A(new_n910), .ZN(new_n913));
  INV_X1    g488(.A(G2067), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n751), .B(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n915), .B(KEYINPUT108), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(new_n772), .ZN(new_n917));
  INV_X1    g492(.A(new_n916), .ZN(new_n918));
  OAI211_X1 g493(.A(new_n913), .B(new_n917), .C1(G1996), .C2(new_n918), .ZN(new_n919));
  XOR2_X1   g494(.A(new_n720), .B(new_n723), .Z(new_n920));
  NAND2_X1  g495(.A1(new_n913), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n912), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(G290), .B(new_n714), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n923), .B1(new_n910), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT61), .ZN(new_n926));
  NOR2_X1   g501(.A1(G299), .A2(KEYINPUT57), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT57), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n928), .B1(new_n566), .B2(new_n568), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT109), .ZN(new_n931));
  INV_X1    g506(.A(G1384), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n931), .B1(new_n842), .B2(new_n932), .ZN(new_n933));
  AOI211_X1 g508(.A(KEYINPUT109), .B(G1384), .C1(new_n840), .C2(new_n841), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT50), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT50), .ZN(new_n936));
  AOI21_X1  g511(.A(G1384), .B1(new_n840), .B2(new_n841), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n907), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n907), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n937), .A2(KEYINPUT45), .ZN(new_n941));
  XNOR2_X1  g516(.A(KEYINPUT56), .B(G2072), .ZN(new_n942));
  AND4_X1   g517(.A1(new_n906), .A2(new_n940), .A3(new_n941), .A4(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT113), .ZN(new_n944));
  AOI22_X1  g519(.A1(new_n685), .A2(new_n939), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n906), .A2(new_n940), .A3(new_n941), .A4(new_n942), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(KEYINPUT113), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n930), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(KEYINPUT109), .B1(G164), .B2(G1384), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n937), .A2(new_n931), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n936), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n937), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n940), .B1(KEYINPUT50), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n685), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n907), .B1(KEYINPUT45), .B2(new_n937), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n955), .A2(new_n944), .A3(new_n906), .A4(new_n942), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n954), .A2(new_n930), .A3(new_n947), .A4(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n926), .B1(new_n948), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n954), .A2(new_n947), .A3(new_n956), .ZN(new_n960));
  INV_X1    g535(.A(new_n930), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n926), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n945), .A2(KEYINPUT117), .A3(new_n930), .A4(new_n947), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT117), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n957), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n962), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n949), .A2(new_n940), .A3(new_n950), .ZN(new_n967));
  XOR2_X1   g542(.A(KEYINPUT58), .B(G1341), .Z(new_n968));
  AND2_X1   g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n940), .A2(new_n941), .ZN(new_n970));
  INV_X1    g545(.A(new_n906), .ZN(new_n971));
  NOR3_X1   g546(.A1(new_n970), .A2(new_n971), .A3(G1996), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n557), .B1(new_n969), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(KEYINPUT59), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT59), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n975), .B(new_n557), .C1(new_n969), .C2(new_n972), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n959), .A2(new_n966), .A3(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT118), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n959), .A2(new_n966), .A3(KEYINPUT118), .A4(new_n977), .ZN(new_n981));
  NOR3_X1   g556(.A1(new_n933), .A2(new_n934), .A3(KEYINPUT50), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n940), .B1(new_n936), .B2(new_n937), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n730), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(KEYINPUT114), .B1(new_n967), .B2(G2067), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n933), .A2(new_n934), .A3(new_n907), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT114), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n986), .A2(new_n987), .A3(new_n914), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n984), .A2(new_n985), .A3(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT60), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OR2_X1    g566(.A1(new_n989), .A2(new_n990), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n992), .A2(new_n598), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n992), .A2(new_n598), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n991), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n980), .A2(new_n981), .A3(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT116), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n989), .A2(KEYINPUT115), .A3(new_n598), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n960), .A2(new_n961), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(KEYINPUT115), .B1(new_n989), .B2(new_n598), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n997), .B(new_n957), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n989), .A2(new_n598), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT115), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1006), .A2(new_n999), .A3(new_n998), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n997), .B1(new_n1007), .B2(new_n957), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1003), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n996), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(G1961), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1011), .B1(new_n982), .B2(new_n983), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n905), .B1(new_n933), .B2(new_n934), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT53), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1014), .A2(G2078), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1013), .A2(new_n955), .A3(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n955), .A2(new_n761), .A3(new_n906), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT121), .ZN(new_n1018));
  AND3_X1   g593(.A1(new_n1017), .A2(new_n1018), .A3(new_n1014), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1018), .B1(new_n1017), .B2(new_n1014), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1012), .B(new_n1016), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G301), .ZN(new_n1022));
  AND3_X1   g597(.A1(new_n1021), .A2(KEYINPUT122), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT122), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n469), .A2(G40), .A3(new_n1015), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1026), .B1(new_n479), .B2(new_n478), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n906), .A2(new_n941), .A3(new_n1027), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1012), .B(new_n1028), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1029));
  OR2_X1    g604(.A1(new_n1029), .A2(new_n1022), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT54), .B1(new_n1025), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n705), .A2(G1976), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n967), .A2(G8), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT52), .ZN(new_n1034));
  INV_X1    g609(.A(G1976), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT52), .B1(G288), .B2(new_n1035), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n967), .A2(G8), .A3(new_n1032), .A4(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT111), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n515), .A2(G61), .ZN(new_n1039));
  OAI21_X1  g614(.A(G651), .B1(new_n1039), .B2(new_n577), .ZN(new_n1040));
  INV_X1    g615(.A(G1981), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1040), .A2(new_n1041), .A3(new_n581), .A4(new_n582), .ZN(new_n1042));
  OAI21_X1  g617(.A(G1981), .B1(new_n580), .B2(new_n583), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1038), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g619(.A(new_n1044), .B(KEYINPUT49), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1045), .A2(G8), .A3(new_n967), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1034), .A2(new_n1037), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G8), .ZN(new_n1048));
  NOR2_X1   g623(.A1(G166), .A2(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g624(.A(KEYINPUT110), .B(KEYINPUT55), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n1049), .B(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n949), .A2(new_n936), .A3(new_n950), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n907), .B1(new_n952), .B2(KEYINPUT50), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1052), .A2(new_n729), .A3(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n701), .B1(new_n970), .B2(new_n971), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1048), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1047), .B1(new_n1051), .B2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n935), .A2(new_n729), .A3(new_n938), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1048), .B1(new_n1058), .B2(new_n1055), .ZN(new_n1059));
  OR3_X1    g634(.A1(new_n1059), .A2(KEYINPUT112), .A3(new_n1051), .ZN(new_n1060));
  OAI21_X1  g635(.A(KEYINPUT112), .B1(new_n1059), .B2(new_n1051), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1057), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1029), .A2(G171), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1064), .B(KEYINPUT54), .C1(new_n1022), .C2(new_n1021), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT45), .B1(new_n949), .B2(new_n950), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n755), .B1(new_n1066), .B2(new_n970), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1052), .A2(new_n784), .A3(new_n1053), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1048), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(G286), .ZN(new_n1070));
  NAND2_X1  g645(.A1(G286), .A2(G8), .ZN(new_n1071));
  XNOR2_X1  g646(.A(new_n1071), .B(KEYINPUT120), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT119), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1073), .B1(new_n1069), .B2(new_n1074), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n1052), .A2(new_n784), .A3(new_n1053), .ZN(new_n1076));
  AOI21_X1  g651(.A(G1966), .B1(new_n1013), .B2(new_n955), .ZN(new_n1077));
  OAI21_X1  g652(.A(G8), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1078), .A2(KEYINPUT119), .ZN(new_n1079));
  OAI211_X1 g654(.A(KEYINPUT51), .B(new_n1070), .C1(new_n1075), .C2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1071), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n1069), .A2(KEYINPUT51), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1063), .A2(new_n1065), .A3(new_n1080), .A4(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1031), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1010), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT62), .ZN(new_n1087));
  OAI21_X1  g662(.A(KEYINPUT51), .B1(new_n1078), .B2(G168), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1069), .A2(new_n1074), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1072), .B1(new_n1078), .B2(KEYINPUT119), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1088), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1087), .B1(new_n1091), .B2(new_n1082), .ZN(new_n1092));
  OR2_X1    g667(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1080), .A2(KEYINPUT62), .A3(new_n1083), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1092), .A2(new_n1093), .A3(new_n1094), .A4(new_n1063), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1056), .A2(new_n1051), .ZN(new_n1096));
  NOR2_X1   g671(.A1(G288), .A2(G1976), .ZN(new_n1097));
  AOI22_X1  g672(.A1(new_n1046), .A2(new_n1097), .B1(new_n1041), .B2(new_n584), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n967), .A2(G8), .ZN(new_n1099));
  OAI22_X1  g674(.A1(new_n1096), .A2(new_n1047), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT63), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1069), .A2(G168), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1101), .B1(new_n1062), .B2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1102), .A2(new_n1101), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1104), .B(new_n1057), .C1(new_n1051), .C2(new_n1056), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1100), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n1095), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n925), .B1(new_n1086), .B2(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(new_n911), .B(KEYINPUT46), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n913), .A2(new_n917), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT47), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1109), .A2(KEYINPUT47), .A3(new_n1110), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT123), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n912), .A2(new_n919), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n721), .A2(new_n723), .ZN(new_n1119));
  OAI22_X1  g694(.A1(new_n1118), .A2(new_n1119), .B1(G2067), .B2(new_n751), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n913), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1113), .A2(KEYINPUT123), .A3(new_n1114), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n923), .A2(KEYINPUT124), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT124), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n922), .A2(new_n1124), .ZN(new_n1125));
  NOR3_X1   g700(.A1(new_n910), .A2(G1986), .A3(G290), .ZN(new_n1126));
  XOR2_X1   g701(.A(new_n1126), .B(KEYINPUT48), .Z(new_n1127));
  NAND3_X1  g702(.A1(new_n1123), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1117), .A2(new_n1121), .A3(new_n1122), .A4(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(KEYINPUT125), .B1(new_n1108), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1129), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT125), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1095), .A2(new_n1106), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1133), .B1(new_n1010), .B2(new_n1085), .ZN(new_n1134));
  OAI211_X1 g709(.A(new_n1131), .B(new_n1132), .C1(new_n1134), .C2(new_n925), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1130), .A2(new_n1135), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g711(.A1(new_n902), .A2(KEYINPUT43), .ZN(new_n1138));
  NAND2_X1  g712(.A1(new_n894), .A2(new_n897), .ZN(new_n1139));
  NAND2_X1  g713(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g714(.A1(new_n853), .A2(new_n855), .ZN(new_n1141));
  INV_X1    g715(.A(G319), .ZN(new_n1142));
  NOR3_X1   g716(.A1(new_n643), .A2(new_n1142), .A3(G227), .ZN(new_n1143));
  OAI21_X1  g717(.A(new_n1143), .B1(new_n678), .B2(new_n679), .ZN(new_n1144));
  INV_X1    g718(.A(KEYINPUT126), .ZN(new_n1145));
  NAND2_X1  g719(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  OAI211_X1 g720(.A(KEYINPUT126), .B(new_n1143), .C1(new_n678), .C2(new_n679), .ZN(new_n1147));
  NAND2_X1  g721(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  AND3_X1   g722(.A1(new_n1140), .A2(new_n1141), .A3(new_n1148), .ZN(G308));
  NAND3_X1  g723(.A1(new_n1140), .A2(new_n1141), .A3(new_n1148), .ZN(G225));
endmodule


