

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U557 ( .A1(G2105), .A2(G2104), .ZN(n543) );
  NAND2_X1 U558 ( .A1(n527), .A2(n752), .ZN(n747) );
  NOR2_X1 U559 ( .A1(G651), .A2(n579), .ZN(n794) );
  XOR2_X1 U560 ( .A(n654), .B(KEYINPUT28), .Z(n525) );
  XOR2_X1 U561 ( .A(KEYINPUT101), .B(n679), .Z(n526) );
  XNOR2_X1 U562 ( .A(n728), .B(KEYINPUT92), .ZN(n527) );
  INV_X1 U563 ( .A(n664), .ZN(n640) );
  XNOR2_X1 U564 ( .A(n673), .B(KEYINPUT32), .ZN(n680) );
  NAND2_X1 U565 ( .A1(n725), .A2(n596), .ZN(n664) );
  OR2_X1 U566 ( .A1(n766), .A2(n595), .ZN(n726) );
  INV_X1 U567 ( .A(KEYINPUT13), .ZN(n624) );
  OR2_X1 U568 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U569 ( .A(n624), .B(KEYINPUT71), .ZN(n625) );
  NOR2_X1 U570 ( .A1(n579), .A2(n535), .ZN(n798) );
  XNOR2_X1 U571 ( .A(n626), .B(n625), .ZN(n627) );
  NOR2_X2 U572 ( .A1(G2105), .A2(n547), .ZN(n888) );
  NOR2_X1 U573 ( .A1(G543), .A2(G651), .ZN(n799) );
  XNOR2_X1 U574 ( .A(KEYINPUT74), .B(KEYINPUT6), .ZN(n532) );
  INV_X1 U575 ( .A(G651), .ZN(n535) );
  NOR2_X1 U576 ( .A1(G543), .A2(n535), .ZN(n528) );
  XOR2_X1 U577 ( .A(KEYINPUT1), .B(n528), .Z(n793) );
  NAND2_X1 U578 ( .A1(G63), .A2(n793), .ZN(n530) );
  XOR2_X1 U579 ( .A(G543), .B(KEYINPUT0), .Z(n579) );
  NAND2_X1 U580 ( .A1(G51), .A2(n794), .ZN(n529) );
  NAND2_X1 U581 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U582 ( .A(n532), .B(n531), .ZN(n540) );
  NAND2_X1 U583 ( .A1(G89), .A2(n799), .ZN(n533) );
  XOR2_X1 U584 ( .A(KEYINPUT73), .B(n533), .Z(n534) );
  XNOR2_X1 U585 ( .A(n534), .B(KEYINPUT4), .ZN(n537) );
  NAND2_X1 U586 ( .A1(G76), .A2(n798), .ZN(n536) );
  NAND2_X1 U587 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U588 ( .A(KEYINPUT5), .B(n538), .Z(n539) );
  NOR2_X1 U589 ( .A1(n540), .A2(n539), .ZN(n542) );
  XNOR2_X1 U590 ( .A(KEYINPUT75), .B(KEYINPUT7), .ZN(n541) );
  XNOR2_X1 U591 ( .A(n542), .B(n541), .ZN(G168) );
  INV_X1 U592 ( .A(G2104), .ZN(n547) );
  NAND2_X1 U593 ( .A1(n888), .A2(G102), .ZN(n546) );
  XOR2_X1 U594 ( .A(KEYINPUT17), .B(n543), .Z(n544) );
  XNOR2_X1 U595 ( .A(n544), .B(KEYINPUT64), .ZN(n865) );
  NAND2_X1 U596 ( .A1(G138), .A2(n865), .ZN(n545) );
  NAND2_X1 U597 ( .A1(n546), .A2(n545), .ZN(n551) );
  AND2_X1 U598 ( .A1(n547), .A2(G2105), .ZN(n892) );
  NAND2_X1 U599 ( .A1(G126), .A2(n892), .ZN(n549) );
  AND2_X1 U600 ( .A1(G2105), .A2(G2104), .ZN(n893) );
  NAND2_X1 U601 ( .A1(G114), .A2(n893), .ZN(n548) );
  NAND2_X1 U602 ( .A1(n549), .A2(n548), .ZN(n550) );
  NOR2_X1 U603 ( .A1(n551), .A2(n550), .ZN(G164) );
  NAND2_X1 U604 ( .A1(G64), .A2(n793), .ZN(n553) );
  NAND2_X1 U605 ( .A1(G52), .A2(n794), .ZN(n552) );
  NAND2_X1 U606 ( .A1(n553), .A2(n552), .ZN(n558) );
  NAND2_X1 U607 ( .A1(G77), .A2(n798), .ZN(n555) );
  NAND2_X1 U608 ( .A1(G90), .A2(n799), .ZN(n554) );
  NAND2_X1 U609 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U610 ( .A(KEYINPUT9), .B(n556), .Z(n557) );
  NOR2_X1 U611 ( .A1(n558), .A2(n557), .ZN(G171) );
  INV_X1 U612 ( .A(G171), .ZN(G301) );
  XOR2_X1 U613 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U614 ( .A1(G75), .A2(n798), .ZN(n560) );
  NAND2_X1 U615 ( .A1(G88), .A2(n799), .ZN(n559) );
  NAND2_X1 U616 ( .A1(n560), .A2(n559), .ZN(n564) );
  NAND2_X1 U617 ( .A1(G62), .A2(n793), .ZN(n562) );
  NAND2_X1 U618 ( .A1(G50), .A2(n794), .ZN(n561) );
  NAND2_X1 U619 ( .A1(n562), .A2(n561), .ZN(n563) );
  NOR2_X1 U620 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U621 ( .A(n565), .B(KEYINPUT83), .Z(G166) );
  INV_X1 U622 ( .A(G166), .ZN(G303) );
  NAND2_X1 U623 ( .A1(G48), .A2(n794), .ZN(n566) );
  XNOR2_X1 U624 ( .A(n566), .B(KEYINPUT82), .ZN(n575) );
  NAND2_X1 U625 ( .A1(G73), .A2(n798), .ZN(n567) );
  XOR2_X1 U626 ( .A(KEYINPUT2), .B(n567), .Z(n568) );
  XNOR2_X1 U627 ( .A(n568), .B(KEYINPUT81), .ZN(n570) );
  NAND2_X1 U628 ( .A1(G61), .A2(n793), .ZN(n569) );
  NAND2_X1 U629 ( .A1(n570), .A2(n569), .ZN(n573) );
  NAND2_X1 U630 ( .A1(n799), .A2(G86), .ZN(n571) );
  XOR2_X1 U631 ( .A(KEYINPUT80), .B(n571), .Z(n572) );
  NOR2_X1 U632 ( .A1(n573), .A2(n572), .ZN(n574) );
  NAND2_X1 U633 ( .A1(n575), .A2(n574), .ZN(G305) );
  NAND2_X1 U634 ( .A1(G49), .A2(n794), .ZN(n577) );
  NAND2_X1 U635 ( .A1(G74), .A2(G651), .ZN(n576) );
  NAND2_X1 U636 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U637 ( .A1(n793), .A2(n578), .ZN(n581) );
  NAND2_X1 U638 ( .A1(n579), .A2(G87), .ZN(n580) );
  NAND2_X1 U639 ( .A1(n581), .A2(n580), .ZN(G288) );
  NAND2_X1 U640 ( .A1(G60), .A2(n793), .ZN(n583) );
  NAND2_X1 U641 ( .A1(G47), .A2(n794), .ZN(n582) );
  NAND2_X1 U642 ( .A1(n583), .A2(n582), .ZN(n586) );
  NAND2_X1 U643 ( .A1(G72), .A2(n798), .ZN(n584) );
  XNOR2_X1 U644 ( .A(KEYINPUT65), .B(n584), .ZN(n585) );
  NOR2_X1 U645 ( .A1(n586), .A2(n585), .ZN(n588) );
  NAND2_X1 U646 ( .A1(n799), .A2(G85), .ZN(n587) );
  NAND2_X1 U647 ( .A1(n588), .A2(n587), .ZN(G290) );
  NOR2_X1 U648 ( .A1(G164), .A2(G1384), .ZN(n725) );
  NAND2_X1 U649 ( .A1(G137), .A2(n865), .ZN(n591) );
  NAND2_X1 U650 ( .A1(G101), .A2(n888), .ZN(n589) );
  XOR2_X1 U651 ( .A(KEYINPUT23), .B(n589), .Z(n590) );
  NAND2_X1 U652 ( .A1(n591), .A2(n590), .ZN(n766) );
  NAND2_X1 U653 ( .A1(G125), .A2(n892), .ZN(n593) );
  NAND2_X1 U654 ( .A1(G113), .A2(n893), .ZN(n592) );
  NAND2_X1 U655 ( .A1(n593), .A2(n592), .ZN(n767) );
  INV_X1 U656 ( .A(G40), .ZN(n594) );
  OR2_X1 U657 ( .A1(n767), .A2(n594), .ZN(n595) );
  XOR2_X1 U658 ( .A(KEYINPUT96), .B(n726), .Z(n596) );
  NAND2_X1 U659 ( .A1(n664), .A2(G8), .ZN(n698) );
  NOR2_X1 U660 ( .A1(G1966), .A2(n698), .ZN(n674) );
  NOR2_X1 U661 ( .A1(G2084), .A2(n664), .ZN(n676) );
  NOR2_X1 U662 ( .A1(n674), .A2(n676), .ZN(n597) );
  XNOR2_X1 U663 ( .A(n597), .B(KEYINPUT100), .ZN(n598) );
  NAND2_X1 U664 ( .A1(n598), .A2(G8), .ZN(n599) );
  XNOR2_X1 U665 ( .A(KEYINPUT30), .B(n599), .ZN(n600) );
  NOR2_X1 U666 ( .A1(G168), .A2(n600), .ZN(n604) );
  NAND2_X1 U667 ( .A1(G1961), .A2(n664), .ZN(n602) );
  XOR2_X1 U668 ( .A(KEYINPUT25), .B(G2078), .Z(n1014) );
  NAND2_X1 U669 ( .A1(n640), .A2(n1014), .ZN(n601) );
  NAND2_X1 U670 ( .A1(n602), .A2(n601), .ZN(n657) );
  AND2_X1 U671 ( .A1(G301), .A2(n657), .ZN(n603) );
  NOR2_X1 U672 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U673 ( .A(n605), .B(KEYINPUT31), .ZN(n661) );
  NAND2_X1 U674 ( .A1(n799), .A2(G92), .ZN(n612) );
  NAND2_X1 U675 ( .A1(G66), .A2(n793), .ZN(n607) );
  NAND2_X1 U676 ( .A1(G54), .A2(n794), .ZN(n606) );
  NAND2_X1 U677 ( .A1(n607), .A2(n606), .ZN(n610) );
  NAND2_X1 U678 ( .A1(n798), .A2(G79), .ZN(n608) );
  XOR2_X1 U679 ( .A(KEYINPUT72), .B(n608), .Z(n609) );
  NOR2_X1 U680 ( .A1(n610), .A2(n609), .ZN(n611) );
  NAND2_X1 U681 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U682 ( .A(KEYINPUT15), .B(n613), .ZN(n931) );
  INV_X1 U683 ( .A(n931), .ZN(n779) );
  NAND2_X1 U684 ( .A1(G1348), .A2(n664), .ZN(n615) );
  NAND2_X1 U685 ( .A1(G2067), .A2(n640), .ZN(n614) );
  NAND2_X1 U686 ( .A1(n615), .A2(n614), .ZN(n618) );
  NOR2_X1 U687 ( .A1(n779), .A2(n618), .ZN(n638) );
  XOR2_X1 U688 ( .A(KEYINPUT26), .B(KEYINPUT98), .Z(n617) );
  NAND2_X1 U689 ( .A1(n640), .A2(G1996), .ZN(n616) );
  XNOR2_X1 U690 ( .A(n617), .B(n616), .ZN(n636) );
  NAND2_X1 U691 ( .A1(n779), .A2(n618), .ZN(n634) );
  NAND2_X1 U692 ( .A1(n793), .A2(G56), .ZN(n619) );
  XOR2_X1 U693 ( .A(KEYINPUT14), .B(n619), .Z(n628) );
  NAND2_X1 U694 ( .A1(n799), .A2(G81), .ZN(n620) );
  XOR2_X1 U695 ( .A(KEYINPUT12), .B(n620), .Z(n623) );
  NAND2_X1 U696 ( .A1(n798), .A2(G68), .ZN(n621) );
  XOR2_X1 U697 ( .A(n621), .B(KEYINPUT70), .Z(n622) );
  NOR2_X1 U698 ( .A1(n623), .A2(n622), .ZN(n626) );
  NOR2_X1 U699 ( .A1(n628), .A2(n627), .ZN(n630) );
  NAND2_X1 U700 ( .A1(n794), .A2(G43), .ZN(n629) );
  NAND2_X1 U701 ( .A1(n630), .A2(n629), .ZN(n943) );
  NAND2_X1 U702 ( .A1(G1341), .A2(n664), .ZN(n631) );
  XNOR2_X1 U703 ( .A(KEYINPUT99), .B(n631), .ZN(n632) );
  NOR2_X1 U704 ( .A1(n943), .A2(n632), .ZN(n633) );
  NAND2_X1 U705 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U706 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U707 ( .A1(n638), .A2(n637), .ZN(n652) );
  NAND2_X1 U708 ( .A1(n640), .A2(G2072), .ZN(n639) );
  XNOR2_X1 U709 ( .A(n639), .B(KEYINPUT27), .ZN(n642) );
  INV_X1 U710 ( .A(G1956), .ZN(n929) );
  NOR2_X1 U711 ( .A1(n929), .A2(n640), .ZN(n641) );
  NOR2_X1 U712 ( .A1(n642), .A2(n641), .ZN(n653) );
  NAND2_X1 U713 ( .A1(G65), .A2(n793), .ZN(n644) );
  NAND2_X1 U714 ( .A1(G53), .A2(n794), .ZN(n643) );
  NAND2_X1 U715 ( .A1(n644), .A2(n643), .ZN(n650) );
  NAND2_X1 U716 ( .A1(n799), .A2(G91), .ZN(n645) );
  XNOR2_X1 U717 ( .A(n645), .B(KEYINPUT66), .ZN(n647) );
  NAND2_X1 U718 ( .A1(G78), .A2(n798), .ZN(n646) );
  NAND2_X1 U719 ( .A1(n647), .A2(n646), .ZN(n648) );
  XOR2_X1 U720 ( .A(KEYINPUT67), .B(n648), .Z(n649) );
  NOR2_X1 U721 ( .A1(n650), .A2(n649), .ZN(n930) );
  NAND2_X1 U722 ( .A1(n653), .A2(n930), .ZN(n651) );
  NAND2_X1 U723 ( .A1(n652), .A2(n651), .ZN(n655) );
  NOR2_X1 U724 ( .A1(n653), .A2(n930), .ZN(n654) );
  NAND2_X1 U725 ( .A1(n655), .A2(n525), .ZN(n656) );
  XNOR2_X1 U726 ( .A(n656), .B(KEYINPUT29), .ZN(n659) );
  NOR2_X1 U727 ( .A1(G301), .A2(n657), .ZN(n658) );
  NOR2_X1 U728 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U729 ( .A1(n661), .A2(n660), .ZN(n675) );
  INV_X1 U730 ( .A(n675), .ZN(n663) );
  AND2_X1 U731 ( .A1(G286), .A2(G8), .ZN(n662) );
  NAND2_X1 U732 ( .A1(n663), .A2(n662), .ZN(n672) );
  INV_X1 U733 ( .A(G8), .ZN(n670) );
  NOR2_X1 U734 ( .A1(G1971), .A2(n698), .ZN(n666) );
  NOR2_X1 U735 ( .A1(G2090), .A2(n664), .ZN(n665) );
  NOR2_X1 U736 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U737 ( .A1(n667), .A2(G303), .ZN(n668) );
  XNOR2_X1 U738 ( .A(n668), .B(KEYINPUT102), .ZN(n669) );
  OR2_X1 U739 ( .A1(n670), .A2(n669), .ZN(n671) );
  AND2_X1 U740 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U741 ( .A1(n675), .A2(n674), .ZN(n678) );
  NAND2_X1 U742 ( .A1(G8), .A2(n676), .ZN(n677) );
  NAND2_X1 U743 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U744 ( .A1(n680), .A2(n526), .ZN(n691) );
  NAND2_X1 U745 ( .A1(G8), .A2(G166), .ZN(n681) );
  NOR2_X1 U746 ( .A1(G2090), .A2(n681), .ZN(n682) );
  XNOR2_X1 U747 ( .A(n682), .B(KEYINPUT105), .ZN(n683) );
  NAND2_X1 U748 ( .A1(n691), .A2(n683), .ZN(n684) );
  XNOR2_X1 U749 ( .A(n684), .B(KEYINPUT106), .ZN(n685) );
  NAND2_X1 U750 ( .A1(n685), .A2(n698), .ZN(n690) );
  NOR2_X1 U751 ( .A1(G1981), .A2(G305), .ZN(n686) );
  XOR2_X1 U752 ( .A(n686), .B(KEYINPUT24), .Z(n687) );
  NOR2_X1 U753 ( .A1(n698), .A2(n687), .ZN(n688) );
  XNOR2_X1 U754 ( .A(KEYINPUT97), .B(n688), .ZN(n689) );
  NAND2_X1 U755 ( .A1(n690), .A2(n689), .ZN(n712) );
  INV_X1 U756 ( .A(n691), .ZN(n695) );
  NOR2_X1 U757 ( .A1(G1976), .A2(G288), .ZN(n697) );
  NOR2_X1 U758 ( .A1(G1971), .A2(G303), .ZN(n692) );
  NOR2_X1 U759 ( .A1(n697), .A2(n692), .ZN(n693) );
  XNOR2_X1 U760 ( .A(n693), .B(KEYINPUT103), .ZN(n694) );
  NOR2_X1 U761 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U762 ( .A1(n696), .A2(n698), .ZN(n704) );
  NAND2_X1 U763 ( .A1(G1976), .A2(G288), .ZN(n937) );
  INV_X1 U764 ( .A(KEYINPUT33), .ZN(n706) );
  INV_X1 U765 ( .A(n697), .ZN(n936) );
  OR2_X1 U766 ( .A1(n936), .A2(n698), .ZN(n699) );
  NOR2_X1 U767 ( .A1(n706), .A2(n699), .ZN(n700) );
  XOR2_X1 U768 ( .A(n700), .B(KEYINPUT104), .Z(n705) );
  AND2_X1 U769 ( .A1(n937), .A2(n705), .ZN(n702) );
  XNOR2_X1 U770 ( .A(G1981), .B(G305), .ZN(n949) );
  INV_X1 U771 ( .A(n949), .ZN(n701) );
  AND2_X1 U772 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U773 ( .A1(n704), .A2(n703), .ZN(n710) );
  INV_X1 U774 ( .A(n705), .ZN(n707) );
  OR2_X1 U775 ( .A1(n707), .A2(n706), .ZN(n708) );
  OR2_X1 U776 ( .A1(n949), .A2(n708), .ZN(n709) );
  NAND2_X1 U777 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U778 ( .A1(n712), .A2(n711), .ZN(n748) );
  XOR2_X1 U779 ( .A(G2067), .B(KEYINPUT37), .Z(n713) );
  XNOR2_X1 U780 ( .A(KEYINPUT89), .B(n713), .ZN(n759) );
  XNOR2_X1 U781 ( .A(KEYINPUT91), .B(KEYINPUT36), .ZN(n724) );
  NAND2_X1 U782 ( .A1(G128), .A2(n892), .ZN(n715) );
  NAND2_X1 U783 ( .A1(G116), .A2(n893), .ZN(n714) );
  NAND2_X1 U784 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U785 ( .A(KEYINPUT35), .B(n716), .ZN(n722) );
  NAND2_X1 U786 ( .A1(n888), .A2(G104), .ZN(n718) );
  BUF_X1 U787 ( .A(n865), .Z(n889) );
  NAND2_X1 U788 ( .A1(G140), .A2(n889), .ZN(n717) );
  NAND2_X1 U789 ( .A1(n718), .A2(n717), .ZN(n720) );
  XOR2_X1 U790 ( .A(KEYINPUT90), .B(KEYINPUT34), .Z(n719) );
  XNOR2_X1 U791 ( .A(n720), .B(n719), .ZN(n721) );
  NAND2_X1 U792 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U793 ( .A(n724), .B(n723), .ZN(n902) );
  NOR2_X1 U794 ( .A1(n759), .A2(n902), .ZN(n1004) );
  NOR2_X1 U795 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U796 ( .A(n727), .B(KEYINPUT88), .ZN(n761) );
  NAND2_X1 U797 ( .A1(n1004), .A2(n761), .ZN(n728) );
  XOR2_X1 U798 ( .A(KEYINPUT94), .B(G1991), .Z(n1020) );
  NAND2_X1 U799 ( .A1(n893), .A2(G107), .ZN(n730) );
  NAND2_X1 U800 ( .A1(G131), .A2(n889), .ZN(n729) );
  NAND2_X1 U801 ( .A1(n730), .A2(n729), .ZN(n733) );
  NAND2_X1 U802 ( .A1(G119), .A2(n892), .ZN(n731) );
  XNOR2_X1 U803 ( .A(KEYINPUT93), .B(n731), .ZN(n732) );
  NOR2_X1 U804 ( .A1(n733), .A2(n732), .ZN(n735) );
  NAND2_X1 U805 ( .A1(n888), .A2(G95), .ZN(n734) );
  AND2_X1 U806 ( .A1(n735), .A2(n734), .ZN(n870) );
  NOR2_X1 U807 ( .A1(n1020), .A2(n870), .ZN(n745) );
  NAND2_X1 U808 ( .A1(G105), .A2(n888), .ZN(n736) );
  XOR2_X1 U809 ( .A(KEYINPUT38), .B(n736), .Z(n741) );
  NAND2_X1 U810 ( .A1(G129), .A2(n892), .ZN(n738) );
  NAND2_X1 U811 ( .A1(G117), .A2(n893), .ZN(n737) );
  NAND2_X1 U812 ( .A1(n738), .A2(n737), .ZN(n739) );
  XOR2_X1 U813 ( .A(KEYINPUT95), .B(n739), .Z(n740) );
  NOR2_X1 U814 ( .A1(n741), .A2(n740), .ZN(n743) );
  NAND2_X1 U815 ( .A1(G141), .A2(n889), .ZN(n742) );
  NAND2_X1 U816 ( .A1(n743), .A2(n742), .ZN(n877) );
  AND2_X1 U817 ( .A1(n877), .A2(G1996), .ZN(n744) );
  NOR2_X1 U818 ( .A1(n745), .A2(n744), .ZN(n994) );
  INV_X1 U819 ( .A(n994), .ZN(n746) );
  NAND2_X1 U820 ( .A1(n761), .A2(n746), .ZN(n752) );
  XNOR2_X1 U821 ( .A(n749), .B(KEYINPUT107), .ZN(n751) );
  XNOR2_X1 U822 ( .A(G1986), .B(G290), .ZN(n940) );
  NAND2_X1 U823 ( .A1(n940), .A2(n761), .ZN(n750) );
  NAND2_X1 U824 ( .A1(n751), .A2(n750), .ZN(n764) );
  NOR2_X1 U825 ( .A1(G1996), .A2(n877), .ZN(n989) );
  INV_X1 U826 ( .A(n752), .ZN(n755) );
  NOR2_X1 U827 ( .A1(G1986), .A2(G290), .ZN(n753) );
  AND2_X1 U828 ( .A1(n1020), .A2(n870), .ZN(n985) );
  NOR2_X1 U829 ( .A1(n753), .A2(n985), .ZN(n754) );
  NOR2_X1 U830 ( .A1(n755), .A2(n754), .ZN(n756) );
  NOR2_X1 U831 ( .A1(n989), .A2(n756), .ZN(n757) );
  XNOR2_X1 U832 ( .A(n757), .B(KEYINPUT39), .ZN(n758) );
  NAND2_X1 U833 ( .A1(n758), .A2(n527), .ZN(n760) );
  NAND2_X1 U834 ( .A1(n759), .A2(n902), .ZN(n1001) );
  NAND2_X1 U835 ( .A1(n760), .A2(n1001), .ZN(n762) );
  NAND2_X1 U836 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U837 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U838 ( .A(n765), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U839 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U840 ( .A(G57), .ZN(G237) );
  NOR2_X1 U841 ( .A1(n766), .A2(n767), .ZN(G160) );
  NAND2_X1 U842 ( .A1(G7), .A2(G661), .ZN(n768) );
  XOR2_X1 U843 ( .A(n768), .B(KEYINPUT10), .Z(n928) );
  NAND2_X1 U844 ( .A1(n928), .A2(G567), .ZN(n769) );
  XNOR2_X1 U845 ( .A(n769), .B(KEYINPUT11), .ZN(n770) );
  XNOR2_X1 U846 ( .A(KEYINPUT69), .B(n770), .ZN(G234) );
  INV_X1 U847 ( .A(G860), .ZN(n776) );
  OR2_X1 U848 ( .A1(n943), .A2(n776), .ZN(G153) );
  NAND2_X1 U849 ( .A1(G868), .A2(G301), .ZN(n772) );
  INV_X1 U850 ( .A(G868), .ZN(n812) );
  NAND2_X1 U851 ( .A1(n779), .A2(n812), .ZN(n771) );
  NAND2_X1 U852 ( .A1(n772), .A2(n771), .ZN(G284) );
  XOR2_X1 U853 ( .A(n930), .B(KEYINPUT68), .Z(G299) );
  NOR2_X1 U854 ( .A1(G299), .A2(G868), .ZN(n773) );
  XNOR2_X1 U855 ( .A(n773), .B(KEYINPUT76), .ZN(n775) );
  NOR2_X1 U856 ( .A1(n812), .A2(G286), .ZN(n774) );
  NOR2_X1 U857 ( .A1(n775), .A2(n774), .ZN(G297) );
  NAND2_X1 U858 ( .A1(n776), .A2(G559), .ZN(n777) );
  NAND2_X1 U859 ( .A1(n777), .A2(n931), .ZN(n778) );
  XNOR2_X1 U860 ( .A(n778), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U861 ( .A1(n779), .A2(n812), .ZN(n780) );
  XNOR2_X1 U862 ( .A(n780), .B(KEYINPUT77), .ZN(n781) );
  NOR2_X1 U863 ( .A1(G559), .A2(n781), .ZN(n783) );
  NOR2_X1 U864 ( .A1(G868), .A2(n943), .ZN(n782) );
  NOR2_X1 U865 ( .A1(n783), .A2(n782), .ZN(G282) );
  NAND2_X1 U866 ( .A1(n892), .A2(G123), .ZN(n784) );
  XNOR2_X1 U867 ( .A(n784), .B(KEYINPUT18), .ZN(n786) );
  NAND2_X1 U868 ( .A1(G111), .A2(n893), .ZN(n785) );
  NAND2_X1 U869 ( .A1(n786), .A2(n785), .ZN(n790) );
  NAND2_X1 U870 ( .A1(n888), .A2(G99), .ZN(n788) );
  NAND2_X1 U871 ( .A1(G135), .A2(n889), .ZN(n787) );
  NAND2_X1 U872 ( .A1(n788), .A2(n787), .ZN(n789) );
  NOR2_X1 U873 ( .A1(n790), .A2(n789), .ZN(n984) );
  XNOR2_X1 U874 ( .A(n984), .B(G2096), .ZN(n791) );
  INV_X1 U875 ( .A(G2100), .ZN(n841) );
  NAND2_X1 U876 ( .A1(n791), .A2(n841), .ZN(G156) );
  NAND2_X1 U877 ( .A1(G559), .A2(n931), .ZN(n792) );
  XNOR2_X1 U878 ( .A(n792), .B(n943), .ZN(n838) );
  NAND2_X1 U879 ( .A1(G67), .A2(n793), .ZN(n796) );
  NAND2_X1 U880 ( .A1(G55), .A2(n794), .ZN(n795) );
  NAND2_X1 U881 ( .A1(n796), .A2(n795), .ZN(n797) );
  XNOR2_X1 U882 ( .A(KEYINPUT78), .B(n797), .ZN(n803) );
  NAND2_X1 U883 ( .A1(G80), .A2(n798), .ZN(n801) );
  NAND2_X1 U884 ( .A1(G93), .A2(n799), .ZN(n800) );
  NAND2_X1 U885 ( .A1(n801), .A2(n800), .ZN(n802) );
  NOR2_X1 U886 ( .A1(n803), .A2(n802), .ZN(n804) );
  XNOR2_X1 U887 ( .A(KEYINPUT79), .B(n804), .ZN(n839) );
  XOR2_X1 U888 ( .A(G299), .B(n839), .Z(n810) );
  XNOR2_X1 U889 ( .A(KEYINPUT19), .B(KEYINPUT84), .ZN(n806) );
  XOR2_X1 U890 ( .A(G288), .B(G303), .Z(n805) );
  XNOR2_X1 U891 ( .A(n806), .B(n805), .ZN(n807) );
  XOR2_X1 U892 ( .A(n807), .B(G290), .Z(n808) );
  XNOR2_X1 U893 ( .A(G305), .B(n808), .ZN(n809) );
  XNOR2_X1 U894 ( .A(n810), .B(n809), .ZN(n907) );
  XNOR2_X1 U895 ( .A(n838), .B(n907), .ZN(n811) );
  NAND2_X1 U896 ( .A1(n811), .A2(G868), .ZN(n814) );
  NAND2_X1 U897 ( .A1(n839), .A2(n812), .ZN(n813) );
  NAND2_X1 U898 ( .A1(n814), .A2(n813), .ZN(G295) );
  NAND2_X1 U899 ( .A1(G2078), .A2(G2084), .ZN(n815) );
  XOR2_X1 U900 ( .A(KEYINPUT20), .B(n815), .Z(n816) );
  NAND2_X1 U901 ( .A1(G2090), .A2(n816), .ZN(n817) );
  XNOR2_X1 U902 ( .A(KEYINPUT21), .B(n817), .ZN(n818) );
  NAND2_X1 U903 ( .A1(n818), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U904 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U905 ( .A1(G69), .A2(G120), .ZN(n819) );
  NOR2_X1 U906 ( .A1(G237), .A2(n819), .ZN(n820) );
  NAND2_X1 U907 ( .A1(G108), .A2(n820), .ZN(n835) );
  NAND2_X1 U908 ( .A1(G567), .A2(n835), .ZN(n827) );
  XOR2_X1 U909 ( .A(KEYINPUT22), .B(KEYINPUT85), .Z(n822) );
  NAND2_X1 U910 ( .A1(G132), .A2(G82), .ZN(n821) );
  XNOR2_X1 U911 ( .A(n822), .B(n821), .ZN(n823) );
  NOR2_X1 U912 ( .A1(n823), .A2(G218), .ZN(n824) );
  XNOR2_X1 U913 ( .A(KEYINPUT86), .B(n824), .ZN(n825) );
  NAND2_X1 U914 ( .A1(n825), .A2(G96), .ZN(n836) );
  NAND2_X1 U915 ( .A1(G2106), .A2(n836), .ZN(n826) );
  NAND2_X1 U916 ( .A1(n827), .A2(n826), .ZN(n861) );
  NAND2_X1 U917 ( .A1(G661), .A2(G483), .ZN(n828) );
  XOR2_X1 U918 ( .A(KEYINPUT87), .B(n828), .Z(n829) );
  NOR2_X1 U919 ( .A1(n861), .A2(n829), .ZN(n834) );
  NAND2_X1 U920 ( .A1(n834), .A2(G36), .ZN(G176) );
  NAND2_X1 U921 ( .A1(G2106), .A2(n928), .ZN(G217) );
  NAND2_X1 U922 ( .A1(G15), .A2(G2), .ZN(n830) );
  XOR2_X1 U923 ( .A(KEYINPUT108), .B(n830), .Z(n831) );
  NAND2_X1 U924 ( .A1(n831), .A2(G661), .ZN(n832) );
  XOR2_X1 U925 ( .A(KEYINPUT109), .B(n832), .Z(G259) );
  NAND2_X1 U926 ( .A1(G3), .A2(G1), .ZN(n833) );
  NAND2_X1 U927 ( .A1(n834), .A2(n833), .ZN(G188) );
  INV_X1 U929 ( .A(G132), .ZN(G219) );
  INV_X1 U930 ( .A(G120), .ZN(G236) );
  INV_X1 U931 ( .A(G96), .ZN(G221) );
  INV_X1 U932 ( .A(G82), .ZN(G220) );
  INV_X1 U933 ( .A(G69), .ZN(G235) );
  NOR2_X1 U934 ( .A1(n836), .A2(n835), .ZN(n837) );
  XOR2_X1 U935 ( .A(n837), .B(KEYINPUT110), .Z(G261) );
  INV_X1 U936 ( .A(G261), .ZN(G325) );
  NOR2_X1 U937 ( .A1(n838), .A2(G860), .ZN(n840) );
  XOR2_X1 U938 ( .A(n840), .B(n839), .Z(G145) );
  XNOR2_X1 U939 ( .A(n841), .B(KEYINPUT43), .ZN(n843) );
  XNOR2_X1 U940 ( .A(KEYINPUT111), .B(G2678), .ZN(n842) );
  XNOR2_X1 U941 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U942 ( .A(KEYINPUT42), .B(G2090), .Z(n845) );
  XNOR2_X1 U943 ( .A(G2067), .B(G2072), .ZN(n844) );
  XNOR2_X1 U944 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U945 ( .A(n847), .B(n846), .Z(n849) );
  XNOR2_X1 U946 ( .A(KEYINPUT112), .B(G2096), .ZN(n848) );
  XNOR2_X1 U947 ( .A(n849), .B(n848), .ZN(n851) );
  XOR2_X1 U948 ( .A(G2078), .B(G2084), .Z(n850) );
  XNOR2_X1 U949 ( .A(n851), .B(n850), .ZN(G227) );
  XNOR2_X1 U950 ( .A(G1971), .B(n929), .ZN(n853) );
  XNOR2_X1 U951 ( .A(G1986), .B(G1961), .ZN(n852) );
  XNOR2_X1 U952 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U953 ( .A(n854), .B(G2474), .Z(n856) );
  XNOR2_X1 U954 ( .A(G1981), .B(G1966), .ZN(n855) );
  XNOR2_X1 U955 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U956 ( .A(KEYINPUT41), .B(G1976), .Z(n858) );
  XNOR2_X1 U957 ( .A(G1996), .B(G1991), .ZN(n857) );
  XNOR2_X1 U958 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U959 ( .A(n860), .B(n859), .ZN(G229) );
  INV_X1 U960 ( .A(n861), .ZN(G319) );
  NAND2_X1 U961 ( .A1(n892), .A2(G124), .ZN(n862) );
  XNOR2_X1 U962 ( .A(n862), .B(KEYINPUT44), .ZN(n864) );
  NAND2_X1 U963 ( .A1(G112), .A2(n893), .ZN(n863) );
  NAND2_X1 U964 ( .A1(n864), .A2(n863), .ZN(n869) );
  NAND2_X1 U965 ( .A1(n888), .A2(G100), .ZN(n867) );
  NAND2_X1 U966 ( .A1(G136), .A2(n865), .ZN(n866) );
  NAND2_X1 U967 ( .A1(n867), .A2(n866), .ZN(n868) );
  NOR2_X1 U968 ( .A1(n869), .A2(n868), .ZN(G162) );
  XOR2_X1 U969 ( .A(n984), .B(G162), .Z(n872) );
  XNOR2_X1 U970 ( .A(G160), .B(n870), .ZN(n871) );
  XNOR2_X1 U971 ( .A(n872), .B(n871), .ZN(n876) );
  XOR2_X1 U972 ( .A(KEYINPUT116), .B(KEYINPUT114), .Z(n874) );
  XNOR2_X1 U973 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n873) );
  XNOR2_X1 U974 ( .A(n874), .B(n873), .ZN(n875) );
  XOR2_X1 U975 ( .A(n876), .B(n875), .Z(n879) );
  XOR2_X1 U976 ( .A(G164), .B(n877), .Z(n878) );
  XNOR2_X1 U977 ( .A(n879), .B(n878), .ZN(n904) );
  NAND2_X1 U978 ( .A1(n888), .A2(G106), .ZN(n881) );
  NAND2_X1 U979 ( .A1(G142), .A2(n889), .ZN(n880) );
  NAND2_X1 U980 ( .A1(n881), .A2(n880), .ZN(n882) );
  XNOR2_X1 U981 ( .A(n882), .B(KEYINPUT45), .ZN(n887) );
  NAND2_X1 U982 ( .A1(G130), .A2(n892), .ZN(n884) );
  NAND2_X1 U983 ( .A1(G118), .A2(n893), .ZN(n883) );
  NAND2_X1 U984 ( .A1(n884), .A2(n883), .ZN(n885) );
  XNOR2_X1 U985 ( .A(KEYINPUT113), .B(n885), .ZN(n886) );
  NAND2_X1 U986 ( .A1(n887), .A2(n886), .ZN(n900) );
  NAND2_X1 U987 ( .A1(n888), .A2(G103), .ZN(n891) );
  NAND2_X1 U988 ( .A1(G139), .A2(n889), .ZN(n890) );
  NAND2_X1 U989 ( .A1(n891), .A2(n890), .ZN(n898) );
  NAND2_X1 U990 ( .A1(G127), .A2(n892), .ZN(n895) );
  NAND2_X1 U991 ( .A1(G115), .A2(n893), .ZN(n894) );
  NAND2_X1 U992 ( .A1(n895), .A2(n894), .ZN(n896) );
  XOR2_X1 U993 ( .A(KEYINPUT47), .B(n896), .Z(n897) );
  NOR2_X1 U994 ( .A1(n898), .A2(n897), .ZN(n899) );
  XOR2_X1 U995 ( .A(KEYINPUT115), .B(n899), .Z(n995) );
  XNOR2_X1 U996 ( .A(n900), .B(n995), .ZN(n901) );
  XNOR2_X1 U997 ( .A(n902), .B(n901), .ZN(n903) );
  XNOR2_X1 U998 ( .A(n904), .B(n903), .ZN(n905) );
  NOR2_X1 U999 ( .A1(G37), .A2(n905), .ZN(n906) );
  XOR2_X1 U1000 ( .A(KEYINPUT117), .B(n906), .Z(G395) );
  XNOR2_X1 U1001 ( .A(G286), .B(n943), .ZN(n908) );
  XNOR2_X1 U1002 ( .A(n908), .B(n907), .ZN(n910) );
  XOR2_X1 U1003 ( .A(n931), .B(G171), .Z(n909) );
  XNOR2_X1 U1004 ( .A(n910), .B(n909), .ZN(n911) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n911), .ZN(G397) );
  NOR2_X1 U1006 ( .A1(G227), .A2(G229), .ZN(n913) );
  XNOR2_X1 U1007 ( .A(KEYINPUT49), .B(KEYINPUT118), .ZN(n912) );
  XNOR2_X1 U1008 ( .A(n913), .B(n912), .ZN(n924) );
  XOR2_X1 U1009 ( .A(G2451), .B(G2430), .Z(n915) );
  XNOR2_X1 U1010 ( .A(G2438), .B(G2443), .ZN(n914) );
  XNOR2_X1 U1011 ( .A(n915), .B(n914), .ZN(n921) );
  XOR2_X1 U1012 ( .A(G2435), .B(G2454), .Z(n917) );
  XNOR2_X1 U1013 ( .A(G1348), .B(G1341), .ZN(n916) );
  XNOR2_X1 U1014 ( .A(n917), .B(n916), .ZN(n919) );
  XOR2_X1 U1015 ( .A(G2446), .B(G2427), .Z(n918) );
  XNOR2_X1 U1016 ( .A(n919), .B(n918), .ZN(n920) );
  XOR2_X1 U1017 ( .A(n921), .B(n920), .Z(n922) );
  NAND2_X1 U1018 ( .A1(G14), .A2(n922), .ZN(n927) );
  NAND2_X1 U1019 ( .A1(G319), .A2(n927), .ZN(n923) );
  NOR2_X1 U1020 ( .A1(n924), .A2(n923), .ZN(n926) );
  NOR2_X1 U1021 ( .A1(G395), .A2(G397), .ZN(n925) );
  NAND2_X1 U1022 ( .A1(n926), .A2(n925), .ZN(G225) );
  INV_X1 U1023 ( .A(G225), .ZN(G308) );
  INV_X1 U1024 ( .A(G108), .ZN(G238) );
  INV_X1 U1025 ( .A(n927), .ZN(G401) );
  INV_X1 U1026 ( .A(n928), .ZN(G223) );
  XNOR2_X1 U1027 ( .A(n930), .B(n929), .ZN(n933) );
  XOR2_X1 U1028 ( .A(n931), .B(G1348), .Z(n932) );
  NOR2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n948) );
  XOR2_X1 U1030 ( .A(G171), .B(G1961), .Z(n935) );
  XOR2_X1 U1031 ( .A(G166), .B(G1971), .Z(n934) );
  NOR2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(n942) );
  NAND2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1034 ( .A(KEYINPUT121), .B(n938), .Z(n939) );
  NOR2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1036 ( .A1(n942), .A2(n941), .ZN(n946) );
  XNOR2_X1 U1037 ( .A(G1341), .B(n943), .ZN(n944) );
  XNOR2_X1 U1038 ( .A(KEYINPUT122), .B(n944), .ZN(n945) );
  NOR2_X1 U1039 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1040 ( .A1(n948), .A2(n947), .ZN(n953) );
  XOR2_X1 U1041 ( .A(G1966), .B(G168), .Z(n950) );
  NOR2_X1 U1042 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1043 ( .A(KEYINPUT57), .B(n951), .ZN(n952) );
  NOR2_X1 U1044 ( .A1(n953), .A2(n952), .ZN(n955) );
  XOR2_X1 U1045 ( .A(G16), .B(KEYINPUT56), .Z(n954) );
  NOR2_X1 U1046 ( .A1(n955), .A2(n954), .ZN(n983) );
  XNOR2_X1 U1047 ( .A(KEYINPUT123), .B(G1961), .ZN(n956) );
  XNOR2_X1 U1048 ( .A(n956), .B(G5), .ZN(n971) );
  XNOR2_X1 U1049 ( .A(G1966), .B(G21), .ZN(n969) );
  XNOR2_X1 U1050 ( .A(G1348), .B(KEYINPUT59), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(n957), .B(G4), .ZN(n961) );
  XNOR2_X1 U1052 ( .A(G1981), .B(G6), .ZN(n959) );
  XNOR2_X1 U1053 ( .A(G19), .B(G1341), .ZN(n958) );
  NOR2_X1 U1054 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n964) );
  XNOR2_X1 U1056 ( .A(G20), .B(G1956), .ZN(n962) );
  XNOR2_X1 U1057 ( .A(KEYINPUT124), .B(n962), .ZN(n963) );
  NOR2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n967) );
  XNOR2_X1 U1059 ( .A(KEYINPUT125), .B(KEYINPUT126), .ZN(n965) );
  XNOR2_X1 U1060 ( .A(n965), .B(KEYINPUT60), .ZN(n966) );
  XNOR2_X1 U1061 ( .A(n967), .B(n966), .ZN(n968) );
  NOR2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1063 ( .A1(n971), .A2(n970), .ZN(n979) );
  XNOR2_X1 U1064 ( .A(KEYINPUT58), .B(KEYINPUT127), .ZN(n977) );
  XOR2_X1 U1065 ( .A(G1986), .B(G24), .Z(n975) );
  XNOR2_X1 U1066 ( .A(G1976), .B(G23), .ZN(n973) );
  XNOR2_X1 U1067 ( .A(G1971), .B(G22), .ZN(n972) );
  NOR2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n976) );
  XOR2_X1 U1070 ( .A(n977), .B(n976), .Z(n978) );
  NOR2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n980) );
  XOR2_X1 U1072 ( .A(KEYINPUT61), .B(n980), .Z(n981) );
  NOR2_X1 U1073 ( .A1(G16), .A2(n981), .ZN(n982) );
  NOR2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n1010) );
  XNOR2_X1 U1075 ( .A(G160), .B(G2084), .ZN(n987) );
  NOR2_X1 U1076 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n992) );
  XOR2_X1 U1078 ( .A(G2090), .B(G162), .Z(n988) );
  NOR2_X1 U1079 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1080 ( .A(n990), .B(KEYINPUT51), .ZN(n991) );
  NOR2_X1 U1081 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1082 ( .A1(n994), .A2(n993), .ZN(n1000) );
  XOR2_X1 U1083 ( .A(G2072), .B(n995), .Z(n997) );
  XOR2_X1 U1084 ( .A(G164), .B(G2078), .Z(n996) );
  NOR2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n998) );
  XOR2_X1 U1086 ( .A(KEYINPUT50), .B(n998), .Z(n999) );
  NOR2_X1 U1087 ( .A1(n1000), .A2(n999), .ZN(n1002) );
  NAND2_X1 U1088 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NOR2_X1 U1089 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1090 ( .A(KEYINPUT52), .B(n1005), .ZN(n1007) );
  INV_X1 U1091 ( .A(KEYINPUT55), .ZN(n1006) );
  NAND2_X1 U1092 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1093 ( .A1(n1008), .A2(G29), .ZN(n1009) );
  NAND2_X1 U1094 ( .A1(n1010), .A2(n1009), .ZN(n1035) );
  XNOR2_X1 U1095 ( .A(G2067), .B(G26), .ZN(n1012) );
  XNOR2_X1 U1096 ( .A(G33), .B(G2072), .ZN(n1011) );
  NOR2_X1 U1097 ( .A1(n1012), .A2(n1011), .ZN(n1019) );
  XOR2_X1 U1098 ( .A(G32), .B(G1996), .Z(n1013) );
  NAND2_X1 U1099 ( .A1(n1013), .A2(G28), .ZN(n1017) );
  XOR2_X1 U1100 ( .A(G27), .B(n1014), .Z(n1015) );
  XNOR2_X1 U1101 ( .A(KEYINPUT119), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1102 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1103 ( .A1(n1019), .A2(n1018), .ZN(n1022) );
  XOR2_X1 U1104 ( .A(G25), .B(n1020), .Z(n1021) );
  NOR2_X1 U1105 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1106 ( .A(KEYINPUT120), .B(n1023), .Z(n1024) );
  XOR2_X1 U1107 ( .A(KEYINPUT53), .B(n1024), .Z(n1026) );
  XNOR2_X1 U1108 ( .A(G2090), .B(G35), .ZN(n1025) );
  NOR2_X1 U1109 ( .A1(n1026), .A2(n1025), .ZN(n1029) );
  XOR2_X1 U1110 ( .A(G2084), .B(G34), .Z(n1027) );
  XNOR2_X1 U1111 ( .A(KEYINPUT54), .B(n1027), .ZN(n1028) );
  NAND2_X1 U1112 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XOR2_X1 U1113 ( .A(KEYINPUT55), .B(n1030), .Z(n1032) );
  INV_X1 U1114 ( .A(G29), .ZN(n1031) );
  NAND2_X1 U1115 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NAND2_X1 U1116 ( .A1(G11), .A2(n1033), .ZN(n1034) );
  NOR2_X1 U1117 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XOR2_X1 U1118 ( .A(n1036), .B(KEYINPUT62), .Z(G150) );
  INV_X1 U1119 ( .A(G150), .ZN(G311) );
endmodule

