

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U550 ( .A1(n675), .A2(n802), .ZN(n713) );
  BUF_X1 U551 ( .A(n666), .Z(n529) );
  AND2_X2 U552 ( .A1(n519), .A2(G2104), .ZN(n882) );
  XNOR2_X1 U553 ( .A(n686), .B(n685), .ZN(n726) );
  INV_X1 U554 ( .A(KEYINPUT90), .ZN(n684) );
  NOR2_X1 U555 ( .A1(n753), .A2(n735), .ZN(n737) );
  OR2_X1 U556 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U557 ( .A(KEYINPUT29), .B(n711), .Z(n514) );
  NOR2_X1 U558 ( .A1(n742), .A2(n740), .ZN(n515) );
  XOR2_X1 U559 ( .A(KEYINPUT71), .B(n571), .Z(n516) );
  OR2_X1 U560 ( .A1(n697), .A2(n696), .ZN(n705) );
  XNOR2_X1 U561 ( .A(n684), .B(KEYINPUT31), .ZN(n685) );
  NOR2_X1 U562 ( .A1(G1966), .A2(n742), .ZN(n728) );
  AND2_X1 U563 ( .A1(n733), .A2(n732), .ZN(n753) );
  INV_X1 U564 ( .A(KEYINPUT93), .ZN(n736) );
  XOR2_X1 U565 ( .A(KEYINPUT72), .B(n578), .Z(n964) );
  NOR2_X1 U566 ( .A1(n527), .A2(n526), .ZN(G160) );
  INV_X1 U567 ( .A(G2105), .ZN(n519) );
  NOR2_X1 U568 ( .A1(G2104), .A2(n519), .ZN(n878) );
  NAND2_X1 U569 ( .A1(G125), .A2(n878), .ZN(n518) );
  AND2_X1 U570 ( .A1(G2105), .A2(G2104), .ZN(n879) );
  NAND2_X1 U571 ( .A1(G113), .A2(n879), .ZN(n517) );
  NAND2_X1 U572 ( .A1(n518), .A2(n517), .ZN(n527) );
  NAND2_X1 U573 ( .A1(G101), .A2(n882), .ZN(n520) );
  XNOR2_X1 U574 ( .A(n520), .B(KEYINPUT23), .ZN(n521) );
  XNOR2_X1 U575 ( .A(KEYINPUT65), .B(n521), .ZN(n525) );
  NOR2_X1 U576 ( .A1(G2105), .A2(G2104), .ZN(n522) );
  XOR2_X1 U577 ( .A(KEYINPUT17), .B(n522), .Z(n666) );
  NAND2_X1 U578 ( .A1(G137), .A2(n666), .ZN(n523) );
  XNOR2_X1 U579 ( .A(n523), .B(KEYINPUT66), .ZN(n524) );
  NAND2_X1 U580 ( .A1(n525), .A2(n524), .ZN(n526) );
  AND2_X1 U581 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U582 ( .A1(G123), .A2(n878), .ZN(n528) );
  XNOR2_X1 U583 ( .A(n528), .B(KEYINPUT18), .ZN(n536) );
  NAND2_X1 U584 ( .A1(G99), .A2(n882), .ZN(n531) );
  NAND2_X1 U585 ( .A1(G135), .A2(n529), .ZN(n530) );
  NAND2_X1 U586 ( .A1(n531), .A2(n530), .ZN(n534) );
  NAND2_X1 U587 ( .A1(G111), .A2(n879), .ZN(n532) );
  XNOR2_X1 U588 ( .A(KEYINPUT77), .B(n532), .ZN(n533) );
  NOR2_X1 U589 ( .A1(n534), .A2(n533), .ZN(n535) );
  NAND2_X1 U590 ( .A1(n536), .A2(n535), .ZN(n936) );
  XNOR2_X1 U591 ( .A(G2096), .B(n936), .ZN(n537) );
  OR2_X1 U592 ( .A1(G2100), .A2(n537), .ZN(G156) );
  INV_X1 U593 ( .A(G860), .ZN(n589) );
  NOR2_X1 U594 ( .A1(G651), .A2(G543), .ZN(n628) );
  NAND2_X1 U595 ( .A1(n628), .A2(G81), .ZN(n538) );
  XNOR2_X1 U596 ( .A(n538), .B(KEYINPUT12), .ZN(n540) );
  XOR2_X1 U597 ( .A(G543), .B(KEYINPUT0), .Z(n614) );
  INV_X1 U598 ( .A(G651), .ZN(n545) );
  NOR2_X1 U599 ( .A1(n614), .A2(n545), .ZN(n629) );
  NAND2_X1 U600 ( .A1(G68), .A2(n629), .ZN(n539) );
  NAND2_X1 U601 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U602 ( .A(n541), .B(KEYINPUT13), .ZN(n544) );
  NOR2_X1 U603 ( .A1(G651), .A2(n614), .ZN(n542) );
  XNOR2_X2 U604 ( .A(KEYINPUT64), .B(n542), .ZN(n634) );
  NAND2_X1 U605 ( .A1(G43), .A2(n634), .ZN(n543) );
  NAND2_X1 U606 ( .A1(n544), .A2(n543), .ZN(n549) );
  NOR2_X1 U607 ( .A1(G543), .A2(n545), .ZN(n546) );
  XOR2_X2 U608 ( .A(KEYINPUT1), .B(n546), .Z(n632) );
  NAND2_X1 U609 ( .A1(n632), .A2(G56), .ZN(n547) );
  XOR2_X1 U610 ( .A(KEYINPUT14), .B(n547), .Z(n548) );
  NOR2_X1 U611 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U612 ( .A(KEYINPUT70), .B(n550), .Z(n968) );
  OR2_X1 U613 ( .A1(n589), .A2(n968), .ZN(G153) );
  INV_X1 U614 ( .A(G132), .ZN(G219) );
  INV_X1 U615 ( .A(G82), .ZN(G220) );
  INV_X1 U616 ( .A(G57), .ZN(G237) );
  INV_X1 U617 ( .A(G69), .ZN(G235) );
  INV_X1 U618 ( .A(G108), .ZN(G238) );
  INV_X1 U619 ( .A(G120), .ZN(G236) );
  NAND2_X1 U620 ( .A1(n628), .A2(G89), .ZN(n551) );
  XNOR2_X1 U621 ( .A(KEYINPUT4), .B(n551), .ZN(n554) );
  NAND2_X1 U622 ( .A1(n629), .A2(G76), .ZN(n552) );
  XOR2_X1 U623 ( .A(KEYINPUT73), .B(n552), .Z(n553) );
  NAND2_X1 U624 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U625 ( .A(n555), .B(KEYINPUT5), .ZN(n560) );
  NAND2_X1 U626 ( .A1(G63), .A2(n632), .ZN(n557) );
  NAND2_X1 U627 ( .A1(G51), .A2(n634), .ZN(n556) );
  NAND2_X1 U628 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U629 ( .A(KEYINPUT6), .B(n558), .Z(n559) );
  NAND2_X1 U630 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U631 ( .A(n561), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U632 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U633 ( .A1(G7), .A2(G661), .ZN(n562) );
  XNOR2_X1 U634 ( .A(n562), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U635 ( .A(G223), .ZN(n819) );
  NAND2_X1 U636 ( .A1(n819), .A2(G567), .ZN(n563) );
  XOR2_X1 U637 ( .A(KEYINPUT11), .B(n563), .Z(G234) );
  NAND2_X1 U638 ( .A1(G90), .A2(n628), .ZN(n565) );
  NAND2_X1 U639 ( .A1(G77), .A2(n629), .ZN(n564) );
  NAND2_X1 U640 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U641 ( .A(KEYINPUT9), .B(n566), .ZN(n570) );
  NAND2_X1 U642 ( .A1(n634), .A2(G52), .ZN(n568) );
  NAND2_X1 U643 ( .A1(G64), .A2(n632), .ZN(n567) );
  AND2_X1 U644 ( .A1(n568), .A2(n567), .ZN(n569) );
  NAND2_X1 U645 ( .A1(n570), .A2(n569), .ZN(G301) );
  NAND2_X1 U646 ( .A1(G66), .A2(n632), .ZN(n571) );
  NAND2_X1 U647 ( .A1(G79), .A2(n629), .ZN(n572) );
  NAND2_X1 U648 ( .A1(n516), .A2(n572), .ZN(n576) );
  NAND2_X1 U649 ( .A1(n628), .A2(G92), .ZN(n574) );
  NAND2_X1 U650 ( .A1(G54), .A2(n634), .ZN(n573) );
  NAND2_X1 U651 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U652 ( .A(n577), .B(KEYINPUT15), .ZN(n578) );
  NOR2_X1 U653 ( .A1(n964), .A2(G868), .ZN(n580) );
  INV_X1 U654 ( .A(G868), .ZN(n650) );
  NOR2_X1 U655 ( .A1(n650), .A2(G301), .ZN(n579) );
  NOR2_X1 U656 ( .A1(n580), .A2(n579), .ZN(G284) );
  NAND2_X1 U657 ( .A1(G65), .A2(n632), .ZN(n582) );
  NAND2_X1 U658 ( .A1(G53), .A2(n634), .ZN(n581) );
  NAND2_X1 U659 ( .A1(n582), .A2(n581), .ZN(n586) );
  NAND2_X1 U660 ( .A1(G91), .A2(n628), .ZN(n584) );
  NAND2_X1 U661 ( .A1(G78), .A2(n629), .ZN(n583) );
  NAND2_X1 U662 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U663 ( .A1(n586), .A2(n585), .ZN(n967) );
  INV_X1 U664 ( .A(n967), .ZN(G299) );
  NOR2_X1 U665 ( .A1(G286), .A2(n650), .ZN(n588) );
  NOR2_X1 U666 ( .A1(G868), .A2(G299), .ZN(n587) );
  NOR2_X1 U667 ( .A1(n588), .A2(n587), .ZN(G297) );
  NAND2_X1 U668 ( .A1(G559), .A2(n589), .ZN(n590) );
  XNOR2_X1 U669 ( .A(n590), .B(KEYINPUT74), .ZN(n591) );
  INV_X1 U670 ( .A(n964), .ZN(n697) );
  NAND2_X1 U671 ( .A1(n591), .A2(n697), .ZN(n592) );
  XNOR2_X1 U672 ( .A(KEYINPUT16), .B(n592), .ZN(G148) );
  NOR2_X1 U673 ( .A1(n964), .A2(n650), .ZN(n593) );
  XOR2_X1 U674 ( .A(KEYINPUT76), .B(n593), .Z(n594) );
  NOR2_X1 U675 ( .A1(G559), .A2(n594), .ZN(n597) );
  NOR2_X1 U676 ( .A1(n968), .A2(G868), .ZN(n595) );
  XOR2_X1 U677 ( .A(KEYINPUT75), .B(n595), .Z(n596) );
  NOR2_X1 U678 ( .A1(n597), .A2(n596), .ZN(G282) );
  NAND2_X1 U679 ( .A1(n697), .A2(G559), .ZN(n598) );
  XNOR2_X1 U680 ( .A(n598), .B(n968), .ZN(n647) );
  NOR2_X1 U681 ( .A1(n647), .A2(G860), .ZN(n606) );
  NAND2_X1 U682 ( .A1(G67), .A2(n632), .ZN(n600) );
  NAND2_X1 U683 ( .A1(G55), .A2(n634), .ZN(n599) );
  NAND2_X1 U684 ( .A1(n600), .A2(n599), .ZN(n604) );
  NAND2_X1 U685 ( .A1(G93), .A2(n628), .ZN(n602) );
  NAND2_X1 U686 ( .A1(G80), .A2(n629), .ZN(n601) );
  NAND2_X1 U687 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U688 ( .A1(n604), .A2(n603), .ZN(n649) );
  XNOR2_X1 U689 ( .A(n649), .B(KEYINPUT78), .ZN(n605) );
  XNOR2_X1 U690 ( .A(n606), .B(n605), .ZN(G145) );
  NAND2_X1 U691 ( .A1(n628), .A2(G86), .ZN(n608) );
  NAND2_X1 U692 ( .A1(G48), .A2(n634), .ZN(n607) );
  NAND2_X1 U693 ( .A1(n608), .A2(n607), .ZN(n611) );
  NAND2_X1 U694 ( .A1(n629), .A2(G73), .ZN(n609) );
  XOR2_X1 U695 ( .A(KEYINPUT2), .B(n609), .Z(n610) );
  NOR2_X1 U696 ( .A1(n611), .A2(n610), .ZN(n613) );
  NAND2_X1 U697 ( .A1(n632), .A2(G61), .ZN(n612) );
  NAND2_X1 U698 ( .A1(n613), .A2(n612), .ZN(G305) );
  NAND2_X1 U699 ( .A1(n614), .A2(G87), .ZN(n616) );
  NAND2_X1 U700 ( .A1(G49), .A2(n634), .ZN(n615) );
  NAND2_X1 U701 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U702 ( .A1(n632), .A2(n617), .ZN(n620) );
  NAND2_X1 U703 ( .A1(G74), .A2(G651), .ZN(n618) );
  XOR2_X1 U704 ( .A(KEYINPUT79), .B(n618), .Z(n619) );
  NAND2_X1 U705 ( .A1(n620), .A2(n619), .ZN(G288) );
  NAND2_X1 U706 ( .A1(n628), .A2(G88), .ZN(n621) );
  XNOR2_X1 U707 ( .A(n621), .B(KEYINPUT80), .ZN(n623) );
  NAND2_X1 U708 ( .A1(G75), .A2(n629), .ZN(n622) );
  NAND2_X1 U709 ( .A1(n623), .A2(n622), .ZN(n627) );
  NAND2_X1 U710 ( .A1(G62), .A2(n632), .ZN(n625) );
  NAND2_X1 U711 ( .A1(G50), .A2(n634), .ZN(n624) );
  NAND2_X1 U712 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U713 ( .A1(n627), .A2(n626), .ZN(G166) );
  NAND2_X1 U714 ( .A1(G85), .A2(n628), .ZN(n631) );
  NAND2_X1 U715 ( .A1(G72), .A2(n629), .ZN(n630) );
  NAND2_X1 U716 ( .A1(n631), .A2(n630), .ZN(n639) );
  NAND2_X1 U717 ( .A1(n632), .A2(G60), .ZN(n633) );
  XOR2_X1 U718 ( .A(KEYINPUT67), .B(n633), .Z(n636) );
  NAND2_X1 U719 ( .A1(G47), .A2(n634), .ZN(n635) );
  NAND2_X1 U720 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U721 ( .A(KEYINPUT68), .B(n637), .ZN(n638) );
  NOR2_X1 U722 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U723 ( .A(n640), .B(KEYINPUT69), .ZN(G290) );
  XNOR2_X1 U724 ( .A(G288), .B(KEYINPUT19), .ZN(n642) );
  XNOR2_X1 U725 ( .A(n967), .B(G166), .ZN(n641) );
  XNOR2_X1 U726 ( .A(n642), .B(n641), .ZN(n643) );
  XOR2_X1 U727 ( .A(n649), .B(n643), .Z(n644) );
  XNOR2_X1 U728 ( .A(G305), .B(n644), .ZN(n645) );
  XNOR2_X1 U729 ( .A(n645), .B(G290), .ZN(n848) );
  XNOR2_X1 U730 ( .A(KEYINPUT81), .B(n848), .ZN(n646) );
  XNOR2_X1 U731 ( .A(n647), .B(n646), .ZN(n648) );
  NOR2_X1 U732 ( .A1(n650), .A2(n648), .ZN(n652) );
  AND2_X1 U733 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U734 ( .A1(n652), .A2(n651), .ZN(G295) );
  NAND2_X1 U735 ( .A1(G2084), .A2(G2078), .ZN(n653) );
  XOR2_X1 U736 ( .A(KEYINPUT20), .B(n653), .Z(n654) );
  NAND2_X1 U737 ( .A1(G2090), .A2(n654), .ZN(n655) );
  XNOR2_X1 U738 ( .A(KEYINPUT21), .B(n655), .ZN(n656) );
  NAND2_X1 U739 ( .A1(n656), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U740 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U741 ( .A1(G236), .A2(G238), .ZN(n658) );
  NOR2_X1 U742 ( .A1(G235), .A2(G237), .ZN(n657) );
  NAND2_X1 U743 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U744 ( .A(KEYINPUT82), .B(n659), .ZN(n825) );
  NAND2_X1 U745 ( .A1(G567), .A2(n825), .ZN(n664) );
  NOR2_X1 U746 ( .A1(G220), .A2(G219), .ZN(n660) );
  XOR2_X1 U747 ( .A(KEYINPUT22), .B(n660), .Z(n661) );
  NOR2_X1 U748 ( .A1(G218), .A2(n661), .ZN(n662) );
  NAND2_X1 U749 ( .A1(G96), .A2(n662), .ZN(n824) );
  NAND2_X1 U750 ( .A1(G2106), .A2(n824), .ZN(n663) );
  NAND2_X1 U751 ( .A1(n664), .A2(n663), .ZN(n826) );
  NAND2_X1 U752 ( .A1(G661), .A2(G483), .ZN(n665) );
  NOR2_X1 U753 ( .A1(n826), .A2(n665), .ZN(n823) );
  NAND2_X1 U754 ( .A1(n823), .A2(G36), .ZN(G176) );
  NAND2_X1 U755 ( .A1(G102), .A2(n882), .ZN(n668) );
  NAND2_X1 U756 ( .A1(G138), .A2(n666), .ZN(n667) );
  NAND2_X1 U757 ( .A1(n668), .A2(n667), .ZN(n672) );
  NAND2_X1 U758 ( .A1(G126), .A2(n878), .ZN(n670) );
  NAND2_X1 U759 ( .A1(G114), .A2(n879), .ZN(n669) );
  NAND2_X1 U760 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U761 ( .A1(n672), .A2(n671), .ZN(G164) );
  XNOR2_X1 U762 ( .A(KEYINPUT83), .B(G166), .ZN(G303) );
  INV_X1 U763 ( .A(G301), .ZN(G171) );
  NOR2_X1 U764 ( .A1(G1976), .A2(G288), .ZN(n973) );
  INV_X1 U765 ( .A(n973), .ZN(n674) );
  INV_X1 U766 ( .A(KEYINPUT33), .ZN(n673) );
  AND2_X1 U767 ( .A1(n674), .A2(n673), .ZN(n739) );
  NAND2_X1 U768 ( .A1(G160), .A2(G40), .ZN(n801) );
  INV_X1 U769 ( .A(n801), .ZN(n675) );
  NOR2_X1 U770 ( .A1(G164), .A2(G1384), .ZN(n802) );
  NAND2_X1 U771 ( .A1(n713), .A2(G8), .ZN(n676) );
  XNOR2_X1 U772 ( .A(n676), .B(KEYINPUT87), .ZN(n750) );
  INV_X1 U773 ( .A(n750), .ZN(n742) );
  NOR2_X1 U774 ( .A1(G2084), .A2(n713), .ZN(n727) );
  NOR2_X1 U775 ( .A1(n728), .A2(n727), .ZN(n677) );
  NAND2_X1 U776 ( .A1(G8), .A2(n677), .ZN(n678) );
  XNOR2_X1 U777 ( .A(KEYINPUT30), .B(n678), .ZN(n679) );
  NOR2_X1 U778 ( .A1(n679), .A2(G168), .ZN(n683) );
  XOR2_X1 U779 ( .A(G1961), .B(KEYINPUT88), .Z(n989) );
  NAND2_X1 U780 ( .A1(n989), .A2(n713), .ZN(n681) );
  INV_X1 U781 ( .A(n713), .ZN(n699) );
  XNOR2_X1 U782 ( .A(G2078), .B(KEYINPUT25), .ZN(n917) );
  NAND2_X1 U783 ( .A1(n699), .A2(n917), .ZN(n680) );
  NAND2_X1 U784 ( .A1(n681), .A2(n680), .ZN(n687) );
  NOR2_X1 U785 ( .A1(G171), .A2(n687), .ZN(n682) );
  NOR2_X1 U786 ( .A1(n683), .A2(n682), .ZN(n686) );
  NAND2_X1 U787 ( .A1(n687), .A2(G171), .ZN(n712) );
  NAND2_X1 U788 ( .A1(n699), .A2(G2072), .ZN(n688) );
  XNOR2_X1 U789 ( .A(n688), .B(KEYINPUT27), .ZN(n690) );
  INV_X1 U790 ( .A(G1956), .ZN(n990) );
  NOR2_X1 U791 ( .A1(n990), .A2(n699), .ZN(n689) );
  NOR2_X1 U792 ( .A1(n690), .A2(n689), .ZN(n706) );
  NOR2_X1 U793 ( .A1(n967), .A2(n706), .ZN(n691) );
  XOR2_X1 U794 ( .A(n691), .B(KEYINPUT28), .Z(n710) );
  INV_X1 U795 ( .A(G1996), .ZN(n918) );
  NOR2_X1 U796 ( .A1(n713), .A2(n918), .ZN(n692) );
  XOR2_X1 U797 ( .A(n692), .B(KEYINPUT26), .Z(n694) );
  NAND2_X1 U798 ( .A1(n713), .A2(G1341), .ZN(n693) );
  NAND2_X1 U799 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U800 ( .A1(n968), .A2(n695), .ZN(n696) );
  NAND2_X1 U801 ( .A1(n697), .A2(n696), .ZN(n703) );
  AND2_X1 U802 ( .A1(n713), .A2(G1348), .ZN(n698) );
  XNOR2_X1 U803 ( .A(n698), .B(KEYINPUT89), .ZN(n701) );
  NAND2_X1 U804 ( .A1(n699), .A2(G2067), .ZN(n700) );
  NAND2_X1 U805 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U806 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U807 ( .A1(n705), .A2(n704), .ZN(n708) );
  NAND2_X1 U808 ( .A1(n967), .A2(n706), .ZN(n707) );
  NAND2_X1 U809 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U810 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U811 ( .A1(n712), .A2(n514), .ZN(n725) );
  NOR2_X1 U812 ( .A1(G2090), .A2(n713), .ZN(n714) );
  XOR2_X1 U813 ( .A(KEYINPUT91), .B(n714), .Z(n716) );
  NOR2_X1 U814 ( .A1(G1971), .A2(n742), .ZN(n715) );
  NOR2_X1 U815 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U816 ( .A1(n717), .A2(G303), .ZN(n719) );
  AND2_X1 U817 ( .A1(n725), .A2(n719), .ZN(n718) );
  NAND2_X1 U818 ( .A1(n726), .A2(n718), .ZN(n723) );
  INV_X1 U819 ( .A(n719), .ZN(n720) );
  OR2_X1 U820 ( .A1(n720), .A2(G286), .ZN(n721) );
  AND2_X1 U821 ( .A1(G8), .A2(n721), .ZN(n722) );
  NAND2_X1 U822 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U823 ( .A(KEYINPUT32), .B(n724), .ZN(n733) );
  AND2_X1 U824 ( .A1(n726), .A2(n725), .ZN(n731) );
  AND2_X1 U825 ( .A1(G8), .A2(n727), .ZN(n729) );
  OR2_X1 U826 ( .A1(n729), .A2(n728), .ZN(n730) );
  OR2_X1 U827 ( .A1(n731), .A2(n730), .ZN(n732) );
  NOR2_X1 U828 ( .A1(G1971), .A2(G303), .ZN(n734) );
  XNOR2_X1 U829 ( .A(KEYINPUT92), .B(n734), .ZN(n735) );
  XNOR2_X1 U830 ( .A(n737), .B(n736), .ZN(n738) );
  NAND2_X1 U831 ( .A1(n739), .A2(n738), .ZN(n748) );
  NAND2_X1 U832 ( .A1(G1976), .A2(G288), .ZN(n974) );
  INV_X1 U833 ( .A(n974), .ZN(n740) );
  NOR2_X1 U834 ( .A1(KEYINPUT33), .A2(n515), .ZN(n746) );
  XOR2_X1 U835 ( .A(G1981), .B(G305), .Z(n980) );
  NOR2_X1 U836 ( .A1(KEYINPUT33), .A2(KEYINPUT93), .ZN(n741) );
  NOR2_X1 U837 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U838 ( .A1(n973), .A2(n743), .ZN(n744) );
  NAND2_X1 U839 ( .A1(n980), .A2(n744), .ZN(n745) );
  NOR2_X1 U840 ( .A1(n746), .A2(n745), .ZN(n747) );
  AND2_X1 U841 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U842 ( .A(n749), .B(KEYINPUT94), .ZN(n759) );
  NOR2_X1 U843 ( .A1(G2090), .A2(G303), .ZN(n751) );
  NAND2_X1 U844 ( .A1(G8), .A2(n751), .ZN(n752) );
  XOR2_X1 U845 ( .A(KEYINPUT95), .B(n752), .Z(n755) );
  INV_X1 U846 ( .A(n753), .ZN(n754) );
  NAND2_X1 U847 ( .A1(n755), .A2(n754), .ZN(n756) );
  XOR2_X1 U848 ( .A(KEYINPUT96), .B(n756), .Z(n757) );
  NOR2_X1 U849 ( .A1(n750), .A2(n757), .ZN(n758) );
  NOR2_X1 U850 ( .A1(n759), .A2(n758), .ZN(n806) );
  NOR2_X1 U851 ( .A1(G1981), .A2(G305), .ZN(n760) );
  XNOR2_X1 U852 ( .A(n760), .B(KEYINPUT24), .ZN(n761) );
  NAND2_X1 U853 ( .A1(n761), .A2(n750), .ZN(n804) );
  NAND2_X1 U854 ( .A1(G141), .A2(n529), .ZN(n763) );
  NAND2_X1 U855 ( .A1(G129), .A2(n878), .ZN(n762) );
  NAND2_X1 U856 ( .A1(n763), .A2(n762), .ZN(n766) );
  NAND2_X1 U857 ( .A1(n882), .A2(G105), .ZN(n764) );
  XOR2_X1 U858 ( .A(KEYINPUT38), .B(n764), .Z(n765) );
  NOR2_X1 U859 ( .A1(n766), .A2(n765), .ZN(n768) );
  NAND2_X1 U860 ( .A1(n879), .A2(G117), .ZN(n767) );
  NAND2_X1 U861 ( .A1(n768), .A2(n767), .ZN(n875) );
  NOR2_X1 U862 ( .A1(G1996), .A2(n875), .ZN(n769) );
  XOR2_X1 U863 ( .A(KEYINPUT97), .B(n769), .Z(n943) );
  NAND2_X1 U864 ( .A1(G119), .A2(n878), .ZN(n771) );
  NAND2_X1 U865 ( .A1(G107), .A2(n879), .ZN(n770) );
  NAND2_X1 U866 ( .A1(n771), .A2(n770), .ZN(n772) );
  XOR2_X1 U867 ( .A(KEYINPUT86), .B(n772), .Z(n776) );
  NAND2_X1 U868 ( .A1(G95), .A2(n882), .ZN(n774) );
  NAND2_X1 U869 ( .A1(G131), .A2(n529), .ZN(n773) );
  AND2_X1 U870 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U871 ( .A1(n776), .A2(n775), .ZN(n892) );
  NAND2_X1 U872 ( .A1(G1991), .A2(n892), .ZN(n778) );
  NAND2_X1 U873 ( .A1(G1996), .A2(n875), .ZN(n777) );
  NAND2_X1 U874 ( .A1(n778), .A2(n777), .ZN(n809) );
  NOR2_X1 U875 ( .A1(G1991), .A2(n892), .ZN(n938) );
  NOR2_X1 U876 ( .A1(G1986), .A2(G290), .ZN(n779) );
  XNOR2_X1 U877 ( .A(KEYINPUT98), .B(n779), .ZN(n780) );
  NOR2_X1 U878 ( .A1(n938), .A2(n780), .ZN(n781) );
  XOR2_X1 U879 ( .A(KEYINPUT99), .B(n781), .Z(n782) );
  NOR2_X1 U880 ( .A1(n809), .A2(n782), .ZN(n783) );
  NOR2_X1 U881 ( .A1(n943), .A2(n783), .ZN(n784) );
  XNOR2_X1 U882 ( .A(KEYINPUT39), .B(n784), .ZN(n796) );
  XNOR2_X1 U883 ( .A(G2067), .B(KEYINPUT37), .ZN(n785) );
  XOR2_X1 U884 ( .A(n785), .B(KEYINPUT84), .Z(n797) );
  NAND2_X1 U885 ( .A1(n882), .A2(G104), .ZN(n786) );
  XOR2_X1 U886 ( .A(KEYINPUT85), .B(n786), .Z(n788) );
  NAND2_X1 U887 ( .A1(n529), .A2(G140), .ZN(n787) );
  NAND2_X1 U888 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U889 ( .A(KEYINPUT34), .B(n789), .ZN(n794) );
  NAND2_X1 U890 ( .A1(G128), .A2(n878), .ZN(n791) );
  NAND2_X1 U891 ( .A1(G116), .A2(n879), .ZN(n790) );
  NAND2_X1 U892 ( .A1(n791), .A2(n790), .ZN(n792) );
  XOR2_X1 U893 ( .A(KEYINPUT35), .B(n792), .Z(n793) );
  NOR2_X1 U894 ( .A1(n794), .A2(n793), .ZN(n795) );
  XOR2_X1 U895 ( .A(KEYINPUT36), .B(n795), .Z(n862) );
  NAND2_X1 U896 ( .A1(n797), .A2(n862), .ZN(n808) );
  NAND2_X1 U897 ( .A1(n796), .A2(n808), .ZN(n799) );
  NOR2_X1 U898 ( .A1(n862), .A2(n797), .ZN(n798) );
  XOR2_X1 U899 ( .A(KEYINPUT100), .B(n798), .Z(n954) );
  NAND2_X1 U900 ( .A1(n799), .A2(n954), .ZN(n800) );
  XOR2_X1 U901 ( .A(KEYINPUT101), .B(n800), .Z(n803) );
  NOR2_X1 U902 ( .A1(n802), .A2(n801), .ZN(n811) );
  NAND2_X1 U903 ( .A1(n803), .A2(n811), .ZN(n807) );
  AND2_X1 U904 ( .A1(n804), .A2(n807), .ZN(n805) );
  NAND2_X1 U905 ( .A1(n806), .A2(n805), .ZN(n816) );
  INV_X1 U906 ( .A(n807), .ZN(n814) );
  XOR2_X1 U907 ( .A(G1986), .B(G290), .Z(n986) );
  INV_X1 U908 ( .A(n808), .ZN(n810) );
  NOR2_X1 U909 ( .A1(n810), .A2(n809), .ZN(n948) );
  NAND2_X1 U910 ( .A1(n986), .A2(n948), .ZN(n812) );
  NAND2_X1 U911 ( .A1(n812), .A2(n811), .ZN(n813) );
  OR2_X1 U912 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U913 ( .A1(n816), .A2(n815), .ZN(n818) );
  XNOR2_X1 U914 ( .A(KEYINPUT40), .B(KEYINPUT102), .ZN(n817) );
  XNOR2_X1 U915 ( .A(n818), .B(n817), .ZN(G329) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n819), .ZN(G217) );
  AND2_X1 U917 ( .A1(G15), .A2(G2), .ZN(n820) );
  NAND2_X1 U918 ( .A1(G661), .A2(n820), .ZN(G259) );
  NAND2_X1 U919 ( .A1(G3), .A2(G1), .ZN(n821) );
  XOR2_X1 U920 ( .A(KEYINPUT105), .B(n821), .Z(n822) );
  NAND2_X1 U921 ( .A1(n823), .A2(n822), .ZN(G188) );
  XOR2_X1 U922 ( .A(G96), .B(KEYINPUT106), .Z(G221) );
  NOR2_X1 U923 ( .A1(n825), .A2(n824), .ZN(G325) );
  XNOR2_X1 U924 ( .A(KEYINPUT107), .B(G325), .ZN(G261) );
  XOR2_X1 U926 ( .A(KEYINPUT108), .B(n826), .Z(G319) );
  XOR2_X1 U927 ( .A(KEYINPUT42), .B(G2090), .Z(n828) );
  XNOR2_X1 U928 ( .A(G2084), .B(G2078), .ZN(n827) );
  XNOR2_X1 U929 ( .A(n828), .B(n827), .ZN(n829) );
  XOR2_X1 U930 ( .A(n829), .B(G2100), .Z(n831) );
  XNOR2_X1 U931 ( .A(G2067), .B(G2072), .ZN(n830) );
  XNOR2_X1 U932 ( .A(n831), .B(n830), .ZN(n835) );
  XOR2_X1 U933 ( .A(G2096), .B(KEYINPUT43), .Z(n833) );
  XNOR2_X1 U934 ( .A(G2678), .B(KEYINPUT109), .ZN(n832) );
  XNOR2_X1 U935 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U936 ( .A(n835), .B(n834), .Z(G227) );
  XOR2_X1 U937 ( .A(G1976), .B(G1956), .Z(n837) );
  XNOR2_X1 U938 ( .A(G1986), .B(G1961), .ZN(n836) );
  XNOR2_X1 U939 ( .A(n837), .B(n836), .ZN(n847) );
  XOR2_X1 U940 ( .A(KEYINPUT112), .B(G2474), .Z(n839) );
  XNOR2_X1 U941 ( .A(G1996), .B(KEYINPUT110), .ZN(n838) );
  XNOR2_X1 U942 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U943 ( .A(G1981), .B(G1971), .Z(n841) );
  XNOR2_X1 U944 ( .A(G1991), .B(G1966), .ZN(n840) );
  XNOR2_X1 U945 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U946 ( .A(n843), .B(n842), .Z(n845) );
  XNOR2_X1 U947 ( .A(KEYINPUT111), .B(KEYINPUT41), .ZN(n844) );
  XNOR2_X1 U948 ( .A(n845), .B(n844), .ZN(n846) );
  XNOR2_X1 U949 ( .A(n847), .B(n846), .ZN(G229) );
  XOR2_X1 U950 ( .A(n848), .B(G286), .Z(n850) );
  XNOR2_X1 U951 ( .A(n964), .B(G171), .ZN(n849) );
  XNOR2_X1 U952 ( .A(n850), .B(n849), .ZN(n851) );
  XNOR2_X1 U953 ( .A(n851), .B(n968), .ZN(n852) );
  NOR2_X1 U954 ( .A1(G37), .A2(n852), .ZN(G397) );
  NAND2_X1 U955 ( .A1(G124), .A2(n878), .ZN(n853) );
  XNOR2_X1 U956 ( .A(n853), .B(KEYINPUT44), .ZN(n855) );
  NAND2_X1 U957 ( .A1(n882), .A2(G100), .ZN(n854) );
  NAND2_X1 U958 ( .A1(n855), .A2(n854), .ZN(n859) );
  NAND2_X1 U959 ( .A1(G136), .A2(n529), .ZN(n857) );
  NAND2_X1 U960 ( .A1(G112), .A2(n879), .ZN(n856) );
  NAND2_X1 U961 ( .A1(n857), .A2(n856), .ZN(n858) );
  NOR2_X1 U962 ( .A1(n859), .A2(n858), .ZN(G162) );
  XOR2_X1 U963 ( .A(KEYINPUT46), .B(KEYINPUT115), .Z(n861) );
  XNOR2_X1 U964 ( .A(KEYINPUT117), .B(KEYINPUT48), .ZN(n860) );
  XNOR2_X1 U965 ( .A(n861), .B(n860), .ZN(n863) );
  XOR2_X1 U966 ( .A(n863), .B(n862), .Z(n865) );
  XNOR2_X1 U967 ( .A(G164), .B(G160), .ZN(n864) );
  XNOR2_X1 U968 ( .A(n865), .B(n864), .ZN(n866) );
  XNOR2_X1 U969 ( .A(G162), .B(n866), .ZN(n877) );
  NAND2_X1 U970 ( .A1(G127), .A2(n878), .ZN(n868) );
  NAND2_X1 U971 ( .A1(G115), .A2(n879), .ZN(n867) );
  NAND2_X1 U972 ( .A1(n868), .A2(n867), .ZN(n869) );
  XNOR2_X1 U973 ( .A(n869), .B(KEYINPUT47), .ZN(n871) );
  NAND2_X1 U974 ( .A1(G103), .A2(n882), .ZN(n870) );
  NAND2_X1 U975 ( .A1(n871), .A2(n870), .ZN(n874) );
  NAND2_X1 U976 ( .A1(n529), .A2(G139), .ZN(n872) );
  XOR2_X1 U977 ( .A(KEYINPUT116), .B(n872), .Z(n873) );
  NOR2_X1 U978 ( .A1(n874), .A2(n873), .ZN(n949) );
  XNOR2_X1 U979 ( .A(n875), .B(n949), .ZN(n876) );
  XNOR2_X1 U980 ( .A(n877), .B(n876), .ZN(n894) );
  NAND2_X1 U981 ( .A1(G130), .A2(n878), .ZN(n881) );
  NAND2_X1 U982 ( .A1(G118), .A2(n879), .ZN(n880) );
  NAND2_X1 U983 ( .A1(n881), .A2(n880), .ZN(n889) );
  XNOR2_X1 U984 ( .A(KEYINPUT114), .B(KEYINPUT45), .ZN(n887) );
  NAND2_X1 U985 ( .A1(n529), .A2(G142), .ZN(n885) );
  NAND2_X1 U986 ( .A1(n882), .A2(G106), .ZN(n883) );
  XOR2_X1 U987 ( .A(KEYINPUT113), .B(n883), .Z(n884) );
  NAND2_X1 U988 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U989 ( .A(n887), .B(n886), .Z(n888) );
  NOR2_X1 U990 ( .A1(n889), .A2(n888), .ZN(n890) );
  XNOR2_X1 U991 ( .A(n890), .B(n936), .ZN(n891) );
  XNOR2_X1 U992 ( .A(n892), .B(n891), .ZN(n893) );
  XNOR2_X1 U993 ( .A(n894), .B(n893), .ZN(n895) );
  NOR2_X1 U994 ( .A1(G37), .A2(n895), .ZN(n896) );
  XNOR2_X1 U995 ( .A(KEYINPUT118), .B(n896), .ZN(G395) );
  XNOR2_X1 U996 ( .A(G2451), .B(G2446), .ZN(n906) );
  XOR2_X1 U997 ( .A(G2430), .B(KEYINPUT104), .Z(n898) );
  XNOR2_X1 U998 ( .A(G2454), .B(G2435), .ZN(n897) );
  XNOR2_X1 U999 ( .A(n898), .B(n897), .ZN(n902) );
  XOR2_X1 U1000 ( .A(G2438), .B(KEYINPUT103), .Z(n900) );
  XNOR2_X1 U1001 ( .A(G1341), .B(G1348), .ZN(n899) );
  XNOR2_X1 U1002 ( .A(n900), .B(n899), .ZN(n901) );
  XOR2_X1 U1003 ( .A(n902), .B(n901), .Z(n904) );
  XNOR2_X1 U1004 ( .A(G2443), .B(G2427), .ZN(n903) );
  XNOR2_X1 U1005 ( .A(n904), .B(n903), .ZN(n905) );
  XNOR2_X1 U1006 ( .A(n906), .B(n905), .ZN(n907) );
  NAND2_X1 U1007 ( .A1(n907), .A2(G14), .ZN(n913) );
  NAND2_X1 U1008 ( .A1(n913), .A2(G319), .ZN(n910) );
  NOR2_X1 U1009 ( .A1(G227), .A2(G229), .ZN(n908) );
  XNOR2_X1 U1010 ( .A(KEYINPUT49), .B(n908), .ZN(n909) );
  NOR2_X1 U1011 ( .A1(n910), .A2(n909), .ZN(n912) );
  NOR2_X1 U1012 ( .A1(G397), .A2(G395), .ZN(n911) );
  NAND2_X1 U1013 ( .A1(n912), .A2(n911), .ZN(G225) );
  INV_X1 U1014 ( .A(G225), .ZN(G308) );
  INV_X1 U1015 ( .A(n913), .ZN(G401) );
  XNOR2_X1 U1016 ( .A(G29), .B(KEYINPUT123), .ZN(n934) );
  XOR2_X1 U1017 ( .A(KEYINPUT55), .B(KEYINPUT122), .Z(n932) );
  XNOR2_X1 U1018 ( .A(G2090), .B(G35), .ZN(n927) );
  XOR2_X1 U1019 ( .A(G1991), .B(G25), .Z(n914) );
  NAND2_X1 U1020 ( .A1(n914), .A2(G28), .ZN(n924) );
  XNOR2_X1 U1021 ( .A(G2067), .B(G26), .ZN(n916) );
  XNOR2_X1 U1022 ( .A(G33), .B(G2072), .ZN(n915) );
  NOR2_X1 U1023 ( .A1(n916), .A2(n915), .ZN(n922) );
  XOR2_X1 U1024 ( .A(n917), .B(G27), .Z(n920) );
  XOR2_X1 U1025 ( .A(n918), .B(G32), .Z(n919) );
  NOR2_X1 U1026 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1027 ( .A1(n922), .A2(n921), .ZN(n923) );
  NOR2_X1 U1028 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1029 ( .A(KEYINPUT53), .B(n925), .ZN(n926) );
  NOR2_X1 U1030 ( .A1(n927), .A2(n926), .ZN(n930) );
  XOR2_X1 U1031 ( .A(G2084), .B(G34), .Z(n928) );
  XNOR2_X1 U1032 ( .A(KEYINPUT54), .B(n928), .ZN(n929) );
  NAND2_X1 U1033 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1034 ( .A(n932), .B(n931), .ZN(n933) );
  NAND2_X1 U1035 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1036 ( .A1(n935), .A2(G11), .ZN(n963) );
  XNOR2_X1 U1037 ( .A(G160), .B(G2084), .ZN(n937) );
  NAND2_X1 U1038 ( .A1(n937), .A2(n936), .ZN(n939) );
  NOR2_X1 U1039 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1040 ( .A(n940), .B(KEYINPUT119), .ZN(n946) );
  XOR2_X1 U1041 ( .A(G2090), .B(G162), .Z(n941) );
  XNOR2_X1 U1042 ( .A(KEYINPUT120), .B(n941), .ZN(n942) );
  NOR2_X1 U1043 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1044 ( .A(KEYINPUT51), .B(n944), .ZN(n945) );
  NOR2_X1 U1045 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1046 ( .A1(n948), .A2(n947), .ZN(n957) );
  XNOR2_X1 U1047 ( .A(G2072), .B(n949), .ZN(n951) );
  XNOR2_X1 U1048 ( .A(G164), .B(G2078), .ZN(n950) );
  NAND2_X1 U1049 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1050 ( .A(n952), .B(KEYINPUT50), .ZN(n953) );
  XNOR2_X1 U1051 ( .A(n953), .B(KEYINPUT121), .ZN(n955) );
  NAND2_X1 U1052 ( .A1(n955), .A2(n954), .ZN(n956) );
  NOR2_X1 U1053 ( .A1(n957), .A2(n956), .ZN(n958) );
  XOR2_X1 U1054 ( .A(KEYINPUT52), .B(n958), .Z(n959) );
  NOR2_X1 U1055 ( .A1(KEYINPUT55), .A2(n959), .ZN(n961) );
  INV_X1 U1056 ( .A(G29), .ZN(n960) );
  NOR2_X1 U1057 ( .A1(n961), .A2(n960), .ZN(n962) );
  NOR2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n1018) );
  XNOR2_X1 U1059 ( .A(G16), .B(KEYINPUT56), .ZN(n988) );
  XNOR2_X1 U1060 ( .A(G303), .B(G1971), .ZN(n966) );
  XNOR2_X1 U1061 ( .A(n964), .B(G1348), .ZN(n965) );
  NOR2_X1 U1062 ( .A1(n966), .A2(n965), .ZN(n979) );
  XNOR2_X1 U1063 ( .A(n967), .B(G1956), .ZN(n972) );
  XNOR2_X1 U1064 ( .A(G301), .B(G1961), .ZN(n970) );
  XNOR2_X1 U1065 ( .A(n968), .B(G1341), .ZN(n969) );
  NOR2_X1 U1066 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n977) );
  NAND2_X1 U1068 ( .A1(n974), .A2(n674), .ZN(n975) );
  XNOR2_X1 U1069 ( .A(KEYINPUT124), .B(n975), .ZN(n976) );
  NOR2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n984) );
  XNOR2_X1 U1072 ( .A(G1966), .B(G168), .ZN(n981) );
  NAND2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1074 ( .A(KEYINPUT57), .B(n982), .Z(n983) );
  NOR2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1077 ( .A1(n988), .A2(n987), .ZN(n1015) );
  INV_X1 U1078 ( .A(G16), .ZN(n1013) );
  XNOR2_X1 U1079 ( .A(n989), .B(G5), .ZN(n1002) );
  XNOR2_X1 U1080 ( .A(G20), .B(n990), .ZN(n994) );
  XNOR2_X1 U1081 ( .A(G1341), .B(G19), .ZN(n992) );
  XNOR2_X1 U1082 ( .A(G1981), .B(G6), .ZN(n991) );
  NOR2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n997) );
  XOR2_X1 U1085 ( .A(KEYINPUT59), .B(G1348), .Z(n995) );
  XNOR2_X1 U1086 ( .A(G4), .B(n995), .ZN(n996) );
  NOR2_X1 U1087 ( .A1(n997), .A2(n996), .ZN(n998) );
  XOR2_X1 U1088 ( .A(KEYINPUT60), .B(n998), .Z(n1000) );
  XNOR2_X1 U1089 ( .A(G1966), .B(G21), .ZN(n999) );
  NOR2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1010) );
  XNOR2_X1 U1092 ( .A(G1986), .B(G24), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(G22), .B(G1971), .ZN(n1003) );
  NOR2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1007) );
  XNOR2_X1 U1095 ( .A(G1976), .B(KEYINPUT125), .ZN(n1005) );
  XNOR2_X1 U1096 ( .A(n1005), .B(G23), .ZN(n1006) );
  NAND2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1098 ( .A(KEYINPUT58), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1100 ( .A(KEYINPUT61), .B(n1011), .ZN(n1012) );
  NAND2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1103 ( .A(KEYINPUT126), .B(n1016), .Z(n1017) );
  NAND2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1105 ( .A(KEYINPUT62), .B(n1019), .Z(G311) );
  INV_X1 U1106 ( .A(G311), .ZN(G150) );
endmodule

