//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 1 0 0 1 0 0 1 1 0 0 0 0 1 1 1 1 1 0 1 0 0 0 1 0 1 1 0 1 1 0 0 1 1 1 0 1 1 0 0 1 0 1 0 1 1 1 0 1 1 1 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n778, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n864, new_n865, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953;
  INV_X1    g000(.A(KEYINPUT77), .ZN(new_n202));
  NOR2_X1   g001(.A1(G169gat), .A2(G176gat), .ZN(new_n203));
  OAI21_X1  g002(.A(KEYINPUT23), .B1(new_n203), .B2(KEYINPUT67), .ZN(new_n204));
  NAND2_X1  g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT67), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT23), .ZN(new_n207));
  OAI211_X1 g006(.A(new_n206), .B(new_n207), .C1(G169gat), .C2(G176gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n204), .A2(new_n205), .A3(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(G183gat), .B2(G190gat), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  AND2_X1   g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214));
  OR2_X1    g013(.A1(KEYINPUT68), .A2(KEYINPUT24), .ZN(new_n215));
  NAND2_X1  g014(.A1(KEYINPUT68), .A2(KEYINPUT24), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n213), .B1(new_n217), .B2(KEYINPUT69), .ZN(new_n218));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219));
  AND2_X1   g018(.A1(KEYINPUT68), .A2(KEYINPUT24), .ZN(new_n220));
  NOR2_X1   g019(.A1(KEYINPUT68), .A2(KEYINPUT24), .ZN(new_n221));
  OAI211_X1 g020(.A(KEYINPUT69), .B(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n210), .B1(new_n218), .B2(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT24), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n219), .A2(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n225), .B1(new_n227), .B2(KEYINPUT66), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT66), .ZN(new_n230));
  AOI22_X1  g029(.A1(new_n229), .A2(new_n230), .B1(new_n211), .B2(KEYINPUT65), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n228), .B(new_n231), .C1(KEYINPUT65), .C2(new_n211), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n209), .A2(KEYINPUT25), .ZN(new_n233));
  AOI22_X1  g032(.A1(new_n224), .A2(KEYINPUT25), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT70), .ZN(new_n235));
  INV_X1    g034(.A(G183gat), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n235), .B1(new_n236), .B2(KEYINPUT27), .ZN(new_n237));
  AOI21_X1  g036(.A(G190gat), .B1(new_n236), .B2(KEYINPUT27), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT27), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n239), .A2(KEYINPUT70), .A3(G183gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n237), .A2(new_n238), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(KEYINPUT71), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT71), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n237), .A2(new_n238), .A3(new_n243), .A4(new_n240), .ZN(new_n244));
  XNOR2_X1  g043(.A(KEYINPUT72), .B(KEYINPUT28), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n242), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n239), .A2(G183gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n238), .A2(KEYINPUT28), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NOR3_X1   g048(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT73), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n251), .B1(G169gat), .B2(G176gat), .ZN(new_n252));
  OAI21_X1  g051(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n250), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  AND2_X1   g053(.A1(new_n250), .A2(KEYINPUT73), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n219), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n249), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT29), .B1(new_n234), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(G226gat), .A2(G233gat), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n202), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G197gat), .B(G204gat), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT22), .ZN(new_n264));
  INV_X1    g063(.A(G211gat), .ZN(new_n265));
  INV_X1    g064(.A(G218gat), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n263), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(G211gat), .B(G218gat), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n269), .A2(new_n263), .A3(new_n267), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n233), .A2(new_n232), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n212), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n209), .B1(new_n277), .B2(new_n222), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT25), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n274), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n256), .B1(new_n246), .B2(new_n248), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  OAI211_X1 g081(.A(KEYINPUT77), .B(new_n260), .C1(new_n282), .C2(KEYINPUT29), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n234), .A2(new_n258), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n260), .B(KEYINPUT76), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n262), .A2(new_n273), .A3(new_n283), .A4(new_n287), .ZN(new_n288));
  OAI22_X1  g087(.A1(new_n259), .A2(new_n286), .B1(new_n260), .B2(new_n282), .ZN(new_n289));
  INV_X1    g088(.A(new_n273), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(G64gat), .B(G92gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n293), .B(KEYINPUT78), .ZN(new_n294));
  XNOR2_X1  g093(.A(G8gat), .B(G36gat), .ZN(new_n295));
  XOR2_X1   g094(.A(new_n294), .B(new_n295), .Z(new_n296));
  NAND2_X1  g095(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n296), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n288), .A2(new_n291), .A3(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n297), .A2(KEYINPUT30), .A3(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT30), .ZN(new_n301));
  NAND4_X1  g100(.A1(new_n288), .A2(new_n301), .A3(new_n291), .A4(new_n298), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(G225gat), .A2(G233gat), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT80), .ZN(new_n305));
  INV_X1    g104(.A(G155gat), .ZN(new_n306));
  INV_X1    g105(.A(G162gat), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT79), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT79), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n311), .A2(G155gat), .A3(G162gat), .ZN(new_n312));
  OAI21_X1  g111(.A(KEYINPUT80), .B1(G155gat), .B2(G162gat), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n308), .A2(new_n310), .A3(new_n312), .A4(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(G148gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(G141gat), .ZN(new_n316));
  INV_X1    g115(.A(G141gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G148gat), .ZN(new_n318));
  AOI22_X1  g117(.A1(new_n316), .A2(new_n318), .B1(new_n311), .B2(KEYINPUT2), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n314), .A2(new_n319), .ZN(new_n320));
  AND2_X1   g119(.A1(KEYINPUT81), .A2(G141gat), .ZN(new_n321));
  NOR2_X1   g120(.A1(KEYINPUT81), .A2(G141gat), .ZN(new_n322));
  OAI21_X1  g121(.A(G148gat), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT2), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n324), .A2(new_n306), .A3(new_n307), .ZN(new_n325));
  AOI22_X1  g124(.A1(new_n323), .A2(new_n316), .B1(new_n309), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(KEYINPUT3), .B1(new_n320), .B2(new_n326), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n317), .A2(G148gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n315), .A2(G141gat), .ZN(new_n329));
  OAI22_X1  g128(.A1(new_n328), .A2(new_n329), .B1(KEYINPUT79), .B2(new_n324), .ZN(new_n330));
  INV_X1    g129(.A(new_n313), .ZN(new_n331));
  NOR3_X1   g130(.A1(KEYINPUT80), .A2(G155gat), .A3(G162gat), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AND2_X1   g132(.A1(new_n310), .A2(new_n312), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n330), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT3), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n325), .A2(new_n309), .ZN(new_n337));
  OR2_X1    g136(.A1(KEYINPUT81), .A2(G141gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(KEYINPUT81), .A2(G141gat), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n315), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n337), .B1(new_n340), .B2(new_n328), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n335), .A2(new_n336), .A3(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(G120gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(G113gat), .ZN(new_n344));
  INV_X1    g143(.A(G113gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(G120gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT1), .ZN(new_n348));
  INV_X1    g147(.A(G134gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(G127gat), .ZN(new_n350));
  INV_X1    g149(.A(G127gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(G134gat), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n347), .A2(new_n348), .A3(new_n350), .A4(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n350), .A2(new_n352), .ZN(new_n354));
  XNOR2_X1  g153(.A(G113gat), .B(G120gat), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n354), .B1(new_n355), .B2(KEYINPUT1), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n327), .A2(new_n342), .A3(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT4), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n320), .A2(new_n326), .ZN(new_n360));
  INV_X1    g159(.A(new_n357), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(KEYINPUT81), .B(G141gat), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n328), .B1(new_n363), .B2(G148gat), .ZN(new_n364));
  INV_X1    g163(.A(new_n337), .ZN(new_n365));
  OAI22_X1  g164(.A1(new_n364), .A2(new_n365), .B1(new_n314), .B2(new_n319), .ZN(new_n366));
  NOR3_X1   g165(.A1(new_n366), .A2(new_n357), .A3(KEYINPUT4), .ZN(new_n367));
  OAI211_X1 g166(.A(new_n304), .B(new_n358), .C1(new_n362), .C2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT5), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n304), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n360), .A2(new_n361), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n366), .A2(new_n357), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n369), .B1(new_n368), .B2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(G1gat), .B(G29gat), .ZN(new_n377));
  INV_X1    g176(.A(G85gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n377), .B(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(KEYINPUT0), .B(G57gat), .ZN(new_n380));
  XOR2_X1   g179(.A(new_n379), .B(new_n380), .Z(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  NOR3_X1   g181(.A1(new_n371), .A2(new_n376), .A3(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n382), .B1(new_n371), .B2(new_n376), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT6), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n383), .A2(KEYINPUT6), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n303), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT92), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n303), .A2(KEYINPUT92), .A3(new_n389), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(G71gat), .B(G99gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n395), .B(KEYINPUT75), .ZN(new_n396));
  XNOR2_X1  g195(.A(G15gat), .B(G43gat), .ZN(new_n397));
  XOR2_X1   g196(.A(new_n396), .B(new_n397), .Z(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(G227gat), .A2(G233gat), .ZN(new_n400));
  XOR2_X1   g199(.A(new_n400), .B(KEYINPUT64), .Z(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n284), .A2(new_n357), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n282), .A2(new_n361), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n402), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n399), .B1(new_n405), .B2(KEYINPUT33), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n403), .A2(new_n404), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n401), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT74), .B1(new_n409), .B2(KEYINPUT32), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT74), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT32), .ZN(new_n412));
  NOR3_X1   g211(.A1(new_n405), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n407), .B1(new_n410), .B2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT33), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n409), .B(KEYINPUT32), .C1(new_n415), .C2(new_n398), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n403), .A2(new_n404), .A3(new_n402), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n417), .B(KEYINPUT34), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n414), .A2(new_n416), .A3(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n409), .A2(KEYINPUT74), .A3(KEYINPUT32), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n411), .B1(new_n405), .B2(new_n412), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n406), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n416), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n418), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AND3_X1   g224(.A1(new_n420), .A2(new_n425), .A3(KEYINPUT93), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT93), .B1(new_n420), .B2(new_n425), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT35), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT29), .ZN(new_n430));
  INV_X1    g229(.A(new_n272), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n269), .B1(new_n267), .B2(new_n263), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n360), .B1(new_n433), .B2(new_n336), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n273), .B1(new_n342), .B2(new_n430), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT83), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT83), .ZN(new_n437));
  AOI21_X1  g236(.A(KEYINPUT29), .B1(new_n271), .B2(new_n272), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n366), .B1(new_n438), .B2(KEYINPUT3), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT29), .B1(new_n360), .B2(new_n336), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n437), .B(new_n439), .C1(new_n440), .C2(new_n273), .ZN(new_n441));
  NAND2_X1  g240(.A1(G228gat), .A2(G233gat), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n436), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n442), .ZN(new_n444));
  OAI211_X1 g243(.A(KEYINPUT83), .B(new_n444), .C1(new_n434), .C2(new_n435), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(G22gat), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n443), .A2(G22gat), .A3(new_n445), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT85), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(G78gat), .B(G106gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(KEYINPUT31), .B(G50gat), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n446), .A2(KEYINPUT85), .A3(new_n447), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n451), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT84), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n443), .A2(G22gat), .A3(new_n445), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n448), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n454), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n457), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(G22gat), .B1(new_n443), .B2(new_n445), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n457), .B(new_n460), .C1(new_n449), .C2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n456), .B1(new_n461), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT86), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT86), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n467), .B(new_n456), .C1(new_n461), .C2(new_n464), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n394), .A2(new_n428), .A3(new_n429), .A4(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n368), .A2(new_n375), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT5), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n381), .B1(new_n472), .B2(new_n370), .ZN(new_n473));
  OAI21_X1  g272(.A(KEYINPUT82), .B1(new_n473), .B2(KEYINPUT6), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT82), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n385), .A2(new_n475), .A3(new_n386), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n474), .A2(new_n384), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(new_n388), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n303), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n419), .B1(new_n414), .B2(new_n416), .ZN(new_n481));
  NOR3_X1   g280(.A1(new_n423), .A2(new_n424), .A3(new_n418), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n469), .A2(new_n480), .A3(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT94), .ZN(new_n485));
  AND3_X1   g284(.A1(new_n484), .A2(new_n485), .A3(KEYINPUT35), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n485), .B1(new_n484), .B2(KEYINPUT35), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n470), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n466), .A2(new_n479), .A3(new_n468), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT36), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n490), .B1(new_n481), .B2(new_n482), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n420), .A2(new_n425), .A3(KEYINPUT36), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT87), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT91), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT37), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n288), .A2(new_n498), .A3(new_n291), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT89), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n292), .A2(KEYINPUT37), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT89), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n288), .A2(new_n502), .A3(new_n498), .A4(new_n291), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n500), .A2(new_n501), .A3(new_n296), .A4(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n497), .B1(new_n504), .B2(KEYINPUT38), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n387), .A2(new_n388), .A3(new_n299), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n298), .B1(new_n499), .B2(KEYINPUT89), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n498), .B1(new_n289), .B2(new_n273), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n262), .A2(new_n290), .A3(new_n283), .A4(new_n287), .ZN(new_n510));
  AOI21_X1  g309(.A(KEYINPUT38), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n508), .A2(new_n503), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n507), .B1(new_n512), .B2(KEYINPUT90), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT90), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n508), .A2(new_n514), .A3(new_n503), .A4(new_n511), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n504), .A2(new_n497), .A3(KEYINPUT38), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n506), .A2(new_n513), .A3(new_n515), .A4(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT39), .ZN(new_n518));
  NOR3_X1   g317(.A1(new_n373), .A2(new_n374), .A3(new_n372), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n358), .B1(new_n362), .B2(new_n367), .ZN(new_n520));
  AOI211_X1 g319(.A(new_n518), .B(new_n519), .C1(new_n372), .C2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT40), .ZN(new_n522));
  XOR2_X1   g321(.A(KEYINPUT88), .B(KEYINPUT39), .Z(new_n523));
  NAND3_X1  g322(.A1(new_n520), .A2(new_n372), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(new_n382), .ZN(new_n525));
  OR3_X1    g324(.A1(new_n521), .A2(new_n522), .A3(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n522), .B1(new_n521), .B2(new_n525), .ZN(new_n527));
  AND2_X1   g326(.A1(new_n384), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n300), .A2(new_n302), .A3(new_n526), .A4(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n517), .A2(new_n469), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n489), .A2(new_n493), .A3(KEYINPUT87), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n496), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n488), .A2(new_n532), .ZN(new_n533));
  XOR2_X1   g332(.A(G190gat), .B(G218gat), .Z(new_n534));
  INV_X1    g333(.A(KEYINPUT41), .ZN(new_n535));
  NAND2_X1  g334(.A1(G232gat), .A2(G233gat), .ZN(new_n536));
  OAI22_X1  g335(.A1(new_n534), .A2(KEYINPUT102), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(G85gat), .A2(G92gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(KEYINPUT7), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT8), .ZN(new_n540));
  AND2_X1   g339(.A1(G99gat), .A2(G106gat), .ZN(new_n541));
  OAI221_X1 g340(.A(new_n539), .B1(new_n540), .B2(new_n541), .C1(G85gat), .C2(G92gat), .ZN(new_n542));
  NOR2_X1   g341(.A1(G99gat), .A2(G106gat), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT101), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n542), .A2(new_n544), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(G43gat), .B(G50gat), .ZN(new_n551));
  OR3_X1    g350(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n552));
  OAI21_X1  g351(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n553));
  AOI22_X1  g352(.A1(new_n552), .A2(new_n553), .B1(G29gat), .B2(G36gat), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n551), .B1(new_n554), .B2(KEYINPUT15), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(KEYINPUT15), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n555), .B1(new_n556), .B2(new_n551), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n537), .B1(new_n550), .B2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(KEYINPUT17), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(new_n549), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(G134gat), .B(G162gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n534), .A2(KEYINPUT102), .ZN(new_n564));
  XOR2_X1   g363(.A(new_n564), .B(KEYINPUT103), .Z(new_n565));
  NAND2_X1  g364(.A1(new_n536), .A2(new_n535), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n565), .B(new_n566), .Z(new_n567));
  OR2_X1    g366(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n563), .A2(new_n567), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(G57gat), .B(G64gat), .ZN(new_n573));
  XOR2_X1   g372(.A(G71gat), .B(G78gat), .Z(new_n574));
  AOI211_X1 g373(.A(new_n572), .B(new_n573), .C1(new_n574), .C2(KEYINPUT99), .ZN(new_n575));
  OR2_X1    g374(.A1(new_n574), .A2(KEYINPUT99), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  XOR2_X1   g376(.A(G15gat), .B(G22gat), .Z(new_n578));
  INV_X1    g377(.A(G1gat), .ZN(new_n579));
  AND2_X1   g378(.A1(new_n579), .A2(KEYINPUT16), .ZN(new_n580));
  OR2_X1    g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n578), .A2(new_n579), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(G8gat), .B1(new_n582), .B2(KEYINPUT96), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n581), .B(new_n582), .C1(KEYINPUT96), .C2(G8gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n577), .B1(new_n588), .B2(KEYINPUT21), .ZN(new_n589));
  XOR2_X1   g388(.A(G127gat), .B(G155gat), .Z(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G183gat), .B(G211gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT100), .ZN(new_n593));
  NAND2_X1  g392(.A1(G231gat), .A2(G233gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(new_n591), .B(new_n595), .Z(new_n596));
  NOR2_X1   g395(.A1(new_n588), .A2(KEYINPUT21), .ZN(new_n597));
  XOR2_X1   g396(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n596), .B(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n571), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n588), .A2(new_n557), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT98), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n587), .B(KEYINPUT97), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n559), .A2(new_n605), .ZN(new_n606));
  AND2_X1   g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(G229gat), .A2(G233gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT18), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n607), .A2(KEYINPUT18), .A3(new_n608), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n604), .B1(new_n588), .B2(new_n557), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n608), .B(KEYINPUT13), .Z(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n611), .A2(new_n612), .A3(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G113gat), .B(G141gat), .ZN(new_n617));
  INV_X1    g416(.A(G197gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(KEYINPUT11), .B(G169gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(KEYINPUT95), .B(KEYINPUT12), .Z(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n616), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n623), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n611), .A2(new_n625), .A3(new_n612), .A4(new_n615), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT108), .ZN(new_n629));
  AND2_X1   g428(.A1(new_n547), .A2(new_n577), .ZN(new_n630));
  OR2_X1    g429(.A1(new_n544), .A2(KEYINPUT104), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n544), .A2(KEYINPUT104), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n542), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT105), .ZN(new_n634));
  INV_X1    g433(.A(new_n577), .ZN(new_n635));
  AOI22_X1  g434(.A1(new_n630), .A2(new_n634), .B1(new_n549), .B2(new_n635), .ZN(new_n636));
  XOR2_X1   g435(.A(KEYINPUT106), .B(KEYINPUT10), .Z(new_n637));
  AND2_X1   g436(.A1(new_n577), .A2(KEYINPUT10), .ZN(new_n638));
  AOI22_X1  g437(.A1(new_n636), .A2(new_n637), .B1(new_n550), .B2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(G230gat), .ZN(new_n640));
  INV_X1    g439(.A(G233gat), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  NOR3_X1   g442(.A1(new_n636), .A2(new_n640), .A3(new_n641), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n629), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  XOR2_X1   g444(.A(G176gat), .B(G204gat), .Z(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(KEYINPUT107), .ZN(new_n647));
  XNOR2_X1  g446(.A(G120gat), .B(G148gat), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n647), .B(new_n648), .Z(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n645), .A2(new_n650), .ZN(new_n651));
  OAI211_X1 g450(.A(new_n629), .B(new_n649), .C1(new_n643), .C2(new_n644), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NOR3_X1   g453(.A1(new_n602), .A2(new_n628), .A3(new_n654), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n533), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n478), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(G1gat), .ZN(G1324gat));
  INV_X1    g458(.A(new_n303), .ZN(new_n660));
  AND2_X1   g459(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(G8gat), .ZN(new_n662));
  OAI21_X1  g461(.A(KEYINPUT42), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  XOR2_X1   g462(.A(KEYINPUT16), .B(G8gat), .Z(new_n664));
  NAND2_X1  g463(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  MUX2_X1   g464(.A(KEYINPUT42), .B(new_n663), .S(new_n665), .Z(G1325gat));
  AOI21_X1  g465(.A(G15gat), .B1(new_n656), .B2(new_n428), .ZN(new_n667));
  INV_X1    g466(.A(new_n493), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n668), .A2(G15gat), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n667), .B1(new_n656), .B2(new_n669), .ZN(G1326gat));
  INV_X1    g469(.A(new_n468), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n460), .B1(new_n449), .B2(new_n462), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(KEYINPUT84), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(new_n463), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n467), .B1(new_n674), .B2(new_n456), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n656), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(KEYINPUT43), .B(G22gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1327gat));
  NOR3_X1   g478(.A1(new_n654), .A2(new_n628), .A3(new_n601), .ZN(new_n680));
  AOI21_X1  g479(.A(KEYINPUT109), .B1(new_n676), .B2(new_n479), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n466), .A2(new_n479), .A3(KEYINPUT109), .A4(new_n468), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(new_n493), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(KEYINPUT110), .B1(new_n684), .B2(new_n530), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT109), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n489), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n687), .A2(new_n493), .A3(new_n682), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n529), .B1(new_n671), .B2(new_n675), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n513), .A2(new_n515), .ZN(new_n690));
  INV_X1    g489(.A(new_n516), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n691), .A2(new_n505), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n689), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT110), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n688), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n488), .B1(new_n685), .B2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n696), .A2(KEYINPUT111), .A3(new_n697), .A4(new_n570), .ZN(new_n698));
  INV_X1    g497(.A(new_n470), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n484), .A2(KEYINPUT35), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(KEYINPUT94), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n484), .A2(new_n485), .A3(KEYINPUT35), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n699), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n532), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n570), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(KEYINPUT44), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n698), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n694), .B1(new_n688), .B2(new_n693), .ZN(new_n708));
  INV_X1    g507(.A(new_n683), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n709), .A2(new_n530), .A3(KEYINPUT110), .A4(new_n687), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n571), .B1(new_n711), .B2(new_n488), .ZN(new_n712));
  AOI21_X1  g511(.A(KEYINPUT111), .B1(new_n712), .B2(new_n697), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n680), .B1(new_n707), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(G29gat), .B1(new_n714), .B2(new_n478), .ZN(new_n715));
  AND3_X1   g514(.A1(new_n533), .A2(new_n570), .A3(new_n680), .ZN(new_n716));
  INV_X1    g515(.A(G29gat), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n716), .A2(new_n717), .A3(new_n657), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT45), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n715), .A2(new_n719), .ZN(G1328gat));
  INV_X1    g519(.A(KEYINPUT46), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n303), .A2(G36gat), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n716), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT112), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n716), .A2(KEYINPUT112), .A3(new_n722), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n721), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT113), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n725), .A2(new_n721), .A3(new_n726), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(G36gat), .B1(new_n714), .B2(new_n303), .ZN(new_n731));
  OAI211_X1 g530(.A(new_n730), .B(new_n731), .C1(new_n728), .C2(new_n729), .ZN(G1329gat));
  INV_X1    g531(.A(G43gat), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n716), .A2(new_n733), .A3(new_n428), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n734), .A2(KEYINPUT47), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n668), .B(new_n680), .C1(new_n707), .C2(new_n713), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n737), .A2(KEYINPUT114), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT114), .ZN(new_n739));
  OAI21_X1  g538(.A(G43gat), .B1(new_n736), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n735), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n734), .B1(new_n737), .B2(new_n733), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT47), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n741), .A2(new_n744), .ZN(G1330gat));
  XNOR2_X1  g544(.A(KEYINPUT116), .B(KEYINPUT48), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n676), .B(new_n680), .C1(new_n707), .C2(new_n713), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n747), .A2(G50gat), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n469), .A2(G50gat), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n716), .A2(new_n749), .ZN(new_n750));
  OAI211_X1 g549(.A(KEYINPUT115), .B(new_n746), .C1(new_n748), .C2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(new_n746), .ZN(new_n752));
  AOI22_X1  g551(.A1(new_n747), .A2(G50gat), .B1(new_n716), .B2(new_n749), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT115), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n752), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n751), .A2(new_n755), .ZN(G1331gat));
  NOR3_X1   g555(.A1(new_n602), .A2(new_n627), .A3(new_n653), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n696), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n657), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g560(.A1(new_n758), .A2(new_n303), .ZN(new_n762));
  NOR2_X1   g561(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n763));
  AND2_X1   g562(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n762), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n765), .B1(new_n762), .B2(new_n763), .ZN(G1333gat));
  NAND3_X1  g565(.A1(new_n759), .A2(G71gat), .A3(new_n668), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(KEYINPUT117), .ZN(new_n768));
  INV_X1    g567(.A(new_n428), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n758), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(G71gat), .B1(new_n770), .B2(KEYINPUT118), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n771), .B1(KEYINPUT118), .B2(new_n770), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n768), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(KEYINPUT50), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT50), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n768), .A2(new_n775), .A3(new_n772), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n774), .A2(new_n776), .ZN(G1334gat));
  NAND2_X1  g576(.A1(new_n759), .A2(new_n676), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g578(.A1(new_n601), .A2(new_n627), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n696), .A2(new_n570), .A3(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT51), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n712), .A2(KEYINPUT51), .A3(new_n780), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  OR2_X1    g586(.A1(new_n787), .A2(KEYINPUT119), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(KEYINPUT119), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n653), .A2(G85gat), .A3(new_n478), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(KEYINPUT120), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n788), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n707), .A2(new_n713), .ZN(new_n793));
  INV_X1    g592(.A(new_n780), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n793), .A2(new_n653), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n657), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n792), .B1(new_n797), .B2(new_n378), .ZN(G1336gat));
  NOR2_X1   g597(.A1(new_n794), .A2(new_n653), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n799), .B1(new_n707), .B2(new_n713), .ZN(new_n800));
  OAI21_X1  g599(.A(G92gat), .B1(new_n800), .B2(new_n303), .ZN(new_n801));
  OR3_X1    g600(.A1(new_n653), .A2(G92gat), .A3(new_n303), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n801), .B1(new_n787), .B2(new_n802), .ZN(new_n803));
  XNOR2_X1  g602(.A(KEYINPUT121), .B(KEYINPUT52), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n801), .B(new_n804), .C1(new_n787), .C2(new_n802), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(G1337gat));
  NOR3_X1   g607(.A1(new_n769), .A2(G99gat), .A3(new_n653), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n788), .A2(new_n789), .A3(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(G99gat), .B1(new_n800), .B2(new_n493), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(G1338gat));
  NOR3_X1   g611(.A1(new_n653), .A2(new_n469), .A3(G106gat), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n814), .B1(new_n783), .B2(new_n785), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n676), .B(new_n799), .C1(new_n707), .C2(new_n713), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n815), .B1(new_n816), .B2(G106gat), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT122), .ZN(new_n818));
  AND3_X1   g617(.A1(new_n817), .A2(new_n818), .A3(KEYINPUT53), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n818), .A2(KEYINPUT53), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n818), .A2(KEYINPUT53), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n817), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n819), .A2(new_n822), .ZN(G1339gat));
  NOR2_X1   g622(.A1(new_n607), .A2(new_n608), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n613), .A2(new_n614), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n621), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n626), .A2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n570), .B1(new_n654), .B2(new_n828), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n639), .A2(new_n642), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n830), .A2(new_n643), .A3(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n649), .B1(new_n643), .B2(new_n831), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n833), .A2(KEYINPUT55), .A3(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT55), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n643), .A2(new_n831), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n650), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n836), .B1(new_n832), .B2(new_n838), .ZN(new_n839));
  OR3_X1    g638(.A1(new_n643), .A2(new_n644), .A3(new_n650), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n835), .A2(new_n839), .A3(new_n627), .A4(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n601), .B1(new_n829), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n835), .A2(new_n839), .A3(new_n840), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n570), .B1(new_n843), .B2(new_n827), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n602), .A2(new_n654), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n628), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT123), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n848), .A2(new_n849), .A3(new_n469), .ZN(new_n850));
  AOI22_X1  g649(.A1(new_n842), .A2(new_n844), .B1(new_n628), .B2(new_n846), .ZN(new_n851));
  OAI21_X1  g650(.A(KEYINPUT123), .B1(new_n851), .B2(new_n676), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n850), .A2(new_n852), .A3(new_n428), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n657), .A2(new_n303), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(G113gat), .B1(new_n855), .B2(new_n628), .ZN(new_n856));
  INV_X1    g655(.A(new_n483), .ZN(new_n857));
  NOR4_X1   g656(.A1(new_n851), .A2(new_n676), .A3(new_n857), .A4(new_n854), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(new_n345), .A3(new_n627), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n856), .A2(new_n859), .ZN(G1340gat));
  OAI21_X1  g659(.A(G120gat), .B1(new_n855), .B2(new_n653), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n858), .A2(new_n343), .A3(new_n654), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(G1341gat));
  NOR3_X1   g662(.A1(new_n855), .A2(new_n351), .A3(new_n600), .ZN(new_n864));
  AOI21_X1  g663(.A(G127gat), .B1(new_n858), .B2(new_n601), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n864), .A2(new_n865), .ZN(G1342gat));
  NAND3_X1  g665(.A1(new_n858), .A2(new_n349), .A3(new_n570), .ZN(new_n867));
  XOR2_X1   g666(.A(new_n867), .B(KEYINPUT56), .Z(new_n868));
  OAI21_X1  g667(.A(G134gat), .B1(new_n855), .B2(new_n571), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(G1343gat));
  NOR2_X1   g669(.A1(new_n668), .A2(new_n854), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n851), .A2(new_n469), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n873), .A2(KEYINPUT57), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(KEYINPUT57), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n872), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n363), .B1(new_n876), .B2(new_n627), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n873), .A2(new_n871), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n878), .A2(G141gat), .A3(new_n628), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT124), .ZN(new_n881));
  OR2_X1    g680(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(KEYINPUT58), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  OAI211_X1 g683(.A(KEYINPUT58), .B(new_n882), .C1(new_n877), .C2(new_n879), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(G1344gat));
  INV_X1    g685(.A(new_n878), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n887), .A2(new_n315), .A3(new_n654), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n315), .B1(new_n876), .B2(new_n654), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT59), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n889), .A2(new_n890), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n888), .B1(new_n891), .B2(new_n892), .ZN(G1345gat));
  AOI21_X1  g692(.A(G155gat), .B1(new_n887), .B2(new_n601), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n600), .A2(new_n306), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(KEYINPUT125), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n894), .B1(new_n876), .B2(new_n896), .ZN(G1346gat));
  NAND3_X1  g696(.A1(new_n887), .A2(new_n307), .A3(new_n570), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n876), .A2(new_n570), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n898), .B1(new_n899), .B2(new_n307), .ZN(G1347gat));
  NOR2_X1   g699(.A1(new_n657), .A2(new_n303), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n850), .A2(new_n852), .A3(new_n428), .A4(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(G169gat), .B1(new_n902), .B2(new_n628), .ZN(new_n903));
  INV_X1    g702(.A(new_n901), .ZN(new_n904));
  NOR4_X1   g703(.A1(new_n851), .A2(new_n676), .A3(new_n857), .A4(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(G169gat), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n905), .A2(new_n906), .A3(new_n627), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n903), .A2(new_n907), .ZN(G1348gat));
  AOI21_X1  g707(.A(G176gat), .B1(new_n905), .B2(new_n654), .ZN(new_n909));
  INV_X1    g708(.A(new_n902), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n654), .A2(G176gat), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(G1349gat));
  AND3_X1   g711(.A1(new_n850), .A2(new_n852), .A3(new_n428), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n913), .A2(KEYINPUT126), .A3(new_n601), .A4(new_n901), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT126), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n915), .B1(new_n902), .B2(new_n600), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n914), .A2(G183gat), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n236), .A2(KEYINPUT27), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n905), .A2(new_n247), .A3(new_n918), .A4(new_n601), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(KEYINPUT60), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT60), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n917), .A2(new_n922), .A3(new_n919), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n921), .A2(new_n923), .ZN(G1350gat));
  INV_X1    g723(.A(G190gat), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n905), .A2(new_n925), .A3(new_n570), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n570), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT61), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n927), .A2(new_n928), .A3(G190gat), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n928), .B1(new_n927), .B2(G190gat), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n926), .B1(new_n930), .B2(new_n931), .ZN(G1351gat));
  NOR2_X1   g731(.A1(new_n668), .A2(new_n904), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n934), .B1(new_n874), .B2(new_n875), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n618), .B1(new_n935), .B2(new_n627), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n851), .A2(new_n469), .A3(new_n934), .ZN(new_n937));
  AND3_X1   g736(.A1(new_n937), .A2(new_n618), .A3(new_n627), .ZN(new_n938));
  OR2_X1    g737(.A1(new_n936), .A2(new_n938), .ZN(G1352gat));
  INV_X1    g738(.A(G204gat), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n937), .A2(new_n940), .A3(new_n654), .ZN(new_n941));
  XOR2_X1   g740(.A(new_n941), .B(KEYINPUT62), .Z(new_n942));
  NAND3_X1  g741(.A1(new_n935), .A2(KEYINPUT127), .A3(new_n654), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(G204gat), .ZN(new_n944));
  AOI21_X1  g743(.A(KEYINPUT127), .B1(new_n935), .B2(new_n654), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n942), .B1(new_n944), .B2(new_n945), .ZN(G1353gat));
  NAND3_X1  g745(.A1(new_n937), .A2(new_n265), .A3(new_n601), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n935), .A2(new_n601), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n948), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n949));
  AOI21_X1  g748(.A(KEYINPUT63), .B1(new_n948), .B2(G211gat), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n947), .B1(new_n949), .B2(new_n950), .ZN(G1354gat));
  AOI21_X1  g750(.A(G218gat), .B1(new_n937), .B2(new_n570), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n571), .A2(new_n266), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n952), .B1(new_n935), .B2(new_n953), .ZN(G1355gat));
endmodule


