//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 1 0 1 0 0 0 1 0 1 1 1 0 0 0 0 1 0 1 0 1 0 0 0 1 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 0 1 0 1 1 0 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n777, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n865, new_n866, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n986, new_n988,
    new_n989, new_n990, new_n991;
  INV_X1    g000(.A(KEYINPUT97), .ZN(new_n202));
  XOR2_X1   g001(.A(G183gat), .B(G211gat), .Z(new_n203));
  INV_X1    g002(.A(G64gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n204), .A2(G57gat), .ZN(new_n205));
  INV_X1    g004(.A(G57gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n206), .A2(G64gat), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT9), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(G71gat), .A2(G78gat), .ZN(new_n209));
  OR2_X1    g008(.A1(G71gat), .A2(G78gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(KEYINPUT93), .B1(new_n204), .B2(G57gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT93), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n213), .A2(new_n206), .A3(G64gat), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n212), .B(new_n214), .C1(new_n206), .C2(G64gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT9), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n209), .B1(new_n210), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n211), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n219), .B(KEYINPUT94), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT21), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G231gat), .ZN(new_n223));
  INV_X1    g022(.A(G233gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  OAI211_X1 g025(.A(new_n220), .B(new_n221), .C1(new_n223), .C2(new_n224), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(G127gat), .B(G155gat), .ZN(new_n229));
  XOR2_X1   g028(.A(new_n229), .B(KEYINPUT95), .Z(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n228), .A2(new_n230), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n203), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n233), .ZN(new_n235));
  INV_X1    g034(.A(new_n203), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n235), .A2(new_n236), .A3(new_n231), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(G15gat), .B(G22gat), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT16), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n239), .B1(new_n240), .B2(G1gat), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n241), .B1(G1gat), .B2(new_n239), .ZN(new_n242));
  INV_X1    g041(.A(G8gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n242), .B(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n244), .B1(new_n220), .B2(new_n221), .ZN(new_n245));
  XOR2_X1   g044(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n238), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n234), .A2(new_n237), .A3(new_n247), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(G29gat), .ZN(new_n252));
  INV_X1    g051(.A(G36gat), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n252), .A2(new_n253), .A3(KEYINPUT14), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT14), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n255), .B1(G29gat), .B2(G36gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT86), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n257), .A2(new_n258), .B1(G29gat), .B2(G36gat), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n259), .B1(new_n258), .B2(new_n257), .ZN(new_n260));
  XNOR2_X1  g059(.A(G43gat), .B(G50gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT15), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  AND2_X1   g063(.A1(new_n254), .A2(new_n256), .ZN(new_n265));
  OR3_X1    g064(.A1(new_n252), .A2(new_n253), .A3(KEYINPUT88), .ZN(new_n266));
  OAI21_X1  g065(.A(KEYINPUT88), .B1(new_n252), .B2(new_n253), .ZN(new_n267));
  AND4_X1   g066(.A1(new_n262), .A2(new_n265), .A3(new_n266), .A4(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT15), .ZN(new_n269));
  INV_X1    g068(.A(G50gat), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n270), .A2(KEYINPUT87), .A3(G43gat), .ZN(new_n271));
  INV_X1    g070(.A(new_n261), .ZN(new_n272));
  OAI211_X1 g071(.A(new_n269), .B(new_n271), .C1(new_n272), .C2(KEYINPUT87), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n268), .A2(KEYINPUT89), .A3(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(KEYINPUT89), .B1(new_n268), .B2(new_n273), .ZN(new_n276));
  OAI211_X1 g075(.A(KEYINPUT17), .B(new_n264), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(G85gat), .A2(G92gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(KEYINPUT7), .ZN(new_n279));
  INV_X1    g078(.A(G99gat), .ZN(new_n280));
  INV_X1    g079(.A(G106gat), .ZN(new_n281));
  OAI21_X1  g080(.A(KEYINPUT8), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(KEYINPUT96), .B(G92gat), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n279), .B(new_n282), .C1(new_n284), .C2(G85gat), .ZN(new_n285));
  XOR2_X1   g084(.A(G99gat), .B(G106gat), .Z(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  AND2_X1   g086(.A1(new_n266), .A2(new_n267), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n273), .A2(new_n288), .A3(new_n262), .A4(new_n265), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT89), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI22_X1  g090(.A1(new_n291), .A2(new_n274), .B1(new_n263), .B2(new_n260), .ZN(new_n292));
  XNOR2_X1  g091(.A(KEYINPUT90), .B(KEYINPUT17), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n277), .B(new_n287), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n264), .B1(new_n275), .B2(new_n276), .ZN(new_n295));
  INV_X1    g094(.A(new_n286), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n285), .B(new_n296), .ZN(new_n297));
  AND2_X1   g096(.A1(G232gat), .A2(G233gat), .ZN(new_n298));
  AOI22_X1  g097(.A1(new_n295), .A2(new_n297), .B1(KEYINPUT41), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n294), .A2(new_n299), .ZN(new_n300));
  XOR2_X1   g099(.A(G190gat), .B(G218gat), .Z(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n301), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n294), .A2(new_n303), .A3(new_n299), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n298), .A2(KEYINPUT41), .ZN(new_n306));
  XNOR2_X1  g105(.A(G134gat), .B(G162gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n306), .B(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n305), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n302), .A2(new_n308), .A3(new_n304), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n202), .B1(new_n251), .B2(new_n313), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n249), .A2(KEYINPUT97), .A3(new_n250), .A4(new_n312), .ZN(new_n315));
  AND2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n277), .B(new_n244), .C1(new_n292), .C2(new_n293), .ZN(new_n317));
  INV_X1    g116(.A(new_n244), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n295), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(G229gat), .A2(G233gat), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n317), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT91), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT18), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT91), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n317), .A2(new_n319), .A3(new_n324), .A4(new_n320), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n322), .A2(new_n323), .A3(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT92), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n317), .A2(new_n319), .A3(KEYINPUT18), .A4(new_n320), .ZN(new_n329));
  XOR2_X1   g128(.A(new_n320), .B(KEYINPUT13), .Z(new_n330));
  INV_X1    g129(.A(new_n319), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n295), .A2(new_n318), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(G113gat), .B(G141gat), .ZN(new_n334));
  INV_X1    g133(.A(G197gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n334), .B(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(KEYINPUT11), .B(G169gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n336), .B(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n338), .B(KEYINPUT12), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n329), .A2(new_n333), .A3(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n322), .A2(KEYINPUT92), .A3(new_n323), .A4(new_n325), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n328), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n326), .A2(new_n333), .A3(new_n329), .ZN(new_n344));
  INV_X1    g143(.A(new_n339), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n220), .A2(new_n287), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT10), .ZN(new_n349));
  AND2_X1   g148(.A1(new_n286), .A2(KEYINPUT98), .ZN(new_n350));
  OR2_X1    g149(.A1(new_n285), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n285), .A2(new_n350), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n351), .A2(new_n218), .A3(new_n211), .A4(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n348), .A2(new_n349), .A3(new_n353), .ZN(new_n354));
  OR3_X1    g153(.A1(new_n220), .A2(new_n349), .A3(new_n287), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(G230gat), .A2(G233gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n348), .A2(new_n353), .ZN(new_n359));
  INV_X1    g158(.A(new_n357), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(G120gat), .B(G148gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(G176gat), .B(G204gat), .ZN(new_n364));
  XOR2_X1   g163(.A(new_n363), .B(new_n364), .Z(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n358), .A2(new_n361), .A3(new_n365), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  AND3_X1   g169(.A1(new_n316), .A2(new_n347), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(G227gat), .A2(G233gat), .ZN(new_n372));
  INV_X1    g171(.A(G127gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT66), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT66), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(G127gat), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n374), .A2(new_n376), .A3(KEYINPUT67), .A4(G134gat), .ZN(new_n377));
  INV_X1    g176(.A(G113gat), .ZN(new_n378));
  INV_X1    g177(.A(G120gat), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT1), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(G113gat), .A2(G120gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AND2_X1   g181(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n374), .A2(new_n376), .A3(G134gat), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT67), .ZN(new_n385));
  INV_X1    g184(.A(G134gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(G127gat), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n384), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(KEYINPUT68), .B(G120gat), .ZN(new_n389));
  OR2_X1    g188(.A1(new_n389), .A2(new_n378), .ZN(new_n390));
  XNOR2_X1  g189(.A(G127gat), .B(G134gat), .ZN(new_n391));
  AND2_X1   g190(.A1(new_n391), .A2(new_n380), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n383), .A2(new_n388), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  NOR2_X1   g192(.A1(G169gat), .A2(G176gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT23), .ZN(new_n395));
  NAND2_X1  g194(.A1(G169gat), .A2(G176gat), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT23), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n397), .B1(G169gat), .B2(G176gat), .ZN(new_n398));
  AND3_X1   g197(.A1(new_n395), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(G183gat), .ZN(new_n402));
  INV_X1    g201(.A(G190gat), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n401), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n399), .A2(KEYINPUT25), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n395), .A2(new_n396), .A3(new_n398), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n405), .B1(G183gat), .B2(G190gat), .ZN(new_n409));
  NAND2_X1  g208(.A1(G183gat), .A2(G190gat), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT24), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT64), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n400), .A2(KEYINPUT64), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n408), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n407), .B1(new_n415), .B2(KEYINPUT25), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n394), .A2(KEYINPUT26), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT26), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n396), .A2(new_n418), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n417), .B(new_n410), .C1(new_n419), .C2(new_n394), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT27), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(G183gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n402), .A2(KEYINPUT27), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT65), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(G190gat), .B1(new_n423), .B2(KEYINPUT65), .ZN(new_n428));
  AOI21_X1  g227(.A(KEYINPUT28), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT28), .ZN(new_n430));
  NOR3_X1   g229(.A1(new_n425), .A2(new_n430), .A3(G190gat), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n421), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n393), .B1(new_n416), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n416), .A2(new_n432), .A3(new_n393), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n433), .B1(KEYINPUT69), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT69), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n416), .A2(new_n432), .A3(new_n436), .A4(new_n393), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n372), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT32), .ZN(new_n439));
  XNOR2_X1  g238(.A(G15gat), .B(G43gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(G71gat), .B(G99gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n440), .B(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT33), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NOR3_X1   g243(.A1(new_n438), .A2(new_n439), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n434), .A2(KEYINPUT69), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n416), .A2(new_n432), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n380), .B(new_n391), .C1(new_n389), .C2(new_n378), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n377), .A2(new_n382), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n387), .A2(new_n385), .ZN(new_n450));
  XNOR2_X1  g249(.A(KEYINPUT66), .B(G127gat), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n450), .B1(new_n451), .B2(G134gat), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n448), .B1(new_n449), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n447), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n446), .A2(new_n454), .A3(new_n372), .A4(new_n437), .ZN(new_n455));
  XNOR2_X1  g254(.A(new_n455), .B(KEYINPUT34), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n445), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n446), .A2(new_n437), .A3(new_n454), .ZN(new_n458));
  INV_X1    g257(.A(new_n372), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n439), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT33), .B1(new_n458), .B2(new_n459), .ZN(new_n461));
  NOR4_X1   g260(.A1(new_n460), .A2(new_n461), .A3(KEYINPUT70), .A4(new_n442), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT70), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n458), .A2(new_n459), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n442), .B1(new_n464), .B2(new_n443), .ZN(new_n465));
  INV_X1    g264(.A(new_n460), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n457), .B1(new_n462), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n442), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n469), .B1(new_n438), .B2(KEYINPUT33), .ZN(new_n470));
  OAI21_X1  g269(.A(KEYINPUT70), .B1(new_n470), .B2(new_n460), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n465), .A2(new_n463), .A3(new_n466), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n445), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n456), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n468), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT36), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n462), .A2(new_n467), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n456), .B1(new_n477), .B2(new_n445), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT36), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n478), .A2(new_n479), .A3(new_n468), .ZN(new_n480));
  NAND2_X1  g279(.A1(G228gat), .A2(G233gat), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT3), .ZN(new_n482));
  XNOR2_X1  g281(.A(G211gat), .B(G218gat), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(G197gat), .B(G204gat), .ZN(new_n485));
  NAND2_X1  g284(.A1(G211gat), .A2(G218gat), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT71), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT22), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n487), .B1(new_n486), .B2(new_n488), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n484), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT72), .ZN(new_n493));
  INV_X1    g292(.A(new_n491), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n494), .A2(new_n483), .A3(new_n485), .A4(new_n489), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n492), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  OAI211_X1 g295(.A(KEYINPUT72), .B(new_n484), .C1(new_n490), .C2(new_n491), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n482), .B1(new_n498), .B2(KEYINPUT29), .ZN(new_n499));
  OR2_X1    g298(.A1(G141gat), .A2(G148gat), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT2), .ZN(new_n501));
  NAND2_X1  g300(.A1(G141gat), .A2(G148gat), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(G162gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(G155gat), .ZN(new_n505));
  INV_X1    g304(.A(G155gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(G162gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n504), .A2(KEYINPUT74), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT74), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(G162gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n501), .B1(new_n513), .B2(G155gat), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n500), .A2(new_n505), .A3(new_n507), .A4(new_n502), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n509), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n481), .B1(new_n499), .B2(new_n516), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n482), .B(new_n509), .C1(new_n514), .C2(new_n515), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(KEYINPUT75), .ZN(new_n519));
  XNOR2_X1  g318(.A(KEYINPUT74), .B(G162gat), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT2), .B1(new_n520), .B2(new_n506), .ZN(new_n521));
  AND4_X1   g320(.A1(new_n505), .A2(new_n500), .A3(new_n507), .A4(new_n502), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT75), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n523), .A2(new_n524), .A3(new_n482), .A4(new_n509), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT29), .B1(new_n519), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT80), .ZN(new_n527));
  AND2_X1   g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n498), .B1(new_n526), .B2(new_n527), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n517), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(G78gat), .B(G106gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(KEYINPUT31), .B(G50gat), .ZN(new_n532));
  XOR2_X1   g331(.A(new_n531), .B(new_n532), .Z(new_n533));
  NOR2_X1   g332(.A1(new_n533), .A2(KEYINPUT81), .ZN(new_n534));
  AOI21_X1  g333(.A(KEYINPUT29), .B1(new_n492), .B2(new_n495), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n516), .B1(new_n535), .B2(KEYINPUT3), .ZN(new_n536));
  INV_X1    g335(.A(new_n498), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n536), .B1(new_n526), .B2(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n534), .B1(new_n538), .B2(new_n481), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n530), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n533), .A2(KEYINPUT81), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(G22gat), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n530), .A2(new_n539), .A3(new_n542), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(G226gat), .A2(G233gat), .ZN(new_n548));
  XOR2_X1   g347(.A(new_n548), .B(KEYINPUT73), .Z(new_n549));
  INV_X1    g348(.A(KEYINPUT29), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n549), .B1(new_n447), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n549), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n552), .B1(new_n416), .B2(new_n432), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n498), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n414), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n404), .B(new_n405), .C1(new_n400), .C2(KEYINPUT64), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n399), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT25), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n408), .A2(new_n558), .ZN(new_n559));
  AOI22_X1  g358(.A1(new_n557), .A2(new_n558), .B1(new_n406), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n431), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n423), .A2(KEYINPUT65), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(new_n403), .ZN(new_n563));
  AOI21_X1  g362(.A(KEYINPUT65), .B1(new_n423), .B2(new_n424), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n430), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n420), .B1(new_n561), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n550), .B1(new_n560), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(new_n552), .ZN(new_n568));
  INV_X1    g367(.A(new_n553), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n568), .A2(new_n537), .A3(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G8gat), .B(G36gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(G64gat), .B(G92gat), .ZN(new_n572));
  XOR2_X1   g371(.A(new_n571), .B(new_n572), .Z(new_n573));
  NAND3_X1  g372(.A1(new_n554), .A2(new_n570), .A3(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT84), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n568), .A2(new_n576), .A3(new_n537), .A4(new_n569), .ZN(new_n577));
  AND2_X1   g376(.A1(new_n577), .A2(KEYINPUT37), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n554), .A2(new_n570), .A3(KEYINPUT84), .ZN(new_n579));
  AOI21_X1  g378(.A(KEYINPUT38), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n554), .A2(new_n570), .ZN(new_n581));
  INV_X1    g380(.A(new_n573), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(KEYINPUT37), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n575), .B1(new_n580), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n519), .A2(new_n525), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n388), .A2(new_n377), .A3(new_n382), .ZN(new_n588));
  AOI22_X1  g387(.A1(KEYINPUT3), .A2(new_n516), .B1(new_n588), .B2(new_n448), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(KEYINPUT4), .B1(new_n453), .B2(new_n516), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT76), .ZN(new_n592));
  AOI22_X1  g391(.A1(new_n521), .A2(new_n522), .B1(new_n508), .B2(new_n503), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT4), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n593), .A2(new_n588), .A3(new_n594), .A4(new_n448), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n591), .A2(new_n592), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(G225gat), .A2(G233gat), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n593), .A2(new_n588), .A3(new_n448), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n598), .A2(KEYINPUT76), .A3(KEYINPUT4), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n590), .A2(new_n596), .A3(new_n597), .A4(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n453), .A2(new_n516), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n597), .B1(new_n601), .B2(new_n598), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT5), .ZN(new_n603));
  OAI21_X1  g402(.A(KEYINPUT77), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n597), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n453), .A2(new_n516), .ZN(new_n606));
  AOI22_X1  g405(.A1(new_n588), .A2(new_n448), .B1(new_n523), .B2(new_n509), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT77), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n608), .A2(new_n609), .A3(KEYINPUT5), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n600), .A2(new_n604), .A3(new_n610), .ZN(new_n611));
  AOI22_X1  g410(.A1(new_n587), .A2(new_n589), .B1(new_n591), .B2(new_n595), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n605), .A2(KEYINPUT5), .ZN(new_n613));
  AOI21_X1  g412(.A(KEYINPUT79), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n591), .A2(new_n595), .ZN(new_n615));
  AND4_X1   g414(.A1(KEYINPUT79), .A2(new_n590), .A3(new_n615), .A4(new_n613), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n611), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(G1gat), .B(G29gat), .Z(new_n618));
  XNOR2_X1  g417(.A(G57gat), .B(G85gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n617), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT6), .ZN(new_n624));
  INV_X1    g423(.A(new_n622), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n611), .B(new_n625), .C1(new_n614), .C2(new_n616), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n623), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n617), .A2(KEYINPUT6), .A3(new_n622), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n581), .A2(KEYINPUT37), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n582), .B1(new_n581), .B2(KEYINPUT37), .ZN(new_n630));
  OAI21_X1  g429(.A(KEYINPUT38), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n586), .A2(new_n627), .A3(new_n628), .A4(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT83), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n597), .B1(new_n590), .B2(new_n615), .ZN(new_n634));
  XNOR2_X1  g433(.A(KEYINPUT82), .B(KEYINPUT39), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n622), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n601), .A2(new_n598), .A3(new_n597), .ZN(new_n637));
  OAI211_X1 g436(.A(KEYINPUT39), .B(new_n637), .C1(new_n612), .C2(new_n597), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n633), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT40), .ZN(new_n640));
  OR2_X1    g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI22_X1  g440(.A1(new_n639), .A2(new_n640), .B1(new_n617), .B2(new_n622), .ZN(new_n642));
  OR3_X1    g441(.A1(new_n581), .A2(KEYINPUT30), .A3(new_n582), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n583), .A2(KEYINPUT30), .A3(new_n574), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n641), .A2(new_n642), .A3(new_n643), .A4(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n547), .B1(new_n632), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n627), .A2(new_n628), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n644), .A2(new_n643), .ZN(new_n648));
  AND3_X1   g447(.A1(new_n647), .A2(new_n648), .A3(new_n547), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n476), .B(new_n480), .C1(new_n646), .C2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n471), .A2(new_n472), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n547), .B1(new_n651), .B2(new_n457), .ZN(new_n652));
  AOI22_X1  g451(.A1(new_n627), .A2(new_n628), .B1(new_n643), .B2(new_n644), .ZN(new_n653));
  XNOR2_X1  g452(.A(KEYINPUT85), .B(KEYINPUT35), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n478), .A2(new_n652), .A3(new_n653), .A4(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT35), .ZN(new_n656));
  OAI211_X1 g455(.A(new_n468), .B(new_n546), .C1(new_n473), .C2(new_n474), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n647), .A2(new_n648), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n650), .A2(new_n655), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n371), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n647), .ZN(new_n662));
  AND2_X1   g461(.A1(new_n662), .A2(KEYINPUT99), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(KEYINPUT99), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n661), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT100), .B(G1gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(G1324gat));
  NOR2_X1   g468(.A1(new_n661), .A2(new_n648), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(KEYINPUT101), .B(KEYINPUT16), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(G8gat), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  OR2_X1    g473(.A1(new_n674), .A2(KEYINPUT42), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(KEYINPUT42), .ZN(new_n676));
  AOI21_X1  g475(.A(KEYINPUT102), .B1(new_n671), .B2(G8gat), .ZN(new_n677));
  AND3_X1   g476(.A1(new_n671), .A2(KEYINPUT102), .A3(G8gat), .ZN(new_n678));
  OAI211_X1 g477(.A(new_n675), .B(new_n676), .C1(new_n677), .C2(new_n678), .ZN(G1325gat));
  NAND2_X1  g478(.A1(new_n476), .A2(new_n480), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(G15gat), .B1(new_n661), .B2(new_n681), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n475), .A2(G15gat), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n682), .B1(new_n661), .B2(new_n683), .ZN(G1326gat));
  NOR2_X1   g483(.A1(new_n661), .A2(new_n546), .ZN(new_n685));
  XOR2_X1   g484(.A(KEYINPUT43), .B(G22gat), .Z(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(G1327gat));
  AND2_X1   g486(.A1(new_n659), .A2(new_n655), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n312), .B1(new_n688), .B2(new_n650), .ZN(new_n689));
  INV_X1    g488(.A(new_n347), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n251), .A2(new_n370), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n694), .A2(new_n252), .A3(new_n665), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT45), .ZN(new_n696));
  AND3_X1   g495(.A1(new_n310), .A2(KEYINPUT104), .A3(new_n311), .ZN(new_n697));
  AOI21_X1  g496(.A(KEYINPUT104), .B1(new_n310), .B2(new_n311), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n700), .A2(KEYINPUT44), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n660), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n702), .B1(new_n689), .B2(new_n703), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n692), .B(KEYINPUT103), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(new_n665), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(G29gat), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n696), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT105), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n696), .A2(KEYINPUT105), .A3(new_n708), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(G1328gat));
  NOR3_X1   g512(.A1(new_n693), .A2(G36gat), .A3(new_n648), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT46), .ZN(new_n715));
  INV_X1    g514(.A(new_n648), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n706), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n715), .B1(new_n718), .B2(new_n253), .ZN(G1329gat));
  NOR3_X1   g518(.A1(new_n693), .A2(G43gat), .A3(new_n475), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n706), .A2(new_n680), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n720), .B1(new_n721), .B2(G43gat), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g522(.A(KEYINPUT108), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT106), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n703), .B1(new_n660), .B2(new_n313), .ZN(new_n726));
  INV_X1    g525(.A(new_n701), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n727), .B1(new_n688), .B2(new_n650), .ZN(new_n728));
  OAI211_X1 g527(.A(new_n547), .B(new_n705), .C1(new_n726), .C2(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n725), .B1(new_n729), .B2(G50gat), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n729), .A2(new_n725), .A3(G50gat), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n546), .A2(G50gat), .ZN(new_n733));
  AOI21_X1  g532(.A(KEYINPUT48), .B1(new_n694), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n731), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n694), .A2(new_n733), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n704), .A2(KEYINPUT107), .A3(new_n547), .A4(new_n705), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n738), .A2(G50gat), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT107), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n729), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n737), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT48), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n724), .B(new_n735), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n741), .A2(G50gat), .A3(new_n738), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n743), .B1(new_n745), .B2(new_n736), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n732), .A2(new_n734), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n747), .A2(new_n730), .ZN(new_n748));
  OAI21_X1  g547(.A(KEYINPUT108), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n744), .A2(new_n749), .ZN(G1331gat));
  AND4_X1   g549(.A1(new_n690), .A2(new_n314), .A3(new_n315), .A4(new_n369), .ZN(new_n751));
  AND3_X1   g550(.A1(new_n660), .A2(new_n751), .A3(KEYINPUT109), .ZN(new_n752));
  AOI21_X1  g551(.A(KEYINPUT109), .B1(new_n660), .B2(new_n751), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  OR2_X1    g553(.A1(new_n665), .A2(KEYINPUT110), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n665), .A2(KEYINPUT110), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(G57gat), .ZN(G1332gat));
  INV_X1    g558(.A(KEYINPUT111), .ZN(new_n760));
  INV_X1    g559(.A(new_n754), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n761), .A2(new_n648), .ZN(new_n762));
  NOR2_X1   g561(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n763));
  OR2_X1    g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AND2_X1   g563(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n754), .B(new_n716), .C1(new_n763), .C2(new_n765), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n760), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n766), .B(new_n760), .C1(new_n762), .C2(new_n763), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n767), .A2(new_n769), .ZN(G1333gat));
  NOR3_X1   g569(.A1(new_n761), .A2(G71gat), .A3(new_n475), .ZN(new_n771));
  INV_X1    g570(.A(G71gat), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n772), .B1(new_n754), .B2(new_n680), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g573(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n774), .B(new_n775), .ZN(G1334gat));
  NAND2_X1  g575(.A1(new_n754), .A2(new_n547), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(G78gat), .ZN(G1335gat));
  NAND3_X1  g577(.A1(new_n689), .A2(new_n690), .A3(new_n251), .ZN(new_n779));
  XOR2_X1   g578(.A(new_n779), .B(KEYINPUT51), .Z(new_n780));
  NOR3_X1   g579(.A1(new_n666), .A2(G85gat), .A3(new_n370), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n251), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n783), .A2(new_n347), .A3(new_n370), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n704), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n665), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(G85gat), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n782), .A2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT113), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n782), .A2(KEYINPUT113), .A3(new_n787), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(G1336gat));
  NOR3_X1   g591(.A1(new_n370), .A2(G92gat), .A3(new_n648), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n780), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n785), .A2(new_n716), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n284), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(KEYINPUT52), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n794), .A2(new_n799), .A3(new_n796), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n800), .ZN(G1337gat));
  INV_X1    g600(.A(new_n475), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n780), .A2(new_n280), .A3(new_n802), .A4(new_n369), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n785), .A2(new_n680), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n803), .B1(new_n805), .B2(new_n280), .ZN(G1338gat));
  NOR3_X1   g605(.A1(new_n370), .A2(G106gat), .A3(new_n546), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n780), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n785), .A2(new_n547), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(G106gat), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(KEYINPUT53), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT53), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n808), .A2(new_n810), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(G1339gat));
  AND4_X1   g614(.A1(new_n690), .A2(new_n314), .A3(new_n315), .A4(new_n370), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n354), .A2(new_n355), .A3(new_n360), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n358), .A2(KEYINPUT54), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n360), .B1(new_n354), .B2(new_n355), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT54), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n365), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n819), .A2(KEYINPUT55), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(new_n368), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n825));
  AND3_X1   g624(.A1(new_n354), .A2(new_n355), .A3(new_n360), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n826), .A2(new_n820), .A3(new_n821), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n356), .A2(new_n821), .A3(new_n357), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n366), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n825), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT114), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT55), .B1(new_n819), .B2(new_n822), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(KEYINPUT114), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n824), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n340), .B1(new_n326), .B2(new_n327), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n332), .A2(new_n331), .A3(new_n330), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n320), .B1(new_n317), .B2(new_n319), .ZN(new_n838));
  OR2_X1    g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AOI22_X1  g638(.A1(new_n836), .A2(new_n342), .B1(new_n338), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n835), .A2(new_n699), .A3(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n835), .A2(new_n347), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n839), .A2(new_n338), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n343), .A2(new_n369), .A3(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT115), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n840), .A2(KEYINPUT115), .A3(new_n369), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n843), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n842), .B1(new_n849), .B2(new_n700), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n817), .B1(new_n850), .B2(new_n783), .ZN(new_n851));
  INV_X1    g650(.A(new_n657), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n854), .A2(new_n648), .A3(new_n757), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n855), .A2(KEYINPUT116), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n855), .A2(KEYINPUT116), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n378), .B(new_n347), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n851), .A2(new_n648), .A3(new_n852), .A4(new_n665), .ZN(new_n859));
  OAI21_X1  g658(.A(G113gat), .B1(new_n859), .B2(new_n690), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n858), .A2(new_n860), .ZN(G1340gat));
  OAI211_X1 g660(.A(new_n389), .B(new_n369), .C1(new_n856), .C2(new_n857), .ZN(new_n862));
  OAI21_X1  g661(.A(G120gat), .B1(new_n859), .B2(new_n370), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(G1341gat));
  NAND2_X1  g663(.A1(new_n783), .A2(new_n451), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n859), .A2(new_n251), .ZN(new_n866));
  OAI22_X1  g665(.A1(new_n855), .A2(new_n865), .B1(new_n866), .B2(new_n451), .ZN(G1342gat));
  OR2_X1    g666(.A1(new_n859), .A2(new_n312), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n313), .A2(new_n648), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n869), .A2(G134gat), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n854), .A2(new_n757), .A3(new_n870), .ZN(new_n871));
  AOI22_X1  g670(.A1(new_n868), .A2(G134gat), .B1(new_n871), .B2(KEYINPUT56), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n871), .A2(KEYINPUT56), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT117), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n871), .A2(KEYINPUT117), .A3(KEYINPUT56), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n872), .B1(new_n875), .B2(new_n876), .ZN(G1343gat));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n851), .A2(new_n878), .A3(new_n547), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT119), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n830), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n833), .A2(KEYINPUT119), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n824), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AOI22_X1  g682(.A1(new_n883), .A2(new_n347), .B1(new_n840), .B2(new_n369), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n841), .B1(new_n884), .B2(new_n313), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n816), .B1(new_n885), .B2(new_n251), .ZN(new_n886));
  OAI21_X1  g685(.A(KEYINPUT57), .B1(new_n886), .B2(new_n546), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n681), .A2(new_n665), .A3(new_n648), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT118), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n888), .B(new_n889), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n879), .A2(new_n887), .A3(new_n347), .A4(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(G141gat), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n680), .B1(new_n755), .B2(new_n756), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n851), .A2(new_n648), .A3(new_n547), .A4(new_n893), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n690), .A2(G141gat), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  OR3_X1    g695(.A1(new_n894), .A2(KEYINPUT120), .A3(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(KEYINPUT120), .B1(new_n894), .B2(new_n896), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n892), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(KEYINPUT58), .ZN(new_n900));
  INV_X1    g699(.A(new_n894), .ZN(new_n901));
  AOI21_X1  g700(.A(KEYINPUT58), .B1(new_n901), .B2(new_n895), .ZN(new_n902));
  AND3_X1   g701(.A1(new_n892), .A2(new_n902), .A3(KEYINPUT121), .ZN(new_n903));
  AOI21_X1  g702(.A(KEYINPUT121), .B1(new_n892), .B2(new_n902), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n900), .B1(new_n903), .B2(new_n904), .ZN(G1344gat));
  INV_X1    g704(.A(G148gat), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n901), .A2(new_n906), .A3(new_n369), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT59), .ZN(new_n908));
  OR2_X1    g707(.A1(new_n884), .A2(new_n313), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n835), .A2(new_n313), .A3(new_n840), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n783), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n878), .B(new_n547), .C1(new_n911), .C2(new_n816), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n878), .B1(new_n851), .B2(new_n547), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n915), .A2(new_n369), .A3(new_n890), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n908), .B1(new_n916), .B2(G148gat), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n879), .A2(new_n887), .A3(new_n890), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n918), .A2(new_n370), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n919), .A2(KEYINPUT59), .A3(new_n906), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n907), .B1(new_n917), .B2(new_n920), .ZN(G1345gat));
  OAI21_X1  g720(.A(G155gat), .B1(new_n918), .B2(new_n251), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n901), .A2(new_n506), .A3(new_n783), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(G1346gat));
  OAI21_X1  g723(.A(new_n513), .B1(new_n918), .B2(new_n700), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n851), .A2(new_n547), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n869), .A2(new_n513), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n926), .A2(new_n893), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n925), .A2(new_n928), .ZN(G1347gat));
  AND2_X1   g728(.A1(new_n851), .A2(new_n666), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n657), .A2(new_n648), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(G169gat), .B1(new_n932), .B2(new_n347), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n853), .A2(new_n648), .A3(new_n757), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n347), .A2(G169gat), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(G1348gat));
  INV_X1    g735(.A(G176gat), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n932), .A2(new_n937), .A3(new_n369), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n757), .A2(new_n648), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n854), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g739(.A(G176gat), .B1(new_n940), .B2(new_n370), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n938), .A2(new_n941), .ZN(G1349gat));
  INV_X1    g741(.A(new_n425), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n932), .A2(new_n943), .A3(new_n783), .ZN(new_n944));
  OAI21_X1  g743(.A(G183gat), .B1(new_n940), .B2(new_n251), .ZN(new_n945));
  XNOR2_X1  g744(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n946));
  AND3_X1   g745(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n946), .B1(new_n944), .B2(new_n945), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n947), .A2(new_n948), .ZN(G1350gat));
  AOI21_X1  g748(.A(new_n403), .B1(new_n934), .B2(new_n313), .ZN(new_n950));
  XNOR2_X1  g749(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  OR2_X1    g751(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NAND4_X1  g752(.A1(new_n930), .A2(new_n403), .A3(new_n699), .A4(new_n931), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n954), .B(KEYINPUT123), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n950), .A2(new_n952), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n953), .A2(new_n955), .A3(new_n956), .ZN(G1351gat));
  NAND2_X1  g756(.A1(new_n939), .A2(new_n681), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n912), .B1(new_n926), .B2(new_n878), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n958), .B1(new_n959), .B2(KEYINPUT125), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT125), .ZN(new_n961));
  OAI211_X1 g760(.A(new_n912), .B(new_n961), .C1(new_n926), .C2(new_n878), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n690), .A2(new_n335), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n960), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n680), .A2(new_n648), .A3(new_n546), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n930), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n335), .B1(new_n966), .B2(new_n690), .ZN(new_n967));
  AND2_X1   g766(.A1(new_n964), .A2(new_n967), .ZN(G1352gat));
  XNOR2_X1  g767(.A(KEYINPUT126), .B(G204gat), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n370), .A2(new_n969), .ZN(new_n970));
  NAND4_X1  g769(.A1(new_n851), .A2(new_n666), .A3(new_n965), .A4(new_n970), .ZN(new_n971));
  OR2_X1    g770(.A1(new_n971), .A2(KEYINPUT127), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(KEYINPUT127), .ZN(new_n973));
  AND3_X1   g772(.A1(new_n972), .A2(KEYINPUT62), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g773(.A(KEYINPUT62), .B1(new_n972), .B2(new_n973), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g775(.A(KEYINPUT125), .B1(new_n913), .B2(new_n914), .ZN(new_n977));
  INV_X1    g776(.A(new_n958), .ZN(new_n978));
  NAND4_X1  g777(.A1(new_n977), .A2(new_n962), .A3(new_n369), .A4(new_n978), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(new_n969), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n976), .A2(new_n980), .ZN(G1353gat));
  OR3_X1    g780(.A1(new_n966), .A2(G211gat), .A3(new_n251), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n958), .A2(new_n251), .ZN(new_n983));
  OAI211_X1 g782(.A(new_n983), .B(new_n912), .C1(new_n878), .C2(new_n926), .ZN(new_n984));
  AND3_X1   g783(.A1(new_n984), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n985));
  AOI21_X1  g784(.A(KEYINPUT63), .B1(new_n984), .B2(G211gat), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n982), .B1(new_n985), .B2(new_n986), .ZN(G1354gat));
  INV_X1    g786(.A(G218gat), .ZN(new_n988));
  NOR2_X1   g787(.A1(new_n312), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n960), .A2(new_n962), .A3(new_n989), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n988), .B1(new_n966), .B2(new_n700), .ZN(new_n991));
  AND2_X1   g790(.A1(new_n990), .A2(new_n991), .ZN(G1355gat));
endmodule


