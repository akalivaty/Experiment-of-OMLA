//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 0 0 0 0 0 0 1 1 0 0 1 1 1 1 1 1 1 0 0 1 1 1 0 0 1 0 1 0 0 0 0 1 0 0 1 0 0 1 0 0 1 0 0 0 0 1 0 0 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:14 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  OR2_X1    g005(.A1(KEYINPUT0), .A2(G128), .ZN(new_n192));
  NAND2_X1  g006(.A1(KEYINPUT0), .A2(G128), .ZN(new_n193));
  AOI22_X1  g007(.A1(new_n189), .A2(new_n191), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  AND3_X1   g008(.A1(new_n189), .A2(new_n191), .A3(new_n193), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G134), .ZN(new_n197));
  OAI21_X1  g011(.A(KEYINPUT64), .B1(new_n197), .B2(G137), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(KEYINPUT11), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(G137), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT11), .ZN(new_n201));
  OAI211_X1 g015(.A(KEYINPUT64), .B(new_n201), .C1(new_n197), .C2(G137), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n199), .A2(new_n200), .A3(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G131), .ZN(new_n204));
  INV_X1    g018(.A(G131), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n199), .A2(new_n205), .A3(new_n200), .A4(new_n202), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n196), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT1), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n189), .A2(new_n191), .A3(new_n208), .A4(G128), .ZN(new_n209));
  INV_X1    g023(.A(G128), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n210), .B1(new_n189), .B2(KEYINPUT1), .ZN(new_n211));
  XNOR2_X1  g025(.A(G143), .B(G146), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n209), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n197), .A2(G137), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT65), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT65), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n200), .A2(new_n216), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n215), .B(G131), .C1(new_n217), .C2(new_n214), .ZN(new_n218));
  AND3_X1   g032(.A1(new_n213), .A2(new_n206), .A3(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n207), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT30), .ZN(new_n221));
  INV_X1    g035(.A(G116), .ZN(new_n222));
  INV_X1    g036(.A(G119), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(KEYINPUT66), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G119), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n222), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n223), .A2(G116), .ZN(new_n228));
  OAI21_X1  g042(.A(KEYINPUT67), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g043(.A(KEYINPUT2), .B(G113), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT67), .ZN(new_n231));
  INV_X1    g045(.A(new_n228), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT66), .B(G119), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n231), .B(new_n232), .C1(new_n233), .C2(new_n222), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n229), .A2(new_n230), .A3(new_n234), .ZN(new_n235));
  OR3_X1    g049(.A1(new_n227), .A2(new_n230), .A3(new_n228), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT30), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n238), .B1(new_n207), .B2(new_n219), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n221), .A2(new_n237), .A3(new_n239), .ZN(new_n240));
  AND2_X1   g054(.A1(new_n235), .A2(new_n236), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n204), .A2(new_n206), .ZN(new_n242));
  INV_X1    g056(.A(new_n196), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n219), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n241), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n240), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G953), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT68), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G953), .ZN(new_n252));
  AOI21_X1  g066(.A(G237), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G210), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT27), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n254), .B(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT26), .ZN(new_n257));
  OR2_X1    g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n257), .ZN(new_n259));
  AND3_X1   g073(.A1(new_n258), .A2(new_n259), .A3(G101), .ZN(new_n260));
  AOI21_X1  g074(.A(G101), .B1(new_n258), .B2(new_n259), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n248), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT28), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n237), .B1(new_n207), .B2(new_n219), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n264), .B1(new_n246), .B2(new_n265), .ZN(new_n266));
  NOR3_X1   g080(.A1(new_n237), .A2(new_n207), .A3(new_n219), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n267), .A2(KEYINPUT28), .ZN(new_n268));
  OAI21_X1  g082(.A(KEYINPUT69), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n246), .A2(new_n264), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT69), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n262), .B1(new_n269), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n263), .B1(new_n273), .B2(KEYINPUT31), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n256), .B(KEYINPUT26), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n275), .B(G101), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n276), .A2(new_n247), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT31), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n274), .A2(new_n279), .ZN(new_n280));
  NOR2_X1   g094(.A1(G472), .A2(G902), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n281), .B(KEYINPUT70), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT71), .B1(new_n280), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT71), .ZN(new_n285));
  AOI211_X1 g099(.A(new_n285), .B(new_n282), .C1(new_n274), .C2(new_n279), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n187), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n269), .A2(new_n262), .A3(new_n272), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n288), .B1(KEYINPUT72), .B2(KEYINPUT29), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n276), .A2(new_n247), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n289), .B(new_n290), .C1(KEYINPUT72), .C2(new_n288), .ZN(new_n291));
  INV_X1    g105(.A(G902), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT29), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n291), .B(new_n292), .C1(new_n293), .C2(new_n288), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G472), .ZN(new_n295));
  INV_X1    g109(.A(new_n265), .ZN(new_n296));
  OAI21_X1  g110(.A(KEYINPUT28), .B1(new_n296), .B2(new_n267), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n271), .B1(new_n297), .B2(new_n270), .ZN(new_n298));
  INV_X1    g112(.A(new_n272), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n276), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n277), .B1(new_n300), .B2(new_n278), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n263), .A2(KEYINPUT31), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n283), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n303), .A2(new_n187), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n287), .A2(new_n295), .A3(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(G217), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n307), .B1(G234), .B2(new_n292), .ZN(new_n308));
  XOR2_X1   g122(.A(KEYINPUT24), .B(G110), .Z(new_n309));
  NOR2_X1   g123(.A1(new_n233), .A2(new_n210), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n223), .A2(G128), .ZN(new_n311));
  NOR3_X1   g125(.A1(new_n310), .A2(KEYINPUT73), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT73), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n224), .A2(new_n226), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G128), .ZN(new_n315));
  INV_X1    g129(.A(new_n311), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n313), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n309), .B1(new_n312), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT74), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI211_X1 g134(.A(KEYINPUT74), .B(new_n309), .C1(new_n312), .C2(new_n317), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G140), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G125), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n324), .A2(KEYINPUT16), .ZN(new_n325));
  XNOR2_X1  g139(.A(G125), .B(G140), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n325), .B1(new_n326), .B2(KEYINPUT16), .ZN(new_n327));
  OR2_X1    g141(.A1(new_n327), .A2(G146), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(G146), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT75), .B1(new_n314), .B2(G128), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT75), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n233), .A2(new_n332), .A3(new_n210), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT23), .ZN(new_n334));
  OAI211_X1 g148(.A(new_n331), .B(new_n333), .C1(new_n334), .C2(new_n310), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n311), .A2(KEYINPUT23), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AND3_X1   g151(.A1(new_n337), .A2(KEYINPUT76), .A3(G110), .ZN(new_n338));
  AOI21_X1  g152(.A(KEYINPUT76), .B1(new_n337), .B2(G110), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n322), .B(new_n330), .C1(new_n338), .C2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(G110), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n335), .A2(new_n341), .A3(new_n336), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(KEYINPUT77), .ZN(new_n343));
  OR3_X1    g157(.A1(new_n312), .A2(new_n317), .A3(new_n309), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT77), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n335), .A2(new_n345), .A3(new_n341), .A4(new_n336), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n343), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n326), .A2(new_n188), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n347), .A2(new_n329), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n250), .A2(new_n252), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n350), .A2(G221), .A3(G234), .ZN(new_n351));
  XOR2_X1   g165(.A(new_n351), .B(KEYINPUT22), .Z(new_n352));
  XOR2_X1   g166(.A(new_n352), .B(G137), .Z(new_n353));
  NAND3_X1  g167(.A1(new_n340), .A2(new_n349), .A3(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n353), .B1(new_n340), .B2(new_n349), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(KEYINPUT25), .B1(new_n357), .B2(new_n292), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n340), .A2(new_n349), .ZN(new_n359));
  INV_X1    g173(.A(new_n353), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(new_n292), .A3(new_n354), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT25), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n308), .B1(new_n358), .B2(new_n364), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n308), .A2(G902), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n357), .A2(new_n366), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n306), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(G210), .B1(G237), .B2(G902), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n229), .A2(new_n234), .ZN(new_n371));
  XNOR2_X1  g185(.A(KEYINPUT83), .B(KEYINPUT5), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n314), .A2(G116), .ZN(new_n374));
  OAI21_X1  g188(.A(G113), .B1(new_n374), .B2(new_n372), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G104), .ZN(new_n378));
  OAI21_X1  g192(.A(KEYINPUT3), .B1(new_n378), .B2(G107), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT3), .ZN(new_n380));
  INV_X1    g194(.A(G107), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n381), .A3(G104), .ZN(new_n382));
  INV_X1    g196(.A(G101), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n378), .A2(G107), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n379), .A2(new_n382), .A3(new_n383), .A4(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n378), .A2(G107), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n381), .A2(G104), .ZN(new_n387));
  OAI21_X1  g201(.A(G101), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n377), .A2(KEYINPUT84), .A3(new_n236), .A4(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n372), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n392), .B1(new_n229), .B2(new_n234), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n236), .B(new_n390), .C1(new_n393), .C2(new_n375), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT84), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n379), .A2(new_n382), .A3(new_n384), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G101), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n398), .A2(KEYINPUT4), .A3(new_n385), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT4), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n397), .A2(new_n400), .A3(G101), .ZN(new_n401));
  AND2_X1   g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT82), .ZN(new_n403));
  AND3_X1   g217(.A1(new_n402), .A2(new_n237), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n403), .B1(new_n402), .B2(new_n237), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n391), .B(new_n396), .C1(new_n404), .C2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT6), .ZN(new_n407));
  XOR2_X1   g221(.A(G110), .B(G122), .Z(new_n408));
  NAND3_X1  g222(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT85), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n406), .A2(new_n408), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n399), .A2(new_n401), .ZN(new_n412));
  OAI21_X1  g226(.A(KEYINPUT82), .B1(new_n241), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n402), .A2(new_n237), .A3(new_n403), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n408), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n415), .A2(new_n416), .A3(new_n391), .A4(new_n396), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n411), .A2(KEYINPUT6), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n410), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(G125), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n213), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n421), .B1(new_n420), .B2(new_n196), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n249), .A2(G224), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n422), .B(new_n423), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n411), .A2(new_n417), .A3(KEYINPUT85), .A4(KEYINPUT6), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n419), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n377), .A2(new_n236), .A3(new_n389), .ZN(new_n427));
  XOR2_X1   g241(.A(new_n408), .B(KEYINPUT8), .Z(new_n428));
  NAND3_X1  g242(.A1(new_n374), .A2(KEYINPUT5), .A3(new_n232), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n376), .A2(new_n429), .ZN(new_n430));
  AND2_X1   g244(.A1(new_n430), .A2(new_n236), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n427), .B(new_n428), .C1(new_n389), .C2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n423), .A2(KEYINPUT7), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n422), .B(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n417), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  AND2_X1   g249(.A1(new_n435), .A2(new_n292), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n370), .B1(new_n426), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n426), .A2(new_n370), .A3(new_n436), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n438), .A2(KEYINPUT86), .A3(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(G237), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n350), .A2(G214), .A3(new_n441), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n442), .A2(new_n190), .ZN(new_n443));
  AOI21_X1  g257(.A(G143), .B1(new_n253), .B2(G214), .ZN(new_n444));
  OAI21_X1  g258(.A(G131), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT17), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n442), .A2(new_n190), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n253), .A2(G143), .A3(G214), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n447), .A2(new_n205), .A3(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n445), .A2(new_n446), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n205), .B1(new_n447), .B2(new_n448), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(KEYINPUT17), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n450), .A2(new_n328), .A3(new_n329), .A4(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(G113), .B(G122), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n454), .B(new_n378), .ZN(new_n455));
  OAI211_X1 g269(.A(KEYINPUT18), .B(G131), .C1(new_n443), .C2(new_n444), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n420), .A2(G140), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n324), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(G146), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n459), .A2(new_n348), .A3(KEYINPUT87), .ZN(new_n460));
  NAND2_X1  g274(.A1(KEYINPUT18), .A2(G131), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n447), .A2(new_n448), .A3(new_n461), .ZN(new_n462));
  OR3_X1    g276(.A1(new_n326), .A2(KEYINPUT87), .A3(new_n188), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n456), .A2(new_n460), .A3(new_n462), .A4(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n453), .A2(new_n455), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n458), .A2(KEYINPUT19), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT19), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n326), .A2(new_n467), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n469), .A2(KEYINPUT88), .A3(new_n188), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n466), .A2(new_n468), .A3(new_n188), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT88), .ZN(new_n472));
  AOI22_X1  g286(.A1(new_n471), .A2(new_n472), .B1(new_n327), .B2(G146), .ZN(new_n473));
  NOR3_X1   g287(.A1(new_n443), .A2(new_n444), .A3(G131), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n470), .B(new_n473), .C1(new_n474), .C2(new_n451), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n464), .ZN(new_n476));
  INV_X1    g290(.A(new_n455), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI211_X1 g292(.A(G475), .B(G902), .C1(new_n465), .C2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT20), .ZN(new_n480));
  OAI21_X1  g294(.A(KEYINPUT89), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n465), .A2(new_n478), .ZN(new_n482));
  INV_X1    g296(.A(G475), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(new_n483), .A3(new_n292), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT89), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(new_n485), .A3(KEYINPUT20), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n479), .A2(new_n480), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n481), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n455), .B1(new_n453), .B2(new_n464), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT90), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT90), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n465), .A2(new_n491), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n490), .B(new_n292), .C1(new_n492), .C2(new_n489), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(G475), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n488), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(G128), .B(G143), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n496), .B(new_n197), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT13), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n498), .B(G134), .C1(new_n190), .C2(G128), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  XOR2_X1   g314(.A(KEYINPUT91), .B(G107), .Z(new_n501));
  XNOR2_X1  g315(.A(G116), .B(G122), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n501), .B(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n499), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(new_n496), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n500), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  OR2_X1    g320(.A1(new_n222), .A2(G122), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n381), .B1(new_n507), .B2(KEYINPUT14), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(new_n502), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n497), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  XOR2_X1   g325(.A(KEYINPUT9), .B(G234), .Z(new_n512));
  NAND3_X1  g326(.A1(new_n512), .A2(G217), .A3(new_n249), .ZN(new_n513));
  XOR2_X1   g327(.A(new_n513), .B(KEYINPUT92), .Z(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n514), .A2(new_n506), .A3(new_n510), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(KEYINPUT93), .A3(new_n292), .ZN(new_n519));
  INV_X1    g333(.A(G478), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n520), .A2(KEYINPUT15), .ZN(new_n521));
  XOR2_X1   g335(.A(new_n519), .B(new_n521), .Z(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(G952), .ZN(new_n524));
  OR2_X1    g338(.A1(new_n524), .A2(KEYINPUT94), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(KEYINPUT94), .ZN(new_n526));
  AOI21_X1  g340(.A(G953), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n528), .B1(G234), .B2(G237), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  AOI211_X1 g344(.A(new_n292), .B(new_n350), .C1(G234), .C2(G237), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  XOR2_X1   g346(.A(KEYINPUT21), .B(G898), .Z(new_n533));
  OAI21_X1  g347(.A(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  XOR2_X1   g348(.A(new_n534), .B(KEYINPUT95), .Z(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NOR3_X1   g350(.A1(new_n495), .A2(new_n523), .A3(new_n536), .ZN(new_n537));
  OR2_X1    g351(.A1(new_n439), .A2(KEYINPUT86), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n512), .A2(new_n292), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n539), .A2(G221), .ZN(new_n540));
  OAI21_X1  g354(.A(G214), .B1(G237), .B2(G902), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT81), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT80), .ZN(new_n544));
  INV_X1    g358(.A(new_n209), .ZN(new_n545));
  OAI21_X1  g359(.A(KEYINPUT1), .B1(new_n190), .B2(G146), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT79), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n189), .A2(KEYINPUT79), .A3(KEYINPUT1), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n548), .A2(G128), .A3(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n212), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n545), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n544), .B1(new_n552), .B2(new_n389), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n210), .B1(new_n546), .B2(new_n547), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n212), .B1(new_n554), .B2(new_n549), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n390), .B(KEYINPUT80), .C1(new_n555), .C2(new_n545), .ZN(new_n556));
  AOI21_X1  g370(.A(KEYINPUT10), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n243), .A2(new_n399), .A3(new_n401), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n390), .A2(KEYINPUT10), .A3(new_n213), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NOR3_X1   g374(.A1(new_n557), .A2(new_n242), .A3(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(G110), .B(G140), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n562), .B(KEYINPUT78), .ZN(new_n563));
  AND2_X1   g377(.A1(new_n350), .A2(G227), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n563), .B(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n543), .B1(new_n561), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n553), .A2(new_n556), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT10), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n242), .ZN(new_n570));
  INV_X1    g384(.A(new_n560), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n565), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n572), .A2(KEYINPUT81), .A3(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n213), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n389), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n567), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n577), .A2(KEYINPUT12), .A3(new_n242), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT12), .ZN(new_n579));
  AOI22_X1  g393(.A1(new_n553), .A2(new_n556), .B1(new_n575), .B2(new_n389), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n579), .B1(new_n580), .B2(new_n570), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n566), .A2(new_n574), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n570), .B1(new_n569), .B2(new_n571), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n565), .B1(new_n584), .B2(new_n561), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(G469), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n586), .A2(new_n587), .A3(new_n292), .ZN(new_n588));
  AOI21_X1  g402(.A(KEYINPUT12), .B1(new_n577), .B2(new_n242), .ZN(new_n589));
  NOR3_X1   g403(.A1(new_n580), .A2(new_n579), .A3(new_n570), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n572), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n584), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n561), .A2(new_n565), .ZN(new_n593));
  AOI22_X1  g407(.A1(new_n591), .A2(new_n565), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(G469), .B1(new_n594), .B2(G902), .ZN(new_n595));
  AOI211_X1 g409(.A(new_n540), .B(new_n542), .C1(new_n588), .C2(new_n595), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n440), .A2(new_n537), .A3(new_n538), .A4(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n369), .A2(new_n597), .ZN(new_n598));
  XOR2_X1   g412(.A(KEYINPUT96), .B(G101), .Z(new_n599));
  XNOR2_X1  g413(.A(new_n598), .B(new_n599), .ZN(G3));
  NAND2_X1  g414(.A1(new_n303), .A2(new_n285), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n282), .B1(new_n274), .B2(new_n279), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(KEYINPUT71), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n540), .B1(new_n588), .B2(new_n595), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n292), .B1(new_n301), .B2(new_n302), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(G472), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n604), .A2(new_n368), .A3(new_n605), .A4(new_n607), .ZN(new_n608));
  AOI22_X1  g422(.A1(new_n518), .A2(new_n292), .B1(KEYINPUT97), .B2(new_n520), .ZN(new_n609));
  OR2_X1    g423(.A1(new_n520), .A2(KEYINPUT97), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT33), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n518), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n516), .A2(KEYINPUT33), .A3(new_n517), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n613), .A2(new_n614), .A3(G478), .A4(new_n292), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(KEYINPUT98), .ZN(new_n617));
  AOI21_X1  g431(.A(KEYINPUT99), .B1(new_n495), .B2(new_n617), .ZN(new_n618));
  AND3_X1   g432(.A1(new_n495), .A2(KEYINPUT99), .A3(new_n617), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n536), .A2(new_n542), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n426), .A2(new_n370), .A3(new_n436), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n620), .B1(new_n621), .B2(new_n437), .ZN(new_n622));
  NOR4_X1   g436(.A1(new_n608), .A2(new_n618), .A3(new_n619), .A4(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(KEYINPUT34), .B(G104), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G6));
  NAND2_X1  g439(.A1(new_n523), .A2(new_n494), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n479), .A2(KEYINPUT89), .A3(new_n480), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n485), .B1(new_n484), .B2(KEYINPUT20), .ZN(new_n628));
  OAI21_X1  g442(.A(KEYINPUT100), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT100), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n481), .A2(new_n630), .A3(new_n486), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n626), .B1(new_n632), .B2(new_n487), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n438), .A2(new_n439), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n633), .A2(new_n634), .A3(new_n620), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n636), .A2(new_n608), .ZN(new_n637));
  XNOR2_X1  g451(.A(KEYINPUT35), .B(G107), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G9));
  NOR2_X1   g453(.A1(new_n360), .A2(KEYINPUT36), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(new_n359), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n366), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n365), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n604), .A2(new_n607), .A3(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT101), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n646), .A2(new_n597), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(KEYINPUT37), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G110), .ZN(G12));
  OAI211_X1 g463(.A(new_n541), .B(new_n605), .C1(new_n621), .C2(new_n437), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n306), .A2(new_n643), .A3(new_n651), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n627), .A2(new_n628), .A3(KEYINPUT100), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n630), .B1(new_n481), .B2(new_n486), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n487), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n626), .ZN(new_n656));
  INV_X1    g470(.A(G900), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n531), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n530), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n655), .A2(new_n656), .A3(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT102), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n633), .A2(KEYINPUT102), .A3(new_n659), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n652), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(new_n210), .ZN(G30));
  NAND2_X1  g480(.A1(new_n440), .A2(new_n538), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT38), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n659), .B(KEYINPUT39), .Z(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n605), .A2(new_n670), .ZN(new_n671));
  AND2_X1   g485(.A1(new_n671), .A2(KEYINPUT40), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n248), .A2(new_n276), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n246), .A2(new_n265), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n292), .B1(new_n262), .B2(new_n674), .ZN(new_n675));
  OAI21_X1  g489(.A(G472), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n287), .A2(new_n305), .A3(new_n676), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n522), .B1(new_n488), .B2(new_n494), .ZN(new_n678));
  OAI211_X1 g492(.A(new_n677), .B(new_n678), .C1(KEYINPUT40), .C2(new_n671), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n668), .A2(new_n672), .A3(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n357), .A2(KEYINPUT25), .A3(new_n292), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n362), .A2(new_n363), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AOI22_X1  g497(.A1(new_n683), .A2(new_n308), .B1(new_n366), .B2(new_n641), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n680), .A2(new_n541), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(KEYINPUT103), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G143), .ZN(G45));
  AND3_X1   g501(.A1(new_n495), .A2(new_n617), .A3(new_n659), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n306), .A2(new_n643), .A3(new_n651), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G146), .ZN(G48));
  NOR3_X1   g504(.A1(new_n622), .A2(new_n619), .A3(new_n618), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n586), .A2(new_n292), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(G469), .ZN(new_n693));
  INV_X1    g507(.A(new_n540), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n693), .A2(new_n694), .A3(new_n588), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n691), .A2(new_n306), .A3(new_n368), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(KEYINPUT41), .B(G113), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G15));
  NAND4_X1  g513(.A1(new_n635), .A2(new_n306), .A3(new_n368), .A4(new_n696), .ZN(new_n700));
  XOR2_X1   g514(.A(KEYINPUT104), .B(G116), .Z(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G18));
  OAI21_X1  g516(.A(new_n541), .B1(new_n621), .B2(new_n437), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n703), .A2(new_n695), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n306), .A2(new_n704), .A3(new_n537), .A4(new_n643), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G119), .ZN(G21));
  INV_X1    g520(.A(new_n368), .ZN(new_n707));
  AOI21_X1  g521(.A(G902), .B1(new_n274), .B2(new_n279), .ZN(new_n708));
  INV_X1    g522(.A(G472), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n303), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  OAI211_X1 g525(.A(new_n678), .B(new_n541), .C1(new_n621), .C2(new_n437), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n712), .A2(new_n695), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n711), .A2(new_n713), .A3(new_n535), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G122), .ZN(G24));
  NOR3_X1   g529(.A1(new_n684), .A2(new_n710), .A3(KEYINPUT105), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT105), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n602), .B1(new_n606), .B2(G472), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n717), .B1(new_n718), .B2(new_n643), .ZN(new_n719));
  OAI211_X1 g533(.A(new_n704), .B(new_n688), .C1(new_n716), .C2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G125), .ZN(G27));
  INV_X1    g535(.A(KEYINPUT106), .ZN(new_n722));
  AND3_X1   g536(.A1(new_n588), .A2(new_n595), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n722), .B1(new_n588), .B2(new_n595), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n694), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT107), .ZN(new_n726));
  OR2_X1    g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n542), .B1(new_n440), .B2(new_n538), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n725), .A2(new_n726), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n727), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT108), .ZN(new_n731));
  INV_X1    g545(.A(new_n369), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n730), .A2(new_n731), .A3(new_n732), .A4(new_n688), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT42), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n727), .A2(new_n728), .A3(new_n688), .A4(new_n729), .ZN(new_n735));
  OAI21_X1  g549(.A(KEYINPUT108), .B1(new_n735), .B2(new_n369), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n733), .A2(new_n734), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n303), .A2(new_n187), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n295), .A2(new_n305), .A3(new_n738), .ZN(new_n739));
  AND2_X1   g553(.A1(new_n739), .A2(new_n368), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n730), .A2(KEYINPUT42), .A3(new_n688), .A4(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n737), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G131), .ZN(G33));
  NAND2_X1  g557(.A1(new_n664), .A2(KEYINPUT109), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n730), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n732), .B1(new_n664), .B2(KEYINPUT109), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(new_n197), .ZN(G36));
  XOR2_X1   g562(.A(new_n594), .B(KEYINPUT45), .Z(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(G469), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT110), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(G469), .A2(G902), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT46), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n752), .A2(KEYINPUT46), .A3(new_n753), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(new_n588), .A3(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n758), .A2(new_n694), .A3(new_n670), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n617), .A2(new_n488), .A3(new_n494), .ZN(new_n761));
  XOR2_X1   g575(.A(new_n761), .B(KEYINPUT43), .Z(new_n762));
  NAND2_X1  g576(.A1(new_n604), .A2(new_n607), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(new_n763), .A3(new_n643), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT44), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OR2_X1    g580(.A1(new_n764), .A2(new_n765), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT111), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n767), .A2(new_n768), .A3(new_n728), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n768), .B1(new_n767), .B2(new_n728), .ZN(new_n770));
  OAI211_X1 g584(.A(new_n760), .B(new_n766), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G137), .ZN(G39));
  NAND2_X1  g586(.A1(new_n758), .A2(new_n694), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(KEYINPUT47), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n304), .B1(new_n604), .B2(new_n187), .ZN(new_n775));
  AND4_X1   g589(.A1(new_n775), .A2(new_n295), .A3(new_n688), .A4(new_n707), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT47), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n758), .A2(new_n777), .A3(new_n694), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n774), .A2(new_n728), .A3(new_n776), .A4(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G140), .ZN(G42));
  NAND2_X1  g594(.A1(new_n774), .A2(new_n778), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n693), .A2(new_n588), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n781), .B1(new_n694), .B2(new_n782), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n762), .A2(new_n529), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n784), .A2(new_n711), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n783), .A2(new_n728), .A3(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n785), .A2(new_n542), .A3(new_n668), .A4(new_n696), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n787), .A2(KEYINPUT50), .ZN(new_n788));
  OR2_X1    g602(.A1(new_n716), .A2(new_n719), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n728), .A2(new_n696), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n784), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n677), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n790), .A2(new_n792), .A3(new_n368), .A4(new_n529), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n793), .A2(new_n495), .A3(new_n617), .ZN(new_n794));
  AOI211_X1 g608(.A(new_n791), .B(new_n794), .C1(new_n787), .C2(KEYINPUT50), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n786), .A2(new_n788), .A3(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT51), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n786), .A2(KEYINPUT51), .A3(new_n788), .A4(new_n795), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n785), .A2(new_n704), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n784), .A2(new_n740), .A3(new_n790), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT48), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n793), .A2(new_n618), .A3(new_n619), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n801), .A2(new_n802), .ZN(new_n805));
  NOR4_X1   g619(.A1(new_n800), .A2(new_n803), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n798), .A2(new_n799), .A3(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT115), .ZN(new_n808));
  XOR2_X1   g622(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n643), .B1(new_n775), .B2(new_n676), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT113), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n712), .A2(new_n725), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n811), .A2(new_n812), .A3(new_n659), .A4(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n813), .A2(new_n677), .A3(new_n684), .A4(new_n659), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(KEYINPUT113), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n720), .B(new_n689), .C1(new_n652), .C2(new_n664), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n808), .B(new_n810), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n818), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n820), .A2(KEYINPUT52), .A3(new_n816), .A4(new_n814), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n684), .B1(new_n775), .B2(new_n295), .ZN(new_n823));
  AOI21_X1  g637(.A(KEYINPUT102), .B1(new_n633), .B2(new_n659), .ZN(new_n824));
  AND4_X1   g638(.A1(KEYINPUT102), .A2(new_n655), .A3(new_n656), .A4(new_n659), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n823), .B(new_n651), .C1(new_n826), .C2(new_n688), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n827), .A2(new_n720), .A3(new_n816), .A4(new_n814), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n808), .B1(new_n828), .B2(new_n810), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n822), .A2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n747), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n597), .B1(new_n646), .B2(new_n369), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n697), .A2(new_n700), .A3(new_n705), .A4(new_n714), .ZN(new_n833));
  INV_X1    g647(.A(new_n620), .ZN(new_n834));
  AOI22_X1  g648(.A1(new_n656), .A2(new_n488), .B1(new_n495), .B2(new_n617), .ZN(new_n835));
  NOR4_X1   g649(.A1(new_n608), .A2(new_n667), .A3(new_n834), .A4(new_n835), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n832), .A2(new_n833), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n789), .A2(new_n688), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n727), .A2(new_n728), .A3(new_n729), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n605), .A2(new_n494), .A3(new_n659), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n823), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n728), .A2(new_n522), .A3(new_n655), .ZN(new_n842));
  OAI22_X1  g656(.A1(new_n838), .A2(new_n839), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n742), .A2(new_n831), .A3(new_n837), .A4(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(KEYINPUT53), .B1(new_n830), .B2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT52), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n828), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(new_n821), .ZN(new_n849));
  NOR4_X1   g663(.A1(new_n843), .A2(new_n832), .A3(new_n833), .A4(new_n836), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n747), .B1(new_n737), .B2(new_n741), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n849), .A2(new_n850), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT54), .B1(new_n846), .B2(new_n853), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n850), .A2(new_n851), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n855), .A2(KEYINPUT53), .A3(new_n849), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(KEYINPUT116), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n852), .B1(new_n830), .B2(new_n845), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT116), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n855), .A2(new_n859), .A3(KEYINPUT53), .A4(new_n849), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n857), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n854), .B1(new_n861), .B2(KEYINPUT54), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n527), .B(KEYINPUT117), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n807), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n864), .B1(G952), .B2(G953), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n368), .A2(new_n694), .A3(new_n541), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(KEYINPUT112), .ZN(new_n867));
  AOI211_X1 g681(.A(new_n761), .B(new_n867), .C1(KEYINPUT49), .C2(new_n782), .ZN(new_n868));
  OR2_X1    g682(.A1(new_n782), .A2(KEYINPUT49), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n868), .A2(new_n668), .A3(new_n792), .A4(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n865), .A2(new_n870), .ZN(G75));
  XNOR2_X1  g685(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n846), .A2(G210), .A3(G902), .A4(new_n853), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT56), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n419), .A2(new_n425), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(new_n424), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n874), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n877), .B1(new_n874), .B2(new_n875), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n873), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n874), .A2(new_n875), .ZN(new_n881));
  INV_X1    g695(.A(new_n877), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n874), .A2(new_n875), .A3(new_n877), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n883), .A2(new_n872), .A3(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n350), .A2(G952), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n880), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(KEYINPUT119), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT119), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n880), .A2(new_n885), .A3(new_n890), .A4(new_n887), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n889), .A2(new_n891), .ZN(G51));
  AND2_X1   g706(.A1(new_n846), .A2(new_n853), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n893), .A2(KEYINPUT120), .A3(KEYINPUT54), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT120), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n846), .A2(new_n853), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT54), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n894), .B(new_n898), .C1(KEYINPUT54), .C2(new_n893), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n753), .B(KEYINPUT57), .Z(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n586), .ZN(new_n902));
  OR3_X1    g716(.A1(new_n896), .A2(new_n292), .A3(new_n752), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n886), .B1(new_n902), .B2(new_n903), .ZN(G54));
  NAND4_X1  g718(.A1(new_n893), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n905));
  INV_X1    g719(.A(new_n482), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n905), .A2(new_n906), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n907), .A2(new_n908), .A3(new_n886), .ZN(G60));
  NAND2_X1  g723(.A1(G478), .A2(G902), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n910), .B(KEYINPUT59), .Z(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n899), .A2(new_n614), .A3(new_n613), .A4(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n613), .A2(new_n614), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n914), .B1(new_n862), .B2(new_n911), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n913), .A2(new_n887), .A3(new_n915), .ZN(G63));
  NAND2_X1  g730(.A1(G217), .A2(G902), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT60), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n896), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n641), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n920), .B(new_n887), .C1(new_n357), .C2(new_n919), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n921), .B(KEYINPUT61), .Z(G66));
  INV_X1    g736(.A(new_n350), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n837), .A2(new_n923), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT121), .Z(new_n925));
  AOI21_X1  g739(.A(new_n249), .B1(new_n533), .B2(G224), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT122), .Z(new_n928));
  OAI21_X1  g742(.A(new_n876), .B1(G898), .B2(new_n350), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n928), .B(new_n929), .ZN(G69));
  NAND2_X1  g744(.A1(new_n771), .A2(new_n820), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT125), .ZN(new_n932));
  INV_X1    g746(.A(new_n712), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n760), .A2(new_n933), .A3(new_n740), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n934), .A2(new_n851), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n932), .A2(new_n350), .A3(new_n779), .A4(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n221), .A2(new_n239), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(new_n469), .Z(new_n938));
  OAI211_X1 g752(.A(new_n936), .B(new_n938), .C1(new_n657), .C2(new_n350), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n938), .B(KEYINPUT123), .Z(new_n940));
  NOR3_X1   g754(.A1(new_n369), .A2(new_n671), .A3(new_n835), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n728), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n771), .A2(new_n779), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n818), .B1(KEYINPUT124), .B2(KEYINPUT62), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n685), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g759(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  OR2_X1    g761(.A1(new_n945), .A2(new_n946), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n943), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n940), .B1(new_n949), .B2(new_n923), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n939), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n350), .B1(G227), .B2(G900), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n952), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n939), .A2(new_n954), .A3(new_n950), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n953), .A2(new_n955), .ZN(G72));
  XNOR2_X1  g770(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n709), .A2(new_n292), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n957), .B(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n959), .B1(new_n949), .B2(new_n837), .ZN(new_n960));
  INV_X1    g774(.A(new_n673), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n887), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n290), .B(KEYINPUT127), .Z(new_n963));
  OAI21_X1  g777(.A(new_n861), .B1(new_n277), .B2(new_n963), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n964), .A2(new_n959), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n932), .A2(new_n779), .A3(new_n837), .A4(new_n935), .ZN(new_n966));
  INV_X1    g780(.A(new_n959), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n262), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  AOI211_X1 g782(.A(new_n962), .B(new_n965), .C1(new_n248), .C2(new_n968), .ZN(G57));
endmodule


