

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U552 ( .A1(n632), .A2(n775), .ZN(n633) );
  NOR2_X1 U553 ( .A1(n615), .A2(n889), .ZN(n617) );
  NOR2_X2 U554 ( .A1(n581), .A2(n548), .ZN(n802) );
  NOR2_X2 U555 ( .A1(n662), .A2(n661), .ZN(n663) );
  INV_X1 U556 ( .A(n912), .ZN(n711) );
  BUF_X2 U557 ( .A(n615), .Z(n683) );
  NAND2_X1 U558 ( .A1(n724), .A2(G138), .ZN(n604) );
  XNOR2_X1 U559 ( .A(n631), .B(KEYINPUT76), .ZN(n775) );
  BUF_X1 U560 ( .A(n609), .Z(n990) );
  BUF_X2 U561 ( .A(n603), .Z(n994) );
  BUF_X1 U562 ( .A(n775), .Z(n1020) );
  XNOR2_X1 U563 ( .A(KEYINPUT108), .B(n769), .ZN(n520) );
  OR2_X1 U564 ( .A1(n722), .A2(n721), .ZN(n521) );
  AND2_X1 U565 ( .A1(n763), .A2(n756), .ZN(n522) );
  NOR2_X1 U566 ( .A1(n711), .A2(n710), .ZN(n523) );
  AND2_X1 U567 ( .A1(n917), .A2(n705), .ZN(n524) );
  XNOR2_X1 U568 ( .A(KEYINPUT32), .B(KEYINPUT105), .ZN(n525) );
  AND2_X1 U569 ( .A1(n704), .A2(n703), .ZN(n526) );
  INV_X1 U570 ( .A(KEYINPUT26), .ZN(n616) );
  NOR2_X1 U571 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U572 ( .A(n663), .B(KEYINPUT29), .ZN(n691) );
  INV_X1 U573 ( .A(n920), .ZN(n703) );
  NAND2_X1 U574 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U575 ( .A(n699), .B(n525), .ZN(n700) );
  NAND2_X1 U576 ( .A1(n714), .A2(n526), .ZN(n706) );
  XNOR2_X1 U577 ( .A(KEYINPUT74), .B(KEYINPUT14), .ZN(n624) );
  INV_X1 U578 ( .A(KEYINPUT17), .ZN(n535) );
  AND2_X1 U579 ( .A1(n528), .A2(G2105), .ZN(n609) );
  INV_X1 U580 ( .A(G2104), .ZN(n528) );
  NOR2_X1 U581 ( .A1(G2105), .A2(n528), .ZN(n603) );
  NOR2_X1 U582 ( .A1(n548), .A2(G543), .ZN(n549) );
  NOR2_X2 U583 ( .A1(G651), .A2(G543), .ZN(n805) );
  NOR2_X1 U584 ( .A1(G651), .A2(n581), .ZN(n809) );
  NOR2_X1 U585 ( .A1(n541), .A2(n540), .ZN(n602) );
  BUF_X1 U586 ( .A(n602), .Z(G160) );
  NAND2_X1 U587 ( .A1(n603), .A2(G101), .ZN(n527) );
  XNOR2_X1 U588 ( .A(KEYINPUT23), .B(n527), .ZN(n531) );
  NAND2_X1 U589 ( .A1(n609), .A2(G125), .ZN(n529) );
  XNOR2_X1 U590 ( .A(KEYINPUT65), .B(n529), .ZN(n530) );
  NOR2_X1 U591 ( .A1(n531), .A2(n530), .ZN(n533) );
  INV_X1 U592 ( .A(KEYINPUT66), .ZN(n532) );
  XNOR2_X1 U593 ( .A(n533), .B(n532), .ZN(n541) );
  NAND2_X1 U594 ( .A1(G2105), .A2(G2104), .ZN(n534) );
  XNOR2_X2 U595 ( .A(n534), .B(KEYINPUT67), .ZN(n991) );
  NAND2_X1 U596 ( .A1(G113), .A2(n991), .ZN(n538) );
  NOR2_X2 U597 ( .A1(G2105), .A2(G2104), .ZN(n536) );
  XNOR2_X2 U598 ( .A(n536), .B(n535), .ZN(n724) );
  NAND2_X1 U599 ( .A1(G137), .A2(n724), .ZN(n537) );
  NAND2_X1 U600 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U601 ( .A(n539), .B(KEYINPUT68), .ZN(n540) );
  XOR2_X1 U602 ( .A(KEYINPUT0), .B(G543), .Z(n581) );
  NAND2_X1 U603 ( .A1(G53), .A2(n809), .ZN(n542) );
  XOR2_X1 U604 ( .A(KEYINPUT72), .B(n542), .Z(n547) );
  INV_X1 U605 ( .A(G651), .ZN(n548) );
  NAND2_X1 U606 ( .A1(G78), .A2(n802), .ZN(n544) );
  NAND2_X1 U607 ( .A1(G91), .A2(n805), .ZN(n543) );
  NAND2_X1 U608 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U609 ( .A(KEYINPUT71), .B(n545), .Z(n546) );
  NOR2_X1 U610 ( .A1(n547), .A2(n546), .ZN(n551) );
  XOR2_X2 U611 ( .A(KEYINPUT1), .B(n549), .Z(n801) );
  NAND2_X1 U612 ( .A1(n801), .A2(G65), .ZN(n550) );
  NAND2_X1 U613 ( .A1(n551), .A2(n550), .ZN(G299) );
  NAND2_X1 U614 ( .A1(G64), .A2(n801), .ZN(n553) );
  NAND2_X1 U615 ( .A1(G52), .A2(n809), .ZN(n552) );
  NAND2_X1 U616 ( .A1(n553), .A2(n552), .ZN(n558) );
  NAND2_X1 U617 ( .A1(G77), .A2(n802), .ZN(n555) );
  NAND2_X1 U618 ( .A1(G90), .A2(n805), .ZN(n554) );
  NAND2_X1 U619 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U620 ( .A(KEYINPUT9), .B(n556), .Z(n557) );
  NOR2_X1 U621 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U622 ( .A(KEYINPUT70), .B(n559), .ZN(G171) );
  NAND2_X1 U623 ( .A1(n805), .A2(G89), .ZN(n560) );
  XNOR2_X1 U624 ( .A(n560), .B(KEYINPUT4), .ZN(n562) );
  NAND2_X1 U625 ( .A1(G76), .A2(n802), .ZN(n561) );
  NAND2_X1 U626 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U627 ( .A(KEYINPUT5), .B(n563), .ZN(n569) );
  NAND2_X1 U628 ( .A1(n809), .A2(G51), .ZN(n564) );
  XOR2_X1 U629 ( .A(KEYINPUT79), .B(n564), .Z(n566) );
  NAND2_X1 U630 ( .A1(n801), .A2(G63), .ZN(n565) );
  NAND2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U632 ( .A(KEYINPUT6), .B(n567), .Z(n568) );
  NAND2_X1 U633 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U634 ( .A(KEYINPUT7), .B(n570), .ZN(G168) );
  NAND2_X1 U635 ( .A1(G75), .A2(n802), .ZN(n572) );
  NAND2_X1 U636 ( .A1(G88), .A2(n805), .ZN(n571) );
  NAND2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n576) );
  NAND2_X1 U638 ( .A1(G62), .A2(n801), .ZN(n574) );
  NAND2_X1 U639 ( .A1(G50), .A2(n809), .ZN(n573) );
  NAND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U641 ( .A1(n576), .A2(n575), .ZN(G166) );
  INV_X1 U642 ( .A(G166), .ZN(G303) );
  XOR2_X1 U643 ( .A(G168), .B(KEYINPUT8), .Z(n577) );
  XNOR2_X1 U644 ( .A(KEYINPUT80), .B(n577), .ZN(G286) );
  NAND2_X1 U645 ( .A1(G49), .A2(n809), .ZN(n579) );
  NAND2_X1 U646 ( .A1(G74), .A2(G651), .ZN(n578) );
  NAND2_X1 U647 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X1 U648 ( .A1(n801), .A2(n580), .ZN(n583) );
  NAND2_X1 U649 ( .A1(n581), .A2(G87), .ZN(n582) );
  NAND2_X1 U650 ( .A1(n583), .A2(n582), .ZN(G288) );
  NAND2_X1 U651 ( .A1(n801), .A2(G61), .ZN(n584) );
  XNOR2_X1 U652 ( .A(n584), .B(KEYINPUT84), .ZN(n586) );
  NAND2_X1 U653 ( .A1(G86), .A2(n805), .ZN(n585) );
  NAND2_X1 U654 ( .A1(n586), .A2(n585), .ZN(n590) );
  XOR2_X1 U655 ( .A(KEYINPUT85), .B(KEYINPUT2), .Z(n588) );
  NAND2_X1 U656 ( .A1(n802), .A2(G73), .ZN(n587) );
  XOR2_X1 U657 ( .A(n588), .B(n587), .Z(n589) );
  NOR2_X1 U658 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U659 ( .A(KEYINPUT86), .B(n591), .ZN(n594) );
  NAND2_X1 U660 ( .A1(n809), .A2(G48), .ZN(n592) );
  XOR2_X1 U661 ( .A(KEYINPUT87), .B(n592), .Z(n593) );
  NAND2_X1 U662 ( .A1(n594), .A2(n593), .ZN(G305) );
  NAND2_X1 U663 ( .A1(G72), .A2(n802), .ZN(n596) );
  NAND2_X1 U664 ( .A1(G85), .A2(n805), .ZN(n595) );
  NAND2_X1 U665 ( .A1(n596), .A2(n595), .ZN(n599) );
  NAND2_X1 U666 ( .A1(G60), .A2(n801), .ZN(n597) );
  XNOR2_X1 U667 ( .A(KEYINPUT69), .B(n597), .ZN(n598) );
  NOR2_X1 U668 ( .A1(n599), .A2(n598), .ZN(n601) );
  NAND2_X1 U669 ( .A1(n809), .A2(G47), .ZN(n600) );
  NAND2_X1 U670 ( .A1(n601), .A2(n600), .ZN(G290) );
  NAND2_X1 U671 ( .A1(n602), .A2(G40), .ZN(n735) );
  INV_X1 U672 ( .A(n735), .ZN(n614) );
  NAND2_X1 U673 ( .A1(G102), .A2(n994), .ZN(n605) );
  NAND2_X1 U674 ( .A1(n605), .A2(n604), .ZN(n606) );
  NAND2_X1 U675 ( .A1(KEYINPUT92), .A2(n606), .ZN(n608) );
  OR2_X1 U676 ( .A1(KEYINPUT92), .A2(n606), .ZN(n607) );
  NAND2_X1 U677 ( .A1(n608), .A2(n607), .ZN(n613) );
  NAND2_X1 U678 ( .A1(G126), .A2(n990), .ZN(n611) );
  NAND2_X1 U679 ( .A1(G114), .A2(n991), .ZN(n610) );
  NAND2_X1 U680 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U681 ( .A1(n613), .A2(n612), .ZN(n772) );
  NOR2_X1 U682 ( .A1(n772), .A2(G1384), .ZN(n734) );
  NAND2_X1 U683 ( .A1(n614), .A2(n734), .ZN(n615) );
  NOR2_X1 U684 ( .A1(G2084), .A2(n683), .ZN(n671) );
  NAND2_X1 U685 ( .A1(G8), .A2(n671), .ZN(n682) );
  INV_X1 U686 ( .A(G1996), .ZN(n889) );
  XNOR2_X1 U687 ( .A(n617), .B(n616), .ZN(n619) );
  NAND2_X1 U688 ( .A1(n683), .A2(G1341), .ZN(n618) );
  NAND2_X1 U689 ( .A1(n619), .A2(n618), .ZN(n632) );
  NAND2_X1 U690 ( .A1(n805), .A2(G81), .ZN(n620) );
  XNOR2_X1 U691 ( .A(n620), .B(KEYINPUT12), .ZN(n622) );
  NAND2_X1 U692 ( .A1(G68), .A2(n802), .ZN(n621) );
  NAND2_X1 U693 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U694 ( .A(n623), .B(KEYINPUT13), .ZN(n627) );
  NAND2_X1 U695 ( .A1(G56), .A2(n801), .ZN(n625) );
  XNOR2_X1 U696 ( .A(n625), .B(n624), .ZN(n626) );
  NAND2_X1 U697 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U698 ( .A(n628), .B(KEYINPUT75), .ZN(n630) );
  NAND2_X1 U699 ( .A1(G43), .A2(n809), .ZN(n629) );
  NAND2_X1 U700 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U701 ( .A(n633), .B(KEYINPUT64), .ZN(n647) );
  NAND2_X1 U702 ( .A1(G79), .A2(n802), .ZN(n635) );
  NAND2_X1 U703 ( .A1(G92), .A2(n805), .ZN(n634) );
  NAND2_X1 U704 ( .A1(n635), .A2(n634), .ZN(n639) );
  NAND2_X1 U705 ( .A1(G66), .A2(n801), .ZN(n637) );
  NAND2_X1 U706 ( .A1(G54), .A2(n809), .ZN(n636) );
  NAND2_X1 U707 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U708 ( .A1(n639), .A2(n638), .ZN(n640) );
  XOR2_X1 U709 ( .A(KEYINPUT15), .B(n640), .Z(n1017) );
  NAND2_X1 U710 ( .A1(n647), .A2(n1017), .ZN(n641) );
  XNOR2_X1 U711 ( .A(n641), .B(KEYINPUT100), .ZN(n645) );
  NOR2_X1 U712 ( .A1(G2067), .A2(n683), .ZN(n643) );
  INV_X1 U713 ( .A(n683), .ZN(n664) );
  NOR2_X1 U714 ( .A1(n664), .A2(G1348), .ZN(n642) );
  NOR2_X1 U715 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U716 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U717 ( .A(n646), .B(KEYINPUT101), .ZN(n649) );
  NOR2_X1 U718 ( .A1(n647), .A2(n1017), .ZN(n648) );
  XNOR2_X1 U719 ( .A(n650), .B(KEYINPUT102), .ZN(n656) );
  NAND2_X1 U720 ( .A1(n664), .A2(G2072), .ZN(n651) );
  XOR2_X1 U721 ( .A(KEYINPUT27), .B(n651), .Z(n653) );
  NAND2_X1 U722 ( .A1(G1956), .A2(n683), .ZN(n652) );
  NAND2_X1 U723 ( .A1(n653), .A2(n652), .ZN(n658) );
  NOR2_X1 U724 ( .A1(G299), .A2(n658), .ZN(n654) );
  XOR2_X1 U725 ( .A(KEYINPUT103), .B(n654), .Z(n655) );
  NOR2_X1 U726 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U727 ( .A(KEYINPUT104), .B(n657), .ZN(n662) );
  NAND2_X1 U728 ( .A1(n658), .A2(G299), .ZN(n659) );
  XNOR2_X1 U729 ( .A(n659), .B(KEYINPUT28), .ZN(n660) );
  XNOR2_X1 U730 ( .A(KEYINPUT99), .B(n660), .ZN(n661) );
  XOR2_X1 U731 ( .A(G1961), .B(KEYINPUT98), .Z(n946) );
  NAND2_X1 U732 ( .A1(n946), .A2(n683), .ZN(n666) );
  XNOR2_X1 U733 ( .A(G2078), .B(KEYINPUT25), .ZN(n892) );
  NAND2_X1 U734 ( .A1(n664), .A2(n892), .ZN(n665) );
  NAND2_X1 U735 ( .A1(n666), .A2(n665), .ZN(n674) );
  NAND2_X1 U736 ( .A1(n674), .A2(G171), .ZN(n689) );
  NAND2_X1 U737 ( .A1(G8), .A2(n683), .ZN(n722) );
  NOR2_X1 U738 ( .A1(n722), .A2(G1966), .ZN(n667) );
  XNOR2_X1 U739 ( .A(n667), .B(KEYINPUT97), .ZN(n669) );
  AND2_X1 U740 ( .A1(n689), .A2(n669), .ZN(n668) );
  NAND2_X1 U741 ( .A1(n691), .A2(n668), .ZN(n680) );
  INV_X1 U742 ( .A(n669), .ZN(n678) );
  NAND2_X1 U743 ( .A1(G8), .A2(n669), .ZN(n670) );
  NOR2_X1 U744 ( .A1(n671), .A2(n670), .ZN(n672) );
  XOR2_X1 U745 ( .A(KEYINPUT30), .B(n672), .Z(n673) );
  NOR2_X1 U746 ( .A1(G168), .A2(n673), .ZN(n676) );
  NOR2_X1 U747 ( .A1(n674), .A2(G171), .ZN(n675) );
  NOR2_X1 U748 ( .A1(n676), .A2(n675), .ZN(n677) );
  XOR2_X1 U749 ( .A(KEYINPUT31), .B(n677), .Z(n694) );
  OR2_X1 U750 ( .A1(n678), .A2(n694), .ZN(n679) );
  NAND2_X1 U751 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U752 ( .A1(n682), .A2(n681), .ZN(n701) );
  NOR2_X1 U753 ( .A1(G1971), .A2(n722), .ZN(n685) );
  NOR2_X1 U754 ( .A1(G2090), .A2(n683), .ZN(n684) );
  NOR2_X1 U755 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U756 ( .A1(n686), .A2(G303), .ZN(n693) );
  INV_X1 U757 ( .A(n693), .ZN(n687) );
  OR2_X1 U758 ( .A1(n687), .A2(G286), .ZN(n688) );
  AND2_X1 U759 ( .A1(G8), .A2(n688), .ZN(n692) );
  AND2_X1 U760 ( .A1(n689), .A2(n692), .ZN(n690) );
  NAND2_X1 U761 ( .A1(n691), .A2(n690), .ZN(n698) );
  INV_X1 U762 ( .A(n692), .ZN(n696) );
  AND2_X1 U763 ( .A1(n694), .A2(n693), .ZN(n695) );
  OR2_X1 U764 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U765 ( .A1(n701), .A2(n700), .ZN(n714) );
  NOR2_X1 U766 ( .A1(G1971), .A2(G303), .ZN(n702) );
  XOR2_X1 U767 ( .A(n702), .B(KEYINPUT106), .Z(n704) );
  NOR2_X1 U768 ( .A1(G1976), .A2(G288), .ZN(n920) );
  NAND2_X1 U769 ( .A1(G1976), .A2(G288), .ZN(n917) );
  INV_X1 U770 ( .A(n722), .ZN(n705) );
  NAND2_X1 U771 ( .A1(n706), .A2(n524), .ZN(n708) );
  INV_X1 U772 ( .A(KEYINPUT33), .ZN(n707) );
  NAND2_X1 U773 ( .A1(n708), .A2(n707), .ZN(n712) );
  XOR2_X1 U774 ( .A(G1981), .B(G305), .Z(n912) );
  NAND2_X1 U775 ( .A1(n920), .A2(KEYINPUT33), .ZN(n709) );
  NOR2_X1 U776 ( .A1(n709), .A2(n722), .ZN(n710) );
  NAND2_X1 U777 ( .A1(n712), .A2(n523), .ZN(n718) );
  NOR2_X1 U778 ( .A1(G2090), .A2(G303), .ZN(n713) );
  NAND2_X1 U779 ( .A1(G8), .A2(n713), .ZN(n715) );
  NAND2_X1 U780 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U781 ( .A1(n716), .A2(n722), .ZN(n717) );
  NAND2_X1 U782 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U783 ( .A(n719), .B(KEYINPUT107), .ZN(n723) );
  NOR2_X1 U784 ( .A1(G1981), .A2(G305), .ZN(n720) );
  XOR2_X1 U785 ( .A(n720), .B(KEYINPUT24), .Z(n721) );
  NAND2_X1 U786 ( .A1(n723), .A2(n521), .ZN(n757) );
  NAND2_X1 U787 ( .A1(G104), .A2(n994), .ZN(n726) );
  NAND2_X1 U788 ( .A1(G140), .A2(n724), .ZN(n725) );
  NAND2_X1 U789 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U790 ( .A(KEYINPUT34), .B(n727), .ZN(n732) );
  NAND2_X1 U791 ( .A1(G128), .A2(n990), .ZN(n729) );
  NAND2_X1 U792 ( .A1(G116), .A2(n991), .ZN(n728) );
  NAND2_X1 U793 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U794 ( .A(KEYINPUT35), .B(n730), .Z(n731) );
  NOR2_X1 U795 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U796 ( .A(KEYINPUT36), .B(n733), .ZN(n1001) );
  XNOR2_X1 U797 ( .A(G2067), .B(KEYINPUT37), .ZN(n765) );
  NOR2_X1 U798 ( .A1(n1001), .A2(n765), .ZN(n882) );
  NOR2_X1 U799 ( .A1(n734), .A2(n735), .ZN(n768) );
  NAND2_X1 U800 ( .A1(n882), .A2(n768), .ZN(n763) );
  NAND2_X1 U801 ( .A1(G105), .A2(n994), .ZN(n736) );
  XOR2_X1 U802 ( .A(KEYINPUT38), .B(n736), .Z(n739) );
  NAND2_X1 U803 ( .A1(n991), .A2(G117), .ZN(n737) );
  XOR2_X1 U804 ( .A(KEYINPUT94), .B(n737), .Z(n738) );
  NOR2_X1 U805 ( .A1(n739), .A2(n738), .ZN(n741) );
  NAND2_X1 U806 ( .A1(n990), .A2(G129), .ZN(n740) );
  NAND2_X1 U807 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U808 ( .A(n742), .B(KEYINPUT95), .ZN(n744) );
  NAND2_X1 U809 ( .A1(G141), .A2(n724), .ZN(n743) );
  NAND2_X1 U810 ( .A1(n744), .A2(n743), .ZN(n1013) );
  NAND2_X1 U811 ( .A1(G1996), .A2(n1013), .ZN(n745) );
  XNOR2_X1 U812 ( .A(n745), .B(KEYINPUT96), .ZN(n754) );
  NAND2_X1 U813 ( .A1(G119), .A2(n990), .ZN(n747) );
  NAND2_X1 U814 ( .A1(G131), .A2(n724), .ZN(n746) );
  NAND2_X1 U815 ( .A1(n747), .A2(n746), .ZN(n750) );
  NAND2_X1 U816 ( .A1(G95), .A2(n994), .ZN(n748) );
  XNOR2_X1 U817 ( .A(KEYINPUT93), .B(n748), .ZN(n749) );
  NOR2_X1 U818 ( .A1(n750), .A2(n749), .ZN(n752) );
  NAND2_X1 U819 ( .A1(n991), .A2(G107), .ZN(n751) );
  NAND2_X1 U820 ( .A1(n752), .A2(n751), .ZN(n1002) );
  NAND2_X1 U821 ( .A1(G1991), .A2(n1002), .ZN(n753) );
  NAND2_X1 U822 ( .A1(n754), .A2(n753), .ZN(n760) );
  INV_X1 U823 ( .A(n760), .ZN(n866) );
  XOR2_X1 U824 ( .A(G1986), .B(G290), .Z(n922) );
  NAND2_X1 U825 ( .A1(n866), .A2(n922), .ZN(n755) );
  NAND2_X1 U826 ( .A1(n768), .A2(n755), .ZN(n756) );
  NAND2_X1 U827 ( .A1(n757), .A2(n522), .ZN(n770) );
  NOR2_X1 U828 ( .A1(G1996), .A2(n1013), .ZN(n869) );
  NOR2_X1 U829 ( .A1(G1986), .A2(G290), .ZN(n758) );
  NOR2_X1 U830 ( .A1(G1991), .A2(n1002), .ZN(n874) );
  NOR2_X1 U831 ( .A1(n758), .A2(n874), .ZN(n759) );
  NOR2_X1 U832 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X1 U833 ( .A1(n869), .A2(n761), .ZN(n762) );
  XNOR2_X1 U834 ( .A(n762), .B(KEYINPUT39), .ZN(n764) );
  NAND2_X1 U835 ( .A1(n764), .A2(n763), .ZN(n766) );
  NAND2_X1 U836 ( .A1(n1001), .A2(n765), .ZN(n875) );
  NAND2_X1 U837 ( .A1(n766), .A2(n875), .ZN(n767) );
  NAND2_X1 U838 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U839 ( .A1(n770), .A2(n520), .ZN(n771) );
  XNOR2_X1 U840 ( .A(n771), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U841 ( .A1(G452), .A2(G94), .ZN(G173) );
  BUF_X1 U842 ( .A(n772), .Z(G164) );
  INV_X1 U843 ( .A(G132), .ZN(G219) );
  INV_X1 U844 ( .A(G82), .ZN(G220) );
  INV_X1 U845 ( .A(G120), .ZN(G236) );
  INV_X1 U846 ( .A(G69), .ZN(G235) );
  INV_X1 U847 ( .A(G108), .ZN(G238) );
  NAND2_X1 U848 ( .A1(G7), .A2(G661), .ZN(n773) );
  XNOR2_X1 U849 ( .A(n773), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U850 ( .A(G223), .B(KEYINPUT73), .ZN(n841) );
  NAND2_X1 U851 ( .A1(n841), .A2(G567), .ZN(n774) );
  XOR2_X1 U852 ( .A(KEYINPUT11), .B(n774), .Z(G234) );
  XOR2_X1 U853 ( .A(G860), .B(KEYINPUT77), .Z(n784) );
  INV_X1 U854 ( .A(n1020), .ZN(n776) );
  NAND2_X1 U855 ( .A1(n784), .A2(n776), .ZN(G153) );
  NAND2_X1 U856 ( .A1(G868), .A2(G171), .ZN(n778) );
  INV_X1 U857 ( .A(G868), .ZN(n822) );
  NAND2_X1 U858 ( .A1(n1017), .A2(n822), .ZN(n777) );
  NAND2_X1 U859 ( .A1(n778), .A2(n777), .ZN(n779) );
  XOR2_X1 U860 ( .A(KEYINPUT78), .B(n779), .Z(G284) );
  XNOR2_X1 U861 ( .A(KEYINPUT81), .B(G868), .ZN(n780) );
  NOR2_X1 U862 ( .A1(G286), .A2(n780), .ZN(n782) );
  NOR2_X1 U863 ( .A1(G868), .A2(G299), .ZN(n781) );
  NOR2_X1 U864 ( .A1(n782), .A2(n781), .ZN(G297) );
  INV_X1 U865 ( .A(n1017), .ZN(n786) );
  INV_X1 U866 ( .A(G559), .ZN(n783) );
  NOR2_X1 U867 ( .A1(n784), .A2(n783), .ZN(n785) );
  NOR2_X1 U868 ( .A1(n786), .A2(n785), .ZN(n787) );
  XOR2_X1 U869 ( .A(n787), .B(KEYINPUT16), .Z(n788) );
  XNOR2_X1 U870 ( .A(KEYINPUT82), .B(n788), .ZN(G148) );
  NOR2_X1 U871 ( .A1(n1020), .A2(G868), .ZN(n791) );
  NAND2_X1 U872 ( .A1(G868), .A2(n1017), .ZN(n789) );
  NOR2_X1 U873 ( .A1(G559), .A2(n789), .ZN(n790) );
  NOR2_X1 U874 ( .A1(n791), .A2(n790), .ZN(G282) );
  NAND2_X1 U875 ( .A1(n990), .A2(G123), .ZN(n792) );
  XNOR2_X1 U876 ( .A(n792), .B(KEYINPUT18), .ZN(n794) );
  NAND2_X1 U877 ( .A1(G99), .A2(n994), .ZN(n793) );
  NAND2_X1 U878 ( .A1(n794), .A2(n793), .ZN(n798) );
  NAND2_X1 U879 ( .A1(G135), .A2(n724), .ZN(n796) );
  NAND2_X1 U880 ( .A1(G111), .A2(n991), .ZN(n795) );
  NAND2_X1 U881 ( .A1(n796), .A2(n795), .ZN(n797) );
  NOR2_X1 U882 ( .A1(n798), .A2(n797), .ZN(n1006) );
  XNOR2_X1 U883 ( .A(n1006), .B(G2096), .ZN(n800) );
  INV_X1 U884 ( .A(G2100), .ZN(n799) );
  NAND2_X1 U885 ( .A1(n800), .A2(n799), .ZN(G156) );
  NAND2_X1 U886 ( .A1(G67), .A2(n801), .ZN(n804) );
  NAND2_X1 U887 ( .A1(G80), .A2(n802), .ZN(n803) );
  NAND2_X1 U888 ( .A1(n804), .A2(n803), .ZN(n808) );
  NAND2_X1 U889 ( .A1(G93), .A2(n805), .ZN(n806) );
  XNOR2_X1 U890 ( .A(KEYINPUT83), .B(n806), .ZN(n807) );
  NOR2_X1 U891 ( .A1(n808), .A2(n807), .ZN(n811) );
  NAND2_X1 U892 ( .A1(n809), .A2(G55), .ZN(n810) );
  NAND2_X1 U893 ( .A1(n811), .A2(n810), .ZN(n821) );
  NAND2_X1 U894 ( .A1(G559), .A2(n1017), .ZN(n812) );
  XNOR2_X1 U895 ( .A(n1020), .B(n812), .ZN(n819) );
  NOR2_X1 U896 ( .A1(n819), .A2(G860), .ZN(n813) );
  XOR2_X1 U897 ( .A(n821), .B(n813), .Z(G145) );
  XNOR2_X1 U898 ( .A(KEYINPUT19), .B(G303), .ZN(n814) );
  XNOR2_X1 U899 ( .A(n814), .B(G290), .ZN(n815) );
  XNOR2_X1 U900 ( .A(n815), .B(G288), .ZN(n816) );
  XNOR2_X1 U901 ( .A(n816), .B(n821), .ZN(n817) );
  XNOR2_X1 U902 ( .A(n817), .B(G305), .ZN(n818) );
  XNOR2_X1 U903 ( .A(n818), .B(G299), .ZN(n1016) );
  XOR2_X1 U904 ( .A(n819), .B(n1016), .Z(n820) );
  NAND2_X1 U905 ( .A1(n820), .A2(G868), .ZN(n824) );
  NAND2_X1 U906 ( .A1(n822), .A2(n821), .ZN(n823) );
  NAND2_X1 U907 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U908 ( .A(KEYINPUT88), .B(n825), .ZN(G295) );
  NAND2_X1 U909 ( .A1(G2078), .A2(G2084), .ZN(n826) );
  XNOR2_X1 U910 ( .A(n826), .B(KEYINPUT20), .ZN(n827) );
  XNOR2_X1 U911 ( .A(n827), .B(KEYINPUT89), .ZN(n828) );
  NAND2_X1 U912 ( .A1(n828), .A2(G2090), .ZN(n829) );
  XNOR2_X1 U913 ( .A(n829), .B(KEYINPUT90), .ZN(n830) );
  XNOR2_X1 U914 ( .A(n830), .B(KEYINPUT21), .ZN(n831) );
  NAND2_X1 U915 ( .A1(n831), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U916 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U917 ( .A1(G235), .A2(G236), .ZN(n832) );
  XNOR2_X1 U918 ( .A(n832), .B(KEYINPUT91), .ZN(n833) );
  NOR2_X1 U919 ( .A1(G238), .A2(n833), .ZN(n834) );
  NAND2_X1 U920 ( .A1(G57), .A2(n834), .ZN(n968) );
  NAND2_X1 U921 ( .A1(n968), .A2(G567), .ZN(n839) );
  NOR2_X1 U922 ( .A1(G220), .A2(G219), .ZN(n835) );
  XOR2_X1 U923 ( .A(KEYINPUT22), .B(n835), .Z(n836) );
  NOR2_X1 U924 ( .A1(G218), .A2(n836), .ZN(n837) );
  NAND2_X1 U925 ( .A1(G96), .A2(n837), .ZN(n969) );
  NAND2_X1 U926 ( .A1(n969), .A2(G2106), .ZN(n838) );
  NAND2_X1 U927 ( .A1(n839), .A2(n838), .ZN(n970) );
  NAND2_X1 U928 ( .A1(G483), .A2(G661), .ZN(n840) );
  NOR2_X1 U929 ( .A1(n970), .A2(n840), .ZN(n845) );
  NAND2_X1 U930 ( .A1(n845), .A2(G36), .ZN(G176) );
  NAND2_X1 U931 ( .A1(n841), .A2(G2106), .ZN(n842) );
  XNOR2_X1 U932 ( .A(n842), .B(KEYINPUT110), .ZN(G217) );
  AND2_X1 U933 ( .A1(G15), .A2(G2), .ZN(n843) );
  NAND2_X1 U934 ( .A1(G661), .A2(n843), .ZN(G259) );
  NAND2_X1 U935 ( .A1(G3), .A2(G1), .ZN(n844) );
  NAND2_X1 U936 ( .A1(n845), .A2(n844), .ZN(G188) );
  NAND2_X1 U938 ( .A1(n990), .A2(G124), .ZN(n846) );
  XNOR2_X1 U939 ( .A(n846), .B(KEYINPUT44), .ZN(n848) );
  NAND2_X1 U940 ( .A1(G136), .A2(n724), .ZN(n847) );
  NAND2_X1 U941 ( .A1(n848), .A2(n847), .ZN(n849) );
  XNOR2_X1 U942 ( .A(n849), .B(KEYINPUT113), .ZN(n851) );
  NAND2_X1 U943 ( .A1(G100), .A2(n994), .ZN(n850) );
  NAND2_X1 U944 ( .A1(n851), .A2(n850), .ZN(n854) );
  NAND2_X1 U945 ( .A1(n991), .A2(G112), .ZN(n852) );
  XOR2_X1 U946 ( .A(KEYINPUT114), .B(n852), .Z(n853) );
  NOR2_X1 U947 ( .A1(n854), .A2(n853), .ZN(G162) );
  INV_X1 U948 ( .A(KEYINPUT55), .ZN(n908) );
  XNOR2_X1 U949 ( .A(KEYINPUT52), .B(KEYINPUT118), .ZN(n884) );
  NAND2_X1 U950 ( .A1(G103), .A2(n994), .ZN(n856) );
  NAND2_X1 U951 ( .A1(G139), .A2(n724), .ZN(n855) );
  NAND2_X1 U952 ( .A1(n856), .A2(n855), .ZN(n862) );
  NAND2_X1 U953 ( .A1(G127), .A2(n990), .ZN(n858) );
  NAND2_X1 U954 ( .A1(G115), .A2(n991), .ZN(n857) );
  NAND2_X1 U955 ( .A1(n858), .A2(n857), .ZN(n859) );
  XNOR2_X1 U956 ( .A(KEYINPUT115), .B(n859), .ZN(n860) );
  XNOR2_X1 U957 ( .A(KEYINPUT47), .B(n860), .ZN(n861) );
  NOR2_X1 U958 ( .A1(n862), .A2(n861), .ZN(n1008) );
  XOR2_X1 U959 ( .A(G2072), .B(n1008), .Z(n864) );
  XOR2_X1 U960 ( .A(G164), .B(G2078), .Z(n863) );
  NOR2_X1 U961 ( .A1(n864), .A2(n863), .ZN(n865) );
  XNOR2_X1 U962 ( .A(KEYINPUT50), .B(n865), .ZN(n867) );
  NAND2_X1 U963 ( .A1(n867), .A2(n866), .ZN(n873) );
  XNOR2_X1 U964 ( .A(G2090), .B(G162), .ZN(n868) );
  XNOR2_X1 U965 ( .A(n868), .B(KEYINPUT117), .ZN(n870) );
  NOR2_X1 U966 ( .A1(n870), .A2(n869), .ZN(n871) );
  XNOR2_X1 U967 ( .A(KEYINPUT51), .B(n871), .ZN(n872) );
  NOR2_X1 U968 ( .A1(n873), .A2(n872), .ZN(n880) );
  NOR2_X1 U969 ( .A1(n874), .A2(n1006), .ZN(n876) );
  NAND2_X1 U970 ( .A1(n876), .A2(n875), .ZN(n878) );
  XOR2_X1 U971 ( .A(G160), .B(G2084), .Z(n877) );
  NOR2_X1 U972 ( .A1(n878), .A2(n877), .ZN(n879) );
  NAND2_X1 U973 ( .A1(n880), .A2(n879), .ZN(n881) );
  NOR2_X1 U974 ( .A1(n882), .A2(n881), .ZN(n883) );
  XNOR2_X1 U975 ( .A(n884), .B(n883), .ZN(n885) );
  NAND2_X1 U976 ( .A1(n908), .A2(n885), .ZN(n886) );
  NAND2_X1 U977 ( .A1(n886), .A2(G29), .ZN(n966) );
  XOR2_X1 U978 ( .A(G2090), .B(G35), .Z(n902) );
  XOR2_X1 U979 ( .A(G1991), .B(G25), .Z(n887) );
  NAND2_X1 U980 ( .A1(n887), .A2(G28), .ZN(n898) );
  XNOR2_X1 U981 ( .A(KEYINPUT119), .B(G2067), .ZN(n888) );
  XNOR2_X1 U982 ( .A(n888), .B(G26), .ZN(n896) );
  XOR2_X1 U983 ( .A(G2072), .B(G33), .Z(n891) );
  XNOR2_X1 U984 ( .A(n889), .B(G32), .ZN(n890) );
  NAND2_X1 U985 ( .A1(n891), .A2(n890), .ZN(n894) );
  XOR2_X1 U986 ( .A(G27), .B(n892), .Z(n893) );
  NOR2_X1 U987 ( .A1(n894), .A2(n893), .ZN(n895) );
  NAND2_X1 U988 ( .A1(n896), .A2(n895), .ZN(n897) );
  NOR2_X1 U989 ( .A1(n898), .A2(n897), .ZN(n899) );
  XOR2_X1 U990 ( .A(KEYINPUT53), .B(n899), .Z(n900) );
  XNOR2_X1 U991 ( .A(n900), .B(KEYINPUT120), .ZN(n901) );
  NAND2_X1 U992 ( .A1(n902), .A2(n901), .ZN(n905) );
  XNOR2_X1 U993 ( .A(G34), .B(G2084), .ZN(n903) );
  XNOR2_X1 U994 ( .A(KEYINPUT54), .B(n903), .ZN(n904) );
  NOR2_X1 U995 ( .A1(n905), .A2(n904), .ZN(n906) );
  XNOR2_X1 U996 ( .A(KEYINPUT121), .B(n906), .ZN(n907) );
  XNOR2_X1 U997 ( .A(n908), .B(n907), .ZN(n910) );
  INV_X1 U998 ( .A(G29), .ZN(n909) );
  NAND2_X1 U999 ( .A1(n910), .A2(n909), .ZN(n911) );
  NAND2_X1 U1000 ( .A1(G11), .A2(n911), .ZN(n964) );
  XNOR2_X1 U1001 ( .A(G16), .B(KEYINPUT56), .ZN(n932) );
  XNOR2_X1 U1002 ( .A(G1966), .B(G168), .ZN(n913) );
  NAND2_X1 U1003 ( .A1(n913), .A2(n912), .ZN(n914) );
  XNOR2_X1 U1004 ( .A(n914), .B(KEYINPUT57), .ZN(n930) );
  XNOR2_X1 U1005 ( .A(G1961), .B(G171), .ZN(n926) );
  XOR2_X1 U1006 ( .A(G299), .B(G1956), .Z(n916) );
  XNOR2_X1 U1007 ( .A(n1017), .B(G1348), .ZN(n915) );
  NAND2_X1 U1008 ( .A1(n916), .A2(n915), .ZN(n924) );
  XNOR2_X1 U1009 ( .A(G166), .B(G1971), .ZN(n918) );
  NAND2_X1 U1010 ( .A1(n918), .A2(n917), .ZN(n919) );
  NOR2_X1 U1011 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1012 ( .A1(n922), .A2(n921), .ZN(n923) );
  NOR2_X1 U1013 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1014 ( .A1(n926), .A2(n925), .ZN(n928) );
  XNOR2_X1 U1015 ( .A(G1341), .B(n1020), .ZN(n927) );
  NOR2_X1 U1016 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1017 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1018 ( .A1(n932), .A2(n931), .ZN(n962) );
  INV_X1 U1019 ( .A(G16), .ZN(n960) );
  XOR2_X1 U1020 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n945) );
  XOR2_X1 U1021 ( .A(G1341), .B(G19), .Z(n933) );
  XNOR2_X1 U1022 ( .A(KEYINPUT123), .B(n933), .ZN(n935) );
  XNOR2_X1 U1023 ( .A(G6), .B(G1981), .ZN(n934) );
  NOR2_X1 U1024 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1025 ( .A(n936), .B(KEYINPUT124), .ZN(n939) );
  XOR2_X1 U1026 ( .A(G1956), .B(KEYINPUT122), .Z(n937) );
  XNOR2_X1 U1027 ( .A(G20), .B(n937), .ZN(n938) );
  NAND2_X1 U1028 ( .A1(n939), .A2(n938), .ZN(n942) );
  XOR2_X1 U1029 ( .A(KEYINPUT59), .B(G1348), .Z(n940) );
  XNOR2_X1 U1030 ( .A(G4), .B(n940), .ZN(n941) );
  NOR2_X1 U1031 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1032 ( .A(n943), .B(KEYINPUT60), .ZN(n944) );
  XNOR2_X1 U1033 ( .A(n945), .B(n944), .ZN(n950) );
  XOR2_X1 U1034 ( .A(n946), .B(G5), .Z(n948) );
  XNOR2_X1 U1035 ( .A(G21), .B(G1966), .ZN(n947) );
  NOR2_X1 U1036 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1037 ( .A1(n950), .A2(n949), .ZN(n957) );
  XNOR2_X1 U1038 ( .A(G1971), .B(G22), .ZN(n952) );
  XNOR2_X1 U1039 ( .A(G24), .B(G1986), .ZN(n951) );
  NOR2_X1 U1040 ( .A1(n952), .A2(n951), .ZN(n954) );
  XOR2_X1 U1041 ( .A(G1976), .B(G23), .Z(n953) );
  NAND2_X1 U1042 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1043 ( .A(KEYINPUT58), .B(n955), .ZN(n956) );
  NOR2_X1 U1044 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1045 ( .A(KEYINPUT61), .B(n958), .ZN(n959) );
  NAND2_X1 U1046 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1047 ( .A1(n962), .A2(n961), .ZN(n963) );
  NOR2_X1 U1048 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1049 ( .A1(n966), .A2(n965), .ZN(n967) );
  XOR2_X1 U1050 ( .A(KEYINPUT62), .B(n967), .Z(G311) );
  XNOR2_X1 U1051 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1052 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1053 ( .A1(n969), .A2(n968), .ZN(G325) );
  INV_X1 U1054 ( .A(G325), .ZN(G261) );
  INV_X1 U1055 ( .A(n970), .ZN(G319) );
  XOR2_X1 U1056 ( .A(KEYINPUT112), .B(G2678), .Z(n972) );
  XNOR2_X1 U1057 ( .A(G2090), .B(G2072), .ZN(n971) );
  XNOR2_X1 U1058 ( .A(n972), .B(n971), .ZN(n976) );
  XOR2_X1 U1059 ( .A(KEYINPUT43), .B(KEYINPUT111), .Z(n974) );
  XNOR2_X1 U1060 ( .A(G2067), .B(KEYINPUT42), .ZN(n973) );
  XNOR2_X1 U1061 ( .A(n974), .B(n973), .ZN(n975) );
  XOR2_X1 U1062 ( .A(n976), .B(n975), .Z(n978) );
  XNOR2_X1 U1063 ( .A(G2096), .B(G2100), .ZN(n977) );
  XNOR2_X1 U1064 ( .A(n978), .B(n977), .ZN(n980) );
  XOR2_X1 U1065 ( .A(G2078), .B(G2084), .Z(n979) );
  XNOR2_X1 U1066 ( .A(n980), .B(n979), .ZN(G227) );
  XOR2_X1 U1067 ( .A(G1986), .B(G1976), .Z(n982) );
  XNOR2_X1 U1068 ( .A(G1966), .B(G1971), .ZN(n981) );
  XNOR2_X1 U1069 ( .A(n982), .B(n981), .ZN(n983) );
  XOR2_X1 U1070 ( .A(n983), .B(G2474), .Z(n985) );
  XNOR2_X1 U1071 ( .A(G1981), .B(G1991), .ZN(n984) );
  XNOR2_X1 U1072 ( .A(n985), .B(n984), .ZN(n989) );
  XOR2_X1 U1073 ( .A(KEYINPUT41), .B(G1996), .Z(n987) );
  XNOR2_X1 U1074 ( .A(G1961), .B(G1956), .ZN(n986) );
  XNOR2_X1 U1075 ( .A(n987), .B(n986), .ZN(n988) );
  XNOR2_X1 U1076 ( .A(n989), .B(n988), .ZN(G229) );
  NAND2_X1 U1077 ( .A1(G130), .A2(n990), .ZN(n993) );
  NAND2_X1 U1078 ( .A1(G118), .A2(n991), .ZN(n992) );
  NAND2_X1 U1079 ( .A1(n993), .A2(n992), .ZN(n999) );
  NAND2_X1 U1080 ( .A1(G106), .A2(n994), .ZN(n996) );
  NAND2_X1 U1081 ( .A1(G142), .A2(n724), .ZN(n995) );
  NAND2_X1 U1082 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1083 ( .A(KEYINPUT45), .B(n997), .Z(n998) );
  NOR2_X1 U1084 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1085 ( .A(G162), .B(n1000), .ZN(n1012) );
  XNOR2_X1 U1086 ( .A(G164), .B(n1001), .ZN(n1005) );
  XNOR2_X1 U1087 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n1003) );
  XNOR2_X1 U1088 ( .A(n1003), .B(n1002), .ZN(n1004) );
  XNOR2_X1 U1089 ( .A(n1005), .B(n1004), .ZN(n1007) );
  XOR2_X1 U1090 ( .A(n1007), .B(n1006), .Z(n1010) );
  XNOR2_X1 U1091 ( .A(G160), .B(n1008), .ZN(n1009) );
  XNOR2_X1 U1092 ( .A(n1010), .B(n1009), .ZN(n1011) );
  XNOR2_X1 U1093 ( .A(n1012), .B(n1011), .ZN(n1014) );
  XOR2_X1 U1094 ( .A(n1014), .B(n1013), .Z(n1015) );
  NOR2_X1 U1095 ( .A1(G37), .A2(n1015), .ZN(G395) );
  INV_X1 U1096 ( .A(G171), .ZN(G301) );
  XOR2_X1 U1097 ( .A(KEYINPUT116), .B(n1016), .Z(n1019) );
  XNOR2_X1 U1098 ( .A(G301), .B(n1017), .ZN(n1018) );
  XNOR2_X1 U1099 ( .A(n1019), .B(n1018), .ZN(n1022) );
  XNOR2_X1 U1100 ( .A(G286), .B(n1020), .ZN(n1021) );
  XNOR2_X1 U1101 ( .A(n1022), .B(n1021), .ZN(n1023) );
  NOR2_X1 U1102 ( .A1(G37), .A2(n1023), .ZN(G397) );
  XOR2_X1 U1103 ( .A(G2443), .B(G2454), .Z(n1025) );
  XNOR2_X1 U1104 ( .A(G1348), .B(G2435), .ZN(n1024) );
  XNOR2_X1 U1105 ( .A(n1025), .B(n1024), .ZN(n1032) );
  XOR2_X1 U1106 ( .A(KEYINPUT109), .B(G2446), .Z(n1027) );
  XNOR2_X1 U1107 ( .A(G1341), .B(G2430), .ZN(n1026) );
  XNOR2_X1 U1108 ( .A(n1027), .B(n1026), .ZN(n1028) );
  XOR2_X1 U1109 ( .A(n1028), .B(G2451), .Z(n1030) );
  XNOR2_X1 U1110 ( .A(G2438), .B(G2427), .ZN(n1029) );
  XNOR2_X1 U1111 ( .A(n1030), .B(n1029), .ZN(n1031) );
  XNOR2_X1 U1112 ( .A(n1032), .B(n1031), .ZN(n1033) );
  NAND2_X1 U1113 ( .A1(n1033), .A2(G14), .ZN(n1039) );
  NAND2_X1 U1114 ( .A1(G319), .A2(n1039), .ZN(n1036) );
  NOR2_X1 U1115 ( .A1(G227), .A2(G229), .ZN(n1034) );
  XNOR2_X1 U1116 ( .A(KEYINPUT49), .B(n1034), .ZN(n1035) );
  NOR2_X1 U1117 ( .A1(n1036), .A2(n1035), .ZN(n1038) );
  NOR2_X1 U1118 ( .A1(G395), .A2(G397), .ZN(n1037) );
  NAND2_X1 U1119 ( .A1(n1038), .A2(n1037), .ZN(G225) );
  INV_X1 U1120 ( .A(G225), .ZN(G308) );
  INV_X1 U1121 ( .A(G57), .ZN(G237) );
  INV_X1 U1122 ( .A(n1039), .ZN(G401) );
endmodule

