//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 0 1 0 1 0 1 0 1 0 1 0 1 0 0 0 1 0 1 1 1 1 0 0 1 1 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n794, new_n795, new_n797, new_n798, new_n799, new_n800, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n845, new_n846,
    new_n847, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913;
  XOR2_X1   g000(.A(G127gat), .B(G134gat), .Z(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT74), .B(KEYINPUT1), .ZN(new_n203));
  INV_X1    g002(.A(G113gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G120gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT72), .B(G120gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n205), .B1(new_n206), .B2(new_n204), .ZN(new_n207));
  AOI211_X1 g006(.A(new_n202), .B(new_n203), .C1(new_n207), .C2(KEYINPUT73), .ZN(new_n208));
  OR2_X1    g007(.A1(new_n207), .A2(KEYINPUT73), .ZN(new_n209));
  XNOR2_X1  g008(.A(G113gat), .B(G120gat), .ZN(new_n210));
  OR2_X1    g009(.A1(new_n210), .A2(KEYINPUT1), .ZN(new_n211));
  AOI22_X1  g010(.A1(new_n208), .A2(new_n209), .B1(new_n211), .B2(new_n202), .ZN(new_n212));
  AND2_X1   g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214));
  XOR2_X1   g013(.A(G141gat), .B(G148gat), .Z(new_n215));
  INV_X1    g014(.A(KEYINPUT2), .ZN(new_n216));
  AOI211_X1 g015(.A(new_n213), .B(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n213), .B1(new_n216), .B2(new_n214), .ZN(new_n218));
  XNOR2_X1  g017(.A(KEYINPUT81), .B(G148gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(G141gat), .ZN(new_n220));
  INV_X1    g019(.A(G141gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G148gat), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n218), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n217), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n212), .B(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(G225gat), .A2(G233gat), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n208), .A2(new_n209), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n211), .A2(new_n202), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n224), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT3), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT3), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n224), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n231), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  AND2_X1   g035(.A1(new_n236), .A2(KEYINPUT4), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n231), .A2(new_n232), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n224), .B(KEYINPUT82), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(new_n212), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT4), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n226), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  OAI211_X1 g042(.A(KEYINPUT5), .B(new_n228), .C1(new_n239), .C2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n236), .A2(KEYINPUT4), .ZN(new_n245));
  AOI22_X1  g044(.A1(new_n245), .A2(new_n241), .B1(KEYINPUT4), .B2(new_n238), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT5), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n246), .A2(new_n247), .A3(new_n226), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n244), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(G1gat), .B(G29gat), .ZN(new_n250));
  INV_X1    g049(.A(G85gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(KEYINPUT0), .B(G57gat), .ZN(new_n253));
  XOR2_X1   g052(.A(new_n252), .B(new_n253), .Z(new_n254));
  NAND2_X1  g053(.A1(new_n249), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT6), .ZN(new_n256));
  INV_X1    g055(.A(new_n254), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n244), .A2(new_n257), .A3(new_n248), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n255), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n249), .A2(KEYINPUT6), .A3(new_n254), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(KEYINPUT83), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT83), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n249), .A2(new_n262), .A3(KEYINPUT6), .A4(new_n254), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n259), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(KEYINPUT78), .B(G197gat), .ZN(new_n265));
  INV_X1    g064(.A(G204gat), .ZN(new_n266));
  OR2_X1    g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n265), .A2(new_n266), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT22), .ZN(new_n269));
  INV_X1    g068(.A(G211gat), .ZN(new_n270));
  INV_X1    g069(.A(G218gat), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n267), .A2(new_n268), .A3(new_n272), .ZN(new_n273));
  XOR2_X1   g072(.A(G211gat), .B(G218gat), .Z(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n275), .B(KEYINPUT79), .ZN(new_n276));
  NOR2_X1   g075(.A1(G169gat), .A2(G176gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(G169gat), .A2(G176gat), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n277), .B1(KEYINPUT23), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT25), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT66), .ZN(new_n282));
  INV_X1    g081(.A(G169gat), .ZN(new_n283));
  INV_X1    g082(.A(G176gat), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  OAI21_X1  g084(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT23), .ZN(new_n288));
  AND2_X1   g087(.A1(new_n281), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(G183gat), .A2(G190gat), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(KEYINPUT24), .B1(new_n291), .B2(KEYINPUT67), .ZN(new_n292));
  INV_X1    g091(.A(G183gat), .ZN(new_n293));
  INV_X1    g092(.A(G190gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT24), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n290), .A2(new_n296), .ZN(new_n297));
  OAI211_X1 g096(.A(new_n292), .B(new_n295), .C1(KEYINPUT67), .C2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n289), .A2(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n279), .B1(KEYINPUT23), .B2(new_n277), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n291), .A2(KEYINPUT65), .A3(KEYINPUT24), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT65), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n302), .B1(new_n290), .B2(new_n296), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n301), .A2(new_n297), .A3(new_n295), .A4(new_n303), .ZN(new_n304));
  AND2_X1   g103(.A1(new_n300), .A2(new_n304), .ZN(new_n305));
  XOR2_X1   g104(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n306));
  OAI21_X1  g105(.A(new_n299), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(KEYINPUT27), .B(G183gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n308), .A2(KEYINPUT28), .A3(new_n294), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  AND2_X1   g109(.A1(KEYINPUT68), .A2(KEYINPUT27), .ZN(new_n311));
  NOR2_X1   g110(.A1(KEYINPUT68), .A2(KEYINPUT27), .ZN(new_n312));
  OAI211_X1 g111(.A(KEYINPUT69), .B(G183gat), .C1(new_n311), .C2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT68), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT27), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(KEYINPUT68), .A2(KEYINPUT27), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n293), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(KEYINPUT69), .B1(new_n315), .B2(G183gat), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n313), .B(new_n294), .C1(new_n318), .C2(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT28), .B1(new_n321), .B2(KEYINPUT70), .ZN(new_n322));
  OAI21_X1  g121(.A(G183gat), .B1(new_n311), .B2(new_n312), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(new_n319), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT70), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n324), .A2(new_n325), .A3(new_n294), .A4(new_n313), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n310), .B1(new_n322), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n278), .ZN(new_n328));
  INV_X1    g127(.A(new_n277), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n328), .B1(new_n329), .B2(KEYINPUT26), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT26), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT71), .B1(new_n287), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT71), .ZN(new_n333));
  AOI211_X1 g132(.A(new_n333), .B(KEYINPUT26), .C1(new_n285), .C2(new_n286), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n330), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(new_n290), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n307), .B1(new_n327), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(G226gat), .ZN(new_n338));
  INV_X1    g137(.A(G233gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n340), .A2(KEYINPUT29), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n337), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n337), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT80), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT80), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n337), .A2(new_n345), .ZN(new_n346));
  AND2_X1   g145(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n340), .ZN(new_n348));
  OAI211_X1 g147(.A(new_n276), .B(new_n342), .C1(new_n347), .C2(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n344), .A2(new_n346), .A3(new_n341), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n343), .A2(new_n340), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n276), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n349), .A2(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(G8gat), .B(G36gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(G64gat), .B(G92gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n356), .B(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n358), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n349), .A2(new_n354), .A3(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n359), .A2(KEYINPUT30), .A3(new_n361), .ZN(new_n362));
  OR3_X1    g161(.A1(new_n355), .A2(KEYINPUT30), .A3(new_n358), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n264), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n235), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n276), .B1(KEYINPUT29), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(G228gat), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n368), .A2(new_n339), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT29), .ZN(new_n370));
  AOI21_X1  g169(.A(KEYINPUT3), .B1(new_n275), .B2(new_n370), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n367), .B(new_n369), .C1(new_n224), .C2(new_n371), .ZN(new_n372));
  OR3_X1    g171(.A1(new_n371), .A2(new_n240), .A3(KEYINPUT84), .ZN(new_n373));
  OAI21_X1  g172(.A(KEYINPUT84), .B1(new_n371), .B2(new_n240), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n367), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n369), .ZN(new_n376));
  AND3_X1   g175(.A1(new_n375), .A2(KEYINPUT85), .A3(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(KEYINPUT85), .B1(new_n375), .B2(new_n376), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n372), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  XOR2_X1   g178(.A(G78gat), .B(G106gat), .Z(new_n380));
  XNOR2_X1  g179(.A(new_n380), .B(G22gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(KEYINPUT31), .B(G50gat), .ZN(new_n382));
  XOR2_X1   g181(.A(new_n381), .B(new_n382), .Z(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n379), .A2(new_n384), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n372), .B(new_n383), .C1(new_n377), .C2(new_n378), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n365), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n321), .A2(KEYINPUT70), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT28), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n390), .A2(new_n326), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n336), .B1(new_n392), .B2(new_n309), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n306), .B1(new_n300), .B2(new_n304), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n394), .B1(new_n298), .B2(new_n289), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n231), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n307), .B(new_n212), .C1(new_n327), .C2(new_n336), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(G227gat), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n399), .A2(new_n339), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT75), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT75), .ZN(new_n402));
  INV_X1    g201(.A(new_n400), .ZN(new_n403));
  AOI211_X1 g202(.A(new_n402), .B(new_n403), .C1(new_n396), .C2(new_n397), .ZN(new_n404));
  OAI21_X1  g203(.A(KEYINPUT32), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT33), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n406), .B1(new_n401), .B2(new_n404), .ZN(new_n407));
  XNOR2_X1  g206(.A(G15gat), .B(G43gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(G71gat), .B(G99gat), .ZN(new_n409));
  XOR2_X1   g208(.A(new_n408), .B(new_n409), .Z(new_n410));
  NAND3_X1  g209(.A1(new_n405), .A2(new_n407), .A3(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n410), .ZN(new_n412));
  OAI221_X1 g211(.A(KEYINPUT32), .B1(new_n406), .B2(new_n412), .C1(new_n401), .C2(new_n404), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n396), .A2(new_n403), .A3(new_n397), .ZN(new_n415));
  XOR2_X1   g214(.A(new_n415), .B(KEYINPUT34), .Z(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n411), .A2(new_n416), .A3(new_n413), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n418), .A2(KEYINPUT36), .A3(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT76), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n418), .A2(KEYINPUT76), .A3(KEYINPUT36), .A4(new_n419), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT77), .ZN(new_n425));
  AND3_X1   g224(.A1(new_n411), .A2(new_n416), .A3(new_n413), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n416), .B1(new_n411), .B2(new_n413), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n425), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n419), .A2(KEYINPUT77), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT36), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n389), .B1(new_n424), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(KEYINPUT86), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT86), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n389), .B(new_n433), .C1(new_n424), .C2(new_n430), .ZN(new_n434));
  INV_X1    g233(.A(new_n355), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT37), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n360), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n437), .B1(new_n436), .B2(new_n435), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(KEYINPUT38), .ZN(new_n439));
  INV_X1    g238(.A(new_n264), .ZN(new_n440));
  INV_X1    g239(.A(new_n352), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n441), .A2(KEYINPUT88), .A3(new_n276), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n342), .B1(new_n347), .B2(new_n348), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(new_n353), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT88), .B1(new_n441), .B2(new_n276), .ZN(new_n446));
  OAI21_X1  g245(.A(KEYINPUT37), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT38), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n447), .A2(new_n437), .A3(new_n448), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n439), .A2(new_n440), .A3(new_n361), .A4(new_n449), .ZN(new_n450));
  OR3_X1    g249(.A1(new_n246), .A2(KEYINPUT39), .A3(new_n226), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n246), .A2(new_n226), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT39), .B1(new_n225), .B2(new_n227), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n451), .B(new_n257), .C1(new_n452), .C2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT87), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT40), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n255), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n459));
  OR3_X1    g258(.A1(new_n364), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n450), .A2(new_n387), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n432), .A2(new_n434), .A3(new_n461), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n426), .A2(new_n427), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n464), .A2(new_n388), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT35), .B1(new_n466), .B2(new_n365), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n428), .A2(new_n429), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n468), .A2(new_n388), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n364), .ZN(new_n470));
  OR2_X1    g269(.A1(new_n440), .A2(KEYINPUT35), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n467), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n462), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT89), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n462), .A2(new_n472), .A3(KEYINPUT89), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT94), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT15), .ZN(new_n478));
  AOI22_X1  g277(.A1(new_n477), .A2(new_n478), .B1(G43gat), .B2(G50gat), .ZN(new_n479));
  XNOR2_X1  g278(.A(KEYINPUT95), .B(G50gat), .ZN(new_n480));
  OAI221_X1 g279(.A(new_n479), .B1(new_n477), .B2(new_n478), .C1(new_n480), .C2(G43gat), .ZN(new_n481));
  AND2_X1   g280(.A1(G43gat), .A2(G50gat), .ZN(new_n482));
  NOR2_X1   g281(.A1(G43gat), .A2(G50gat), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT15), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(G29gat), .A2(G36gat), .ZN(new_n485));
  OR3_X1    g284(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n486));
  OAI21_X1  g285(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n481), .A2(new_n484), .A3(new_n485), .A4(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n489), .B(KEYINPUT96), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n486), .A2(KEYINPUT93), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n487), .B1(new_n486), .B2(KEYINPUT93), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n485), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n484), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n496), .B(KEYINPUT97), .ZN(new_n497));
  XNOR2_X1  g296(.A(G15gat), .B(G22gat), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n498), .A2(G1gat), .ZN(new_n499));
  INV_X1    g298(.A(G1gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT16), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n501), .B(KEYINPUT98), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n499), .B1(new_n502), .B2(new_n498), .ZN(new_n503));
  XOR2_X1   g302(.A(KEYINPUT100), .B(G8gat), .Z(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT99), .ZN(new_n506));
  AOI211_X1 g305(.A(new_n506), .B(new_n499), .C1(new_n498), .C2(new_n502), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n502), .A2(new_n506), .A3(new_n498), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(G8gat), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n505), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(KEYINPUT101), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(KEYINPUT102), .B1(new_n497), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n512), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n513), .B(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(G229gat), .A2(G233gat), .ZN(new_n516));
  XOR2_X1   g315(.A(new_n516), .B(KEYINPUT13), .Z(new_n517));
  INV_X1    g316(.A(KEYINPUT17), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n497), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n510), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n490), .A2(KEYINPUT17), .A3(new_n495), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n522), .A2(new_n516), .A3(new_n514), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT18), .ZN(new_n524));
  AOI22_X1  g323(.A1(new_n515), .A2(new_n517), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G169gat), .B(G197gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n526), .B(new_n221), .ZN(new_n527));
  XNOR2_X1  g326(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(KEYINPUT91), .B(G113gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  XOR2_X1   g330(.A(KEYINPUT92), .B(KEYINPUT12), .Z(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  AND2_X1   g332(.A1(new_n522), .A2(new_n514), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n534), .A2(KEYINPUT18), .A3(new_n516), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n525), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n533), .B1(new_n525), .B2(new_n535), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n475), .A2(new_n476), .A3(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT9), .ZN(new_n542));
  INV_X1    g341(.A(G71gat), .ZN(new_n543));
  INV_X1    g342(.A(G78gat), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT103), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n545), .A2(new_n546), .ZN(new_n548));
  XOR2_X1   g347(.A(G57gat), .B(G64gat), .Z(new_n549));
  NAND3_X1  g348(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  XOR2_X1   g349(.A(G71gat), .B(G78gat), .Z(new_n551));
  OR2_X1    g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n551), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT21), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  XOR2_X1   g355(.A(new_n556), .B(KEYINPUT104), .Z(new_n557));
  OAI21_X1  g356(.A(new_n511), .B1(new_n555), .B2(new_n554), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(KEYINPUT105), .B(KEYINPUT106), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(G231gat), .A2(G233gat), .ZN(new_n562));
  INV_X1    g361(.A(G127gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(G155gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n561), .B(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G183gat), .B(G211gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  OR2_X1    g368(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n566), .A2(new_n569), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(G92gat), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n251), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(KEYINPUT108), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT108), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n576), .B1(new_n251), .B2(new_n573), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n575), .A2(KEYINPUT7), .A3(new_n577), .ZN(new_n578));
  OR3_X1    g377(.A1(new_n574), .A2(KEYINPUT108), .A3(KEYINPUT7), .ZN(new_n579));
  NAND2_X1  g378(.A1(G99gat), .A2(G106gat), .ZN(new_n580));
  AOI22_X1  g379(.A1(KEYINPUT8), .A2(new_n580), .B1(new_n251), .B2(new_n573), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n578), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G99gat), .B(G106gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT109), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n578), .A2(new_n579), .A3(new_n583), .A4(new_n581), .ZN(new_n587));
  AND2_X1   g386(.A1(new_n587), .A2(new_n585), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n519), .A2(new_n521), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G232gat), .A2(G233gat), .ZN(new_n592));
  XOR2_X1   g391(.A(new_n592), .B(KEYINPUT107), .Z(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  AOI22_X1  g393(.A1(new_n497), .A2(new_n589), .B1(KEYINPUT41), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  XOR2_X1   g395(.A(G134gat), .B(G162gat), .Z(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n594), .A2(KEYINPUT41), .ZN(new_n599));
  XNOR2_X1  g398(.A(G190gat), .B(G218gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n598), .A2(new_n602), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n572), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(G120gat), .B(G148gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(G176gat), .B(G204gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n589), .A2(new_n554), .ZN(new_n611));
  OR2_X1    g410(.A1(new_n584), .A2(new_n554), .ZN(new_n612));
  AOI21_X1  g411(.A(KEYINPUT10), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n589), .A2(KEYINPUT10), .A3(new_n553), .A4(new_n552), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  OR2_X1    g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(G230gat), .A2(G233gat), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n617), .B(KEYINPUT110), .Z(new_n618));
  AND2_X1   g417(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n611), .A2(new_n612), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n620), .A2(new_n617), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n610), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n621), .A2(new_n610), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n617), .B1(new_n613), .B2(new_n615), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n541), .A2(new_n607), .A3(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n628), .A2(new_n264), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(new_n500), .ZN(G1324gat));
  INV_X1    g429(.A(new_n364), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n541), .A2(new_n631), .A3(new_n607), .A4(new_n627), .ZN(new_n632));
  XOR2_X1   g431(.A(KEYINPUT16), .B(G8gat), .Z(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NOR3_X1   g433(.A1(new_n632), .A2(KEYINPUT42), .A3(new_n634), .ZN(new_n635));
  OR2_X1    g434(.A1(new_n632), .A2(new_n634), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT42), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n637), .B1(new_n632), .B2(G8gat), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n635), .B1(new_n636), .B2(new_n638), .ZN(G1325gat));
  INV_X1    g438(.A(new_n628), .ZN(new_n640));
  INV_X1    g439(.A(new_n424), .ZN(new_n641));
  INV_X1    g440(.A(new_n430), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  AND3_X1   g443(.A1(new_n640), .A2(G15gat), .A3(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n468), .ZN(new_n646));
  AOI21_X1  g445(.A(G15gat), .B1(new_n640), .B2(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n645), .A2(new_n647), .ZN(G1326gat));
  NOR2_X1   g447(.A1(new_n628), .A2(new_n387), .ZN(new_n649));
  XOR2_X1   g448(.A(KEYINPUT43), .B(G22gat), .Z(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(G1327gat));
  AND2_X1   g450(.A1(new_n570), .A2(new_n571), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n652), .A2(new_n605), .A3(new_n626), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n541), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n264), .A2(G29gat), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(KEYINPUT111), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT111), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n541), .A2(new_n658), .A3(new_n653), .A4(new_n655), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT45), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AND2_X1   g461(.A1(new_n606), .A2(KEYINPUT44), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n475), .A2(new_n476), .A3(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n461), .A2(new_n643), .A3(new_n389), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n605), .B1(new_n472), .B2(new_n665), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n666), .A2(KEYINPUT44), .ZN(new_n667));
  AND2_X1   g466(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT113), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n572), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n570), .A2(KEYINPUT113), .A3(new_n571), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(KEYINPUT112), .B1(new_n537), .B2(new_n538), .ZN(new_n674));
  INV_X1    g473(.A(new_n538), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT112), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n675), .A2(new_n676), .A3(new_n536), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n673), .A2(new_n626), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n668), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(G29gat), .B1(new_n680), .B2(new_n264), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n657), .A2(new_n659), .A3(KEYINPUT45), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n662), .A2(new_n681), .A3(new_n682), .ZN(G1328gat));
  OAI21_X1  g482(.A(G36gat), .B1(new_n680), .B2(new_n364), .ZN(new_n684));
  OR2_X1    g483(.A1(new_n364), .A2(G36gat), .ZN(new_n685));
  OAI21_X1  g484(.A(KEYINPUT46), .B1(new_n654), .B2(new_n685), .ZN(new_n686));
  OR3_X1    g485(.A1(new_n654), .A2(KEYINPUT46), .A3(new_n685), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n684), .A2(new_n686), .A3(new_n687), .ZN(G1329gat));
  NAND4_X1  g487(.A1(new_n664), .A2(new_n644), .A3(new_n667), .A4(new_n679), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(G43gat), .ZN(new_n690));
  INV_X1    g489(.A(G43gat), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n646), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n690), .B1(new_n654), .B2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT47), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(G1330gat));
  NAND4_X1  g494(.A1(new_n664), .A2(new_n388), .A3(new_n667), .A4(new_n679), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(new_n480), .ZN(new_n697));
  OR2_X1    g496(.A1(new_n387), .A2(new_n480), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n697), .B1(new_n654), .B2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT48), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(G1331gat));
  NAND2_X1  g500(.A1(new_n652), .A2(new_n605), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n702), .A2(new_n627), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(new_n678), .ZN(new_n704));
  OR2_X1    g503(.A1(new_n704), .A2(KEYINPUT114), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(KEYINPUT114), .ZN(new_n706));
  AOI22_X1  g505(.A1(new_n705), .A2(new_n706), .B1(new_n472), .B2(new_n665), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(new_n440), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g508(.A1(new_n705), .A2(new_n706), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n472), .A2(new_n665), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n712), .A2(new_n364), .ZN(new_n713));
  NOR2_X1   g512(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n714));
  AND2_X1   g513(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n716), .B1(new_n713), .B2(new_n714), .ZN(G1333gat));
  OAI21_X1  g516(.A(new_n543), .B1(new_n712), .B2(new_n468), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT50), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n644), .A2(G71gat), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n718), .B(new_n719), .C1(new_n712), .C2(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n712), .A2(new_n720), .ZN(new_n722));
  AOI21_X1  g521(.A(G71gat), .B1(new_n707), .B2(new_n646), .ZN(new_n723));
  OAI21_X1  g522(.A(KEYINPUT50), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n721), .A2(new_n724), .ZN(G1334gat));
  NAND2_X1  g524(.A1(new_n707), .A2(new_n388), .ZN(new_n726));
  XNOR2_X1  g525(.A(KEYINPUT115), .B(G78gat), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(G1335gat));
  INV_X1    g527(.A(new_n678), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n729), .A2(new_n652), .A3(new_n627), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n668), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(G85gat), .B1(new_n731), .B2(new_n264), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n666), .A2(new_n572), .A3(new_n678), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT51), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n440), .A2(new_n251), .A3(new_n626), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n732), .B1(new_n734), .B2(new_n735), .ZN(G1336gat));
  NAND4_X1  g535(.A1(new_n664), .A2(new_n631), .A3(new_n667), .A4(new_n730), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(G92gat), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT52), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n627), .A2(new_n364), .A3(G92gat), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n738), .B(new_n739), .C1(new_n734), .C2(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(KEYINPUT116), .A2(KEYINPUT51), .ZN(new_n743));
  OR2_X1    g542(.A1(new_n733), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n733), .A2(new_n743), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n741), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n746), .B1(G92gat), .B2(new_n737), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n742), .B1(new_n747), .B2(new_n739), .ZN(G1337gat));
  OAI21_X1  g547(.A(G99gat), .B1(new_n731), .B2(new_n643), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n468), .A2(new_n627), .A3(G99gat), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT117), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n749), .B1(new_n734), .B2(new_n751), .ZN(G1338gat));
  NAND4_X1  g551(.A1(new_n664), .A2(new_n388), .A3(new_n667), .A4(new_n730), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(G106gat), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT53), .ZN(new_n755));
  OR3_X1    g554(.A1(new_n627), .A2(new_n387), .A3(G106gat), .ZN(new_n756));
  OAI211_X1 g555(.A(new_n754), .B(new_n755), .C1(new_n734), .C2(new_n756), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n753), .A2(KEYINPUT118), .A3(G106gat), .ZN(new_n758));
  AOI21_X1  g557(.A(KEYINPUT118), .B1(new_n753), .B2(G106gat), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n756), .B1(new_n744), .B2(new_n745), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n757), .B1(new_n761), .B2(new_n755), .ZN(G1339gat));
  OAI211_X1 g561(.A(KEYINPUT54), .B(new_n624), .C1(new_n616), .C2(new_n618), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT54), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n616), .A2(new_n764), .A3(new_n618), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n763), .A2(KEYINPUT55), .A3(new_n610), .A4(new_n765), .ZN(new_n766));
  AND3_X1   g565(.A1(new_n766), .A2(KEYINPUT119), .A3(new_n625), .ZN(new_n767));
  AOI21_X1  g566(.A(KEYINPUT119), .B1(new_n766), .B2(new_n625), .ZN(new_n768));
  AND2_X1   g567(.A1(new_n765), .A2(new_n610), .ZN(new_n769));
  AOI21_X1  g568(.A(KEYINPUT55), .B1(new_n769), .B2(new_n763), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n767), .A2(new_n768), .A3(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n674), .A2(new_n677), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n515), .A2(new_n517), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n534), .A2(new_n516), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n531), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n536), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(new_n626), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n606), .B1(new_n772), .B2(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n606), .A2(new_n771), .A3(new_n776), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n672), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n607), .A2(new_n627), .A3(new_n678), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n264), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n466), .A2(new_n631), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n786), .A2(new_n204), .A3(new_n729), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n783), .A2(new_n364), .A3(new_n469), .ZN(new_n788));
  OAI21_X1  g587(.A(G113gat), .B1(new_n788), .B2(new_n539), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n787), .A2(new_n789), .ZN(G1340gat));
  OAI21_X1  g589(.A(G120gat), .B1(new_n788), .B2(new_n627), .ZN(new_n791));
  OR2_X1    g590(.A1(new_n627), .A2(new_n206), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n791), .B1(new_n785), .B2(new_n792), .ZN(G1341gat));
  AOI21_X1  g592(.A(G127gat), .B1(new_n786), .B2(new_n652), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n788), .A2(new_n563), .A3(new_n672), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n794), .A2(new_n795), .ZN(G1342gat));
  OR3_X1    g595(.A1(new_n785), .A2(G134gat), .A3(new_n605), .ZN(new_n797));
  OR2_X1    g596(.A1(new_n797), .A2(KEYINPUT56), .ZN(new_n798));
  OAI21_X1  g597(.A(G134gat), .B1(new_n788), .B2(new_n605), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(KEYINPUT56), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(G1343gat));
  NAND2_X1  g600(.A1(new_n781), .A2(new_n782), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n388), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n643), .A2(new_n440), .A3(new_n364), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n805), .A2(new_n221), .A3(new_n540), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT58), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT57), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n387), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n766), .A2(new_n625), .ZN(new_n811));
  XOR2_X1   g610(.A(KEYINPUT120), .B(KEYINPUT55), .Z(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n813), .B1(new_n769), .B2(new_n763), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n539), .A2(new_n811), .A3(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(new_n777), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n605), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n652), .B1(new_n817), .B2(new_n779), .ZN(new_n818));
  INV_X1    g617(.A(new_n782), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n810), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n387), .B1(new_n781), .B2(new_n782), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n820), .B1(new_n821), .B2(KEYINPUT57), .ZN(new_n822));
  INV_X1    g621(.A(new_n804), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n822), .A2(new_n540), .A3(new_n823), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n824), .A2(KEYINPUT121), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT121), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n822), .A2(new_n826), .A3(new_n540), .A4(new_n823), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(G141gat), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n808), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n822), .A2(new_n729), .A3(new_n823), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(G141gat), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n806), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(KEYINPUT58), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n829), .A2(new_n833), .ZN(G1344gat));
  NAND3_X1  g633(.A1(new_n805), .A2(new_n219), .A3(new_n626), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n822), .A2(new_n823), .ZN(new_n836));
  AOI211_X1 g635(.A(KEYINPUT59), .B(new_n219), .C1(new_n836), .C2(new_n626), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT59), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n803), .A2(KEYINPUT57), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n702), .A2(new_n540), .A3(new_n626), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n809), .B(new_n388), .C1(new_n818), .C2(new_n840), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n839), .A2(new_n626), .A3(new_n823), .A4(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n838), .B1(new_n842), .B2(G148gat), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n835), .B1(new_n837), .B2(new_n843), .ZN(G1345gat));
  AOI21_X1  g643(.A(G155gat), .B1(new_n805), .B2(new_n652), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n673), .A2(G155gat), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n846), .B(KEYINPUT122), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n845), .B1(new_n836), .B2(new_n847), .ZN(G1346gat));
  AOI21_X1  g647(.A(G162gat), .B1(new_n805), .B2(new_n606), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n606), .A2(G162gat), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n849), .B1(new_n836), .B2(new_n850), .ZN(G1347gat));
  NOR2_X1   g650(.A1(new_n440), .A2(new_n364), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n802), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n469), .ZN(new_n854));
  OAI21_X1  g653(.A(G169gat), .B1(new_n854), .B2(new_n539), .ZN(new_n855));
  AND3_X1   g654(.A1(new_n802), .A2(new_n465), .A3(new_n852), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n856), .A2(new_n283), .A3(new_n729), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n855), .A2(new_n857), .ZN(G1348gat));
  OAI21_X1  g657(.A(G176gat), .B1(new_n854), .B2(new_n627), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n856), .A2(new_n284), .A3(new_n626), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(KEYINPUT123), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT123), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n859), .A2(new_n863), .A3(new_n860), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n862), .A2(new_n864), .ZN(G1349gat));
  INV_X1    g664(.A(KEYINPUT124), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n866), .A2(KEYINPUT60), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n856), .A2(new_n308), .A3(new_n652), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n802), .A2(new_n469), .A3(new_n673), .A4(new_n852), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(G183gat), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n867), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n866), .A2(KEYINPUT60), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n871), .B(new_n872), .ZN(G1350gat));
  NAND3_X1  g672(.A1(new_n853), .A2(new_n469), .A3(new_n606), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT61), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n874), .A2(new_n875), .A3(G190gat), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(KEYINPUT125), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n874), .A2(G190gat), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(KEYINPUT61), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT125), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n874), .A2(new_n880), .A3(new_n875), .A4(G190gat), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n877), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n856), .A2(new_n294), .A3(new_n606), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(G1351gat));
  NAND2_X1  g683(.A1(new_n643), .A2(new_n852), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n841), .B(new_n886), .C1(new_n821), .C2(new_n809), .ZN(new_n887));
  OAI21_X1  g686(.A(G197gat), .B1(new_n887), .B2(new_n539), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n803), .A2(new_n885), .ZN(new_n889));
  INV_X1    g688(.A(G197gat), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n889), .A2(new_n890), .A3(new_n729), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n888), .A2(new_n891), .ZN(G1352gat));
  INV_X1    g691(.A(KEYINPUT127), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n627), .A2(G204gat), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n821), .A2(new_n886), .A3(new_n894), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(KEYINPUT126), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n893), .B1(new_n896), .B2(KEYINPUT62), .ZN(new_n897));
  OR2_X1    g696(.A1(new_n895), .A2(KEYINPUT126), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT62), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n895), .A2(KEYINPUT126), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n898), .A2(KEYINPUT127), .A3(new_n899), .A4(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n896), .A2(KEYINPUT62), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n839), .A2(new_n626), .A3(new_n841), .ZN(new_n903));
  OAI21_X1  g702(.A(G204gat), .B1(new_n903), .B2(new_n885), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n897), .A2(new_n901), .A3(new_n902), .A4(new_n904), .ZN(G1353gat));
  NAND3_X1  g704(.A1(new_n889), .A2(new_n270), .A3(new_n652), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n887), .A2(new_n572), .ZN(new_n907));
  AOI21_X1  g706(.A(KEYINPUT63), .B1(new_n907), .B2(G211gat), .ZN(new_n908));
  OAI211_X1 g707(.A(KEYINPUT63), .B(G211gat), .C1(new_n887), .C2(new_n572), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n906), .B1(new_n908), .B2(new_n910), .ZN(G1354gat));
  NOR3_X1   g710(.A1(new_n887), .A2(new_n271), .A3(new_n605), .ZN(new_n912));
  AOI21_X1  g711(.A(G218gat), .B1(new_n889), .B2(new_n606), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n912), .A2(new_n913), .ZN(G1355gat));
endmodule


