//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 1 0 1 0 0 0 1 0 0 1 0 0 0 0 1 0 0 0 0 1 1 0 1 0 1 1 0 1 0 1 1 0 1 1 0 0 0 0 0 0 0 1 1 0 1 0 0 1 0 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:26 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G353));
  NOR2_X1   g0005(.A1(G97), .A2(G107), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT65), .Z(G355));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT0), .ZN(new_n216));
  OAI21_X1  g0016(.A(G50), .B1(G58), .B2(G68), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(new_n211), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  AND2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OR2_X1    g0024(.A1(new_n224), .A2(KEYINPUT66), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(KEYINPUT66), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n228));
  NAND4_X1  g0028(.A1(new_n225), .A2(new_n226), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(new_n213), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n216), .B(new_n221), .C1(new_n230), .C2(KEYINPUT1), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XOR2_X1   g0032(.A(G226), .B(G232), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT68), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT69), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n234), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n202), .A2(G68), .ZN(new_n247));
  INV_X1    g0047(.A(G68), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G50), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G58), .B(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n246), .B(new_n252), .ZN(G351));
  INV_X1    g0053(.A(KEYINPUT75), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G41), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(G1), .A3(G13), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n210), .B1(G41), .B2(G45), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n256), .A2(KEYINPUT70), .A3(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  AOI21_X1  g0059(.A(KEYINPUT70), .B1(new_n256), .B2(new_n257), .ZN(new_n260));
  OAI21_X1  g0060(.A(G238), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT3), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G33), .ZN(new_n265));
  NAND4_X1  g0065(.A1(new_n263), .A2(new_n265), .A3(G232), .A4(G1698), .ZN(new_n266));
  INV_X1    g0066(.A(G1698), .ZN(new_n267));
  NAND4_X1  g0067(.A1(new_n263), .A2(new_n265), .A3(G226), .A4(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G97), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n266), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n219), .B1(G33), .B2(G41), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G41), .ZN(new_n273));
  INV_X1    g0073(.A(G45), .ZN(new_n274));
  AOI21_X1  g0074(.A(G1), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n275), .A2(new_n256), .A3(G274), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT74), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n275), .A2(new_n256), .A3(KEYINPUT74), .A4(G274), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n261), .A2(new_n272), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(KEYINPUT13), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT13), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n261), .A2(new_n272), .A3(new_n280), .A4(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n282), .A2(G190), .A3(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n210), .A2(G13), .A3(G20), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n248), .ZN(new_n288));
  XNOR2_X1  g0088(.A(new_n288), .B(KEYINPUT12), .ZN(new_n289));
  NOR2_X1   g0089(.A1(G20), .A2(G33), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n290), .A2(G50), .B1(G20), .B2(new_n248), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n262), .A2(G20), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G77), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n291), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n219), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n295), .A2(KEYINPUT11), .A3(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n287), .A2(new_n297), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n210), .A2(G20), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n299), .A2(G68), .A3(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n289), .A2(new_n298), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(KEYINPUT11), .B1(new_n295), .B2(new_n297), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n285), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G200), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n306), .B1(new_n282), .B2(new_n284), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n254), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n282), .A2(new_n284), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G200), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n310), .A2(KEYINPUT75), .A3(new_n304), .A4(new_n285), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G226), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n256), .A2(new_n257), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT70), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n313), .B1(new_n316), .B2(new_n258), .ZN(new_n317));
  INV_X1    g0117(.A(new_n276), .ZN(new_n318));
  OAI21_X1  g0118(.A(KEYINPUT71), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(G226), .B1(new_n259), .B2(new_n260), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT71), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n320), .A2(new_n321), .A3(new_n276), .ZN(new_n322));
  XNOR2_X1  g0122(.A(KEYINPUT3), .B(G33), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n323), .A2(G222), .A3(new_n267), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n323), .A2(G223), .A3(G1698), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n324), .B(new_n325), .C1(new_n294), .C2(new_n323), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n271), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n319), .A2(new_n322), .A3(new_n327), .ZN(new_n328));
  XNOR2_X1  g0128(.A(KEYINPUT73), .B(G200), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n297), .ZN(new_n331));
  INV_X1    g0131(.A(G58), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT8), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT8), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G58), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n336), .A2(new_n292), .B1(G150), .B2(new_n290), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n203), .A2(G20), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n331), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n331), .A2(new_n286), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n300), .A2(G50), .ZN(new_n342));
  OAI22_X1  g0142(.A1(new_n341), .A2(new_n342), .B1(G50), .B2(new_n286), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(KEYINPUT9), .B1(new_n340), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT9), .ZN(new_n346));
  NOR3_X1   g0146(.A1(new_n339), .A2(new_n343), .A3(new_n346), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n319), .A2(new_n322), .A3(G190), .A4(new_n327), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n330), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(KEYINPUT10), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT10), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n330), .A2(new_n348), .A3(new_n352), .A4(new_n349), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n304), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT14), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n316), .A2(new_n258), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n357), .A2(G238), .B1(new_n278), .B2(new_n279), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n283), .B1(new_n358), .B2(new_n272), .ZN(new_n359));
  AND4_X1   g0159(.A1(new_n283), .A2(new_n261), .A3(new_n272), .A4(new_n280), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n356), .B(G169), .C1(new_n359), .C2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n282), .A2(G179), .A3(new_n284), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n356), .B1(new_n309), .B2(G169), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n355), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n312), .A2(new_n354), .A3(new_n365), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n263), .A2(new_n265), .A3(G232), .A4(new_n267), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n263), .A2(new_n265), .A3(G238), .A4(G1698), .ZN(new_n368));
  INV_X1    g0168(.A(G107), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n367), .B(new_n368), .C1(new_n369), .C2(new_n323), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n271), .ZN(new_n371));
  OAI21_X1  g0171(.A(G244), .B1(new_n259), .B2(new_n260), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n371), .A2(new_n372), .A3(new_n276), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n329), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n318), .B1(new_n357), .B2(G244), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n375), .A2(G190), .A3(new_n371), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT72), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n336), .A2(new_n290), .B1(G20), .B2(G77), .ZN(new_n378));
  XOR2_X1   g0178(.A(KEYINPUT15), .B(G87), .Z(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n292), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n331), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n300), .A2(G77), .ZN(new_n382));
  OAI22_X1  g0182(.A1(new_n341), .A2(new_n382), .B1(G77), .B2(new_n286), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n377), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  XNOR2_X1  g0184(.A(KEYINPUT8), .B(G58), .ZN(new_n385));
  INV_X1    g0185(.A(new_n290), .ZN(new_n386));
  OAI22_X1  g0186(.A1(new_n385), .A2(new_n386), .B1(new_n211), .B2(new_n294), .ZN(new_n387));
  XNOR2_X1  g0187(.A(KEYINPUT15), .B(G87), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n388), .A2(new_n293), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n297), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n382), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n299), .A2(new_n391), .B1(new_n294), .B2(new_n287), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n390), .A2(KEYINPUT72), .A3(new_n392), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n374), .A2(new_n376), .A3(new_n384), .A4(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n384), .A2(new_n393), .ZN(new_n395));
  INV_X1    g0195(.A(G169), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n373), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(G179), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n375), .A2(new_n398), .A3(new_n371), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n395), .A2(new_n397), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n394), .A2(new_n400), .ZN(new_n401));
  OR2_X1    g0201(.A1(new_n328), .A2(G179), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n339), .A2(new_n343), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n403), .B1(new_n328), .B2(new_n396), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n401), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(G223), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n406), .A2(G1698), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n407), .A2(new_n263), .A3(new_n265), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(KEYINPUT76), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n323), .A2(G226), .A3(G1698), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT76), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n323), .A2(new_n411), .A3(new_n407), .ZN(new_n412));
  NAND2_X1  g0212(.A1(G33), .A2(G87), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n409), .A2(new_n410), .A3(new_n412), .A4(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n271), .ZN(new_n415));
  INV_X1    g0215(.A(G190), .ZN(new_n416));
  INV_X1    g0216(.A(G232), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n276), .B1(new_n314), .B2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n415), .A2(new_n416), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n418), .B1(new_n414), .B2(new_n271), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n420), .B1(G200), .B2(new_n421), .ZN(new_n422));
  AND2_X1   g0222(.A1(new_n336), .A2(new_n300), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n423), .A2(new_n299), .B1(new_n287), .B2(new_n385), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT7), .ZN(new_n426));
  NOR3_X1   g0226(.A1(new_n323), .A2(new_n426), .A3(G20), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n263), .A2(new_n265), .ZN(new_n428));
  AOI21_X1  g0228(.A(KEYINPUT7), .B1(new_n428), .B2(new_n211), .ZN(new_n429));
  OAI21_X1  g0229(.A(G68), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n332), .A2(new_n248), .ZN(new_n431));
  OAI21_X1  g0231(.A(G20), .B1(new_n431), .B2(new_n201), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n290), .A2(G159), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n432), .A2(KEYINPUT16), .A3(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n331), .B1(new_n430), .B2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT16), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n426), .B1(new_n323), .B2(G20), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n428), .A2(KEYINPUT7), .A3(new_n211), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n248), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n432), .A2(new_n433), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n437), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n425), .B1(new_n436), .B2(new_n442), .ZN(new_n443));
  AND3_X1   g0243(.A1(new_n422), .A2(KEYINPUT17), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(KEYINPUT17), .B1(new_n422), .B2(new_n443), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n441), .ZN(new_n447));
  AOI21_X1  g0247(.A(KEYINPUT16), .B1(new_n430), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n297), .B1(new_n440), .B2(new_n434), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n424), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  OR2_X1    g0250(.A1(new_n421), .A2(G169), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT77), .ZN(new_n452));
  AND4_X1   g0252(.A1(new_n452), .A2(new_n415), .A3(new_n398), .A4(new_n419), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n452), .B1(new_n421), .B2(new_n398), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n450), .B(new_n451), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(KEYINPUT18), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n415), .A2(new_n398), .A3(new_n419), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(KEYINPUT77), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n421), .A2(new_n452), .A3(new_n398), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT18), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n460), .A2(new_n461), .A3(new_n450), .A4(new_n451), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n405), .A2(new_n446), .A3(new_n456), .A4(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n366), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n274), .A2(G1), .ZN(new_n465));
  AND2_X1   g0265(.A1(KEYINPUT5), .A2(G41), .ZN(new_n466));
  NOR2_X1   g0266(.A1(KEYINPUT5), .A2(G41), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n468), .A2(G270), .A3(new_n256), .ZN(new_n469));
  XNOR2_X1  g0269(.A(KEYINPUT5), .B(G41), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n470), .A2(new_n256), .A3(G274), .A4(new_n465), .ZN(new_n471));
  AND2_X1   g0271(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n264), .A2(G33), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n474));
  OAI21_X1  g0274(.A(G303), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n263), .A2(new_n265), .A3(G264), .A4(G1698), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n263), .A2(new_n265), .A3(G257), .A4(new_n267), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n271), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n472), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n210), .A2(G33), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n286), .A2(new_n481), .A3(new_n219), .A4(new_n296), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(G116), .ZN(new_n484));
  INV_X1    g0284(.A(G116), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n287), .A2(new_n485), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n296), .A2(new_n219), .B1(G20), .B2(new_n485), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G283), .ZN(new_n488));
  INV_X1    g0288(.A(G97), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n488), .B(new_n211), .C1(G33), .C2(new_n489), .ZN(new_n490));
  AND3_X1   g0290(.A1(new_n487), .A2(KEYINPUT20), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(KEYINPUT20), .B1(new_n487), .B2(new_n490), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n484), .B(new_n486), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n480), .A2(G169), .A3(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT21), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AND3_X1   g0296(.A1(new_n472), .A2(G179), .A3(new_n479), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n493), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n472), .A2(new_n479), .A3(G190), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n491), .A2(new_n492), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n486), .B1(new_n482), .B2(new_n485), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n469), .A2(new_n471), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n503), .B1(new_n271), .B2(new_n478), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n499), .B(new_n502), .C1(new_n504), .C2(new_n306), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n480), .A2(new_n493), .A3(KEYINPUT21), .A4(G169), .ZN(new_n506));
  AND4_X1   g0306(.A1(new_n496), .A2(new_n498), .A3(new_n505), .A4(new_n506), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n263), .A2(new_n265), .A3(new_n211), .A4(G87), .ZN(new_n508));
  XNOR2_X1  g0308(.A(KEYINPUT82), .B(KEYINPUT22), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT22), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n511), .A2(KEYINPUT82), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n323), .A2(new_n211), .A3(G87), .A4(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(G33), .A2(G116), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n514), .A2(G20), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT23), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(new_n211), .B2(G107), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n369), .A2(KEYINPUT23), .A3(G20), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n515), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n510), .A2(new_n513), .A3(new_n519), .ZN(new_n520));
  XOR2_X1   g0320(.A(KEYINPUT83), .B(KEYINPUT24), .Z(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n521), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n510), .A2(new_n513), .A3(new_n519), .A4(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n297), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n287), .A2(KEYINPUT25), .A3(new_n369), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT25), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n528), .B1(new_n286), .B2(G107), .ZN(new_n529));
  AOI22_X1  g0329(.A1(G107), .A2(new_n483), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n263), .A2(new_n265), .A3(G257), .A4(G1698), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n263), .A2(new_n265), .A3(G250), .A4(new_n267), .ZN(new_n532));
  NAND2_X1  g0332(.A1(G33), .A2(G294), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n271), .B1(new_n465), .B2(new_n470), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n534), .A2(new_n271), .B1(new_n535), .B2(G264), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n536), .A2(G190), .A3(new_n471), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n534), .A2(new_n271), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n535), .A2(G264), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n538), .A2(new_n539), .A3(new_n471), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(G200), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n526), .A2(new_n530), .A3(new_n537), .A4(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n379), .A2(new_n286), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n323), .A2(new_n211), .A3(G68), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT19), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n211), .B1(new_n269), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(G87), .B2(new_n207), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n211), .A2(G33), .A3(G97), .ZN(new_n548));
  AND3_X1   g0348(.A1(new_n548), .A2(KEYINPUT81), .A3(new_n545), .ZN(new_n549));
  AOI21_X1  g0349(.A(KEYINPUT81), .B1(new_n548), .B2(new_n545), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n544), .B(new_n547), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n543), .B1(new_n551), .B2(new_n297), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n483), .A2(new_n379), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT80), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(new_n274), .B2(G1), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n210), .A2(KEYINPUT80), .A3(G45), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n256), .A2(new_n556), .A3(G250), .A4(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n256), .A2(G274), .A3(new_n465), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n263), .A2(new_n265), .A3(G244), .A4(G1698), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n263), .A2(new_n265), .A3(G238), .A4(new_n267), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n561), .A2(new_n562), .A3(new_n514), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n560), .B1(new_n271), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n398), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n563), .A2(new_n271), .ZN(new_n566));
  INV_X1    g0366(.A(new_n560), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n396), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n554), .A2(new_n565), .A3(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(G87), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n482), .A2(new_n571), .ZN(new_n572));
  AOI211_X1 g0372(.A(new_n543), .B(new_n572), .C1(new_n551), .C2(new_n297), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n564), .A2(G190), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n568), .A2(new_n329), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  AND2_X1   g0376(.A1(new_n570), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n536), .A2(new_n398), .A3(new_n471), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n540), .A2(new_n396), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n331), .B1(new_n522), .B2(new_n524), .ZN(new_n580));
  INV_X1    g0380(.A(new_n530), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n578), .B(new_n579), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n507), .A2(new_n542), .A3(new_n577), .A4(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT79), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n263), .A2(new_n265), .A3(G244), .A4(new_n267), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT4), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n323), .A2(KEYINPUT4), .A3(G244), .A4(new_n267), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n323), .A2(G250), .A3(G1698), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n587), .A2(new_n588), .A3(new_n488), .A4(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n271), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n468), .A2(new_n256), .ZN(new_n592));
  INV_X1    g0392(.A(G257), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n471), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n396), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n594), .B1(new_n590), .B2(new_n271), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n398), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n386), .A2(new_n294), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT6), .ZN(new_n601));
  AND2_X1   g0401(.A1(G97), .A2(G107), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n601), .B1(new_n602), .B2(new_n206), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n369), .A2(KEYINPUT6), .A3(G97), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n600), .B1(new_n605), .B2(G20), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n438), .A2(new_n439), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n606), .A2(KEYINPUT78), .B1(new_n607), .B2(G107), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT78), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n211), .B1(new_n603), .B2(new_n604), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n609), .B1(new_n610), .B2(new_n600), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n331), .B1(new_n608), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n287), .A2(new_n489), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n482), .B2(new_n489), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n597), .B(new_n599), .C1(new_n612), .C2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n607), .A2(G107), .ZN(new_n616));
  INV_X1    g0416(.A(new_n600), .ZN(new_n617));
  NOR3_X1   g0417(.A1(new_n601), .A2(new_n489), .A3(G107), .ZN(new_n618));
  XNOR2_X1  g0418(.A(G97), .B(G107), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n618), .B1(new_n601), .B2(new_n619), .ZN(new_n620));
  OAI211_X1 g0420(.A(KEYINPUT78), .B(new_n617), .C1(new_n620), .C2(new_n211), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n616), .A2(new_n621), .A3(new_n611), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n614), .B1(new_n622), .B2(new_n297), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n598), .A2(G200), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n591), .A2(new_n416), .A3(new_n595), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n584), .B1(new_n615), .B2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n615), .A2(new_n626), .A3(new_n584), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n583), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n464), .A2(new_n630), .ZN(G372));
  NAND2_X1  g0431(.A1(new_n456), .A2(new_n462), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n310), .A2(new_n304), .A3(new_n285), .ZN(new_n634));
  INV_X1    g0434(.A(new_n400), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n365), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT85), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n446), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n637), .A2(new_n638), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n633), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n642), .A2(new_n354), .B1(new_n402), .B2(new_n404), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n498), .A2(new_n506), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n496), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n582), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n647), .A2(KEYINPUT84), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT84), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n582), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n646), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  AND4_X1   g0451(.A1(new_n615), .A2(new_n577), .A3(new_n626), .A4(new_n542), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n570), .ZN(new_n654));
  INV_X1    g0454(.A(new_n615), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n655), .A2(new_n577), .A3(KEYINPUT26), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT26), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n570), .A2(new_n576), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n657), .B1(new_n615), .B2(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n654), .B1(new_n656), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n653), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n464), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n643), .A2(new_n662), .ZN(G369));
  NAND4_X1  g0463(.A1(new_n496), .A2(new_n505), .A3(new_n498), .A4(new_n506), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n210), .A2(new_n211), .A3(G13), .ZN(new_n665));
  OAI21_X1  g0465(.A(G213), .B1(new_n665), .B2(KEYINPUT27), .ZN(new_n666));
  AOI21_X1  g0466(.A(KEYINPUT86), .B1(new_n665), .B2(KEYINPUT27), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n665), .A2(KEYINPUT86), .A3(KEYINPUT27), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n666), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(G343), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n502), .A2(new_n671), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n664), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n645), .A2(new_n672), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(G330), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n671), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(new_n580), .B2(new_n581), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n542), .A2(new_n582), .A3(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n680), .B1(new_n582), .B2(new_n671), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n645), .A2(new_n671), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(new_n680), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n648), .A2(new_n650), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n684), .B1(new_n685), .B2(new_n671), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n682), .A2(new_n686), .ZN(G399));
  INV_X1    g0487(.A(new_n214), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(G41), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR3_X1   g0490(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(G1), .A3(new_n691), .ZN(new_n692));
  OAI22_X1  g0492(.A1(new_n692), .A2(KEYINPUT87), .B1(new_n217), .B2(new_n690), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n693), .B1(KEYINPUT87), .B2(new_n692), .ZN(new_n694));
  XOR2_X1   g0494(.A(new_n694), .B(KEYINPUT28), .Z(new_n695));
  NAND4_X1  g0495(.A1(new_n497), .A2(new_n598), .A3(new_n536), .A4(new_n564), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT30), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n564), .A2(new_n536), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n699), .A2(KEYINPUT30), .A3(new_n497), .A4(new_n598), .ZN(new_n700));
  NOR3_X1   g0500(.A1(new_n504), .A2(G179), .A3(new_n564), .ZN(new_n701));
  AOI22_X1  g0501(.A1(new_n591), .A2(new_n595), .B1(new_n536), .B2(new_n471), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n698), .A2(new_n700), .A3(new_n703), .ZN(new_n704));
  XOR2_X1   g0504(.A(KEYINPUT88), .B(KEYINPUT31), .Z(new_n705));
  NAND3_X1  g0505(.A1(new_n704), .A2(new_n678), .A3(new_n705), .ZN(new_n706));
  AOI22_X1  g0506(.A1(new_n696), .A2(new_n697), .B1(new_n701), .B2(new_n702), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n671), .B1(new_n707), .B2(new_n700), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n706), .B1(KEYINPUT31), .B2(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n709), .B1(new_n630), .B2(new_n671), .ZN(new_n710));
  INV_X1    g0510(.A(G330), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT89), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n644), .A2(new_n713), .A3(new_n582), .A4(new_n496), .ZN(new_n714));
  OAI21_X1  g0514(.A(KEYINPUT89), .B1(new_n645), .B2(new_n647), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n652), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n678), .B1(new_n716), .B2(new_n660), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT29), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI211_X1 g0519(.A(KEYINPUT29), .B(new_n678), .C1(new_n653), .C2(new_n660), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n712), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n695), .B1(new_n721), .B2(G1), .ZN(G364));
  INV_X1    g0522(.A(G13), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G20), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n210), .B1(new_n724), .B2(G45), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n689), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n219), .B1(G20), .B2(new_n396), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n211), .A2(new_n398), .ZN(new_n731));
  NOR2_X1   g0531(.A1(G190), .A2(G200), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(G311), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n428), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n211), .A2(G179), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(new_n732), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  AND2_X1   g0538(.A1(new_n738), .A2(G329), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n731), .A2(G190), .A3(new_n306), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  AOI211_X1 g0541(.A(new_n735), .B(new_n739), .C1(G322), .C2(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n329), .A2(G190), .A3(new_n736), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G303), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n329), .A2(new_n416), .A3(new_n736), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n746), .B1(G283), .B2(new_n748), .ZN(new_n749));
  NOR3_X1   g0549(.A1(new_n416), .A2(G179), .A3(G200), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n211), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n731), .A2(G200), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n416), .ZN(new_n754));
  AOI22_X1  g0554(.A1(G294), .A2(new_n752), .B1(new_n754), .B2(G326), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n753), .A2(G190), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  XOR2_X1   g0557(.A(KEYINPUT33), .B(G317), .Z(new_n758));
  OAI211_X1 g0558(.A(new_n749), .B(new_n755), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n323), .B1(new_n733), .B2(new_n294), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n760), .B1(G58), .B2(new_n741), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n751), .A2(new_n489), .ZN(new_n762));
  INV_X1    g0562(.A(G159), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n737), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n762), .B1(KEYINPUT32), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n744), .A2(G87), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n748), .A2(G107), .ZN(new_n768));
  AND4_X1   g0568(.A1(new_n761), .A2(new_n766), .A3(new_n767), .A4(new_n768), .ZN(new_n769));
  AOI22_X1  g0569(.A1(G50), .A2(new_n754), .B1(new_n756), .B2(G68), .ZN(new_n770));
  OAI211_X1 g0570(.A(new_n769), .B(new_n770), .C1(KEYINPUT32), .C2(new_n765), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n730), .B1(new_n759), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G13), .A2(G33), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(G20), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n729), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n688), .A2(new_n428), .ZN(new_n777));
  AOI22_X1  g0577(.A1(G355), .A2(new_n777), .B1(new_n485), .B2(new_n688), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n688), .A2(new_n323), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n779), .B1(G45), .B2(new_n217), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n252), .A2(new_n274), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n778), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n728), .B(new_n772), .C1(new_n776), .C2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n775), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n783), .B1(new_n675), .B2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(KEYINPUT90), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n676), .B(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n728), .B1(new_n675), .B2(G330), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n785), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT91), .ZN(G396));
  NAND2_X1  g0590(.A1(new_n661), .A2(new_n671), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n400), .A2(new_n678), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n394), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n794), .B1(new_n395), .B2(new_n678), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n793), .B1(new_n795), .B2(new_n635), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n791), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n796), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n661), .A2(new_n671), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(new_n711), .B2(new_n710), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n797), .A2(new_n712), .A3(new_n799), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n801), .A2(new_n728), .A3(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n733), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n741), .A2(G143), .B1(new_n804), .B2(G159), .ZN(new_n805));
  INV_X1    g0605(.A(G150), .ZN(new_n806));
  INV_X1    g0606(.A(G137), .ZN(new_n807));
  INV_X1    g0607(.A(new_n754), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n805), .B1(new_n757), .B2(new_n806), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n809), .B(KEYINPUT93), .Z(new_n810));
  OR2_X1    g0610(.A1(new_n810), .A2(KEYINPUT34), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(KEYINPUT34), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n747), .A2(new_n248), .ZN(new_n813));
  INV_X1    g0613(.A(G132), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n323), .B1(new_n737), .B2(new_n814), .C1(new_n751), .C2(new_n332), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n813), .B(new_n815), .C1(G50), .C2(new_n744), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n811), .A2(new_n812), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n748), .A2(G87), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(new_n734), .B2(new_n737), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT92), .ZN(new_n820));
  INV_X1    g0620(.A(G303), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n808), .A2(new_n821), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n762), .B(new_n822), .C1(G283), .C2(new_n756), .ZN(new_n823));
  INV_X1    g0623(.A(G294), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n428), .B1(new_n733), .B2(new_n485), .C1(new_n824), .C2(new_n740), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(G107), .B2(new_n744), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n820), .A2(new_n823), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n730), .B1(new_n817), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n729), .A2(new_n773), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n728), .B(new_n828), .C1(new_n294), .C2(new_n829), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(new_n774), .B2(new_n798), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n803), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT94), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n803), .A2(KEYINPUT94), .A3(new_n831), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(G384));
  NOR2_X1   g0636(.A1(new_n724), .A2(new_n210), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT40), .ZN(new_n838));
  INV_X1    g0638(.A(new_n455), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n422), .A2(new_n443), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n450), .A2(new_n670), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(KEYINPUT37), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT37), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n455), .A2(new_n844), .A3(new_n840), .A4(new_n841), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n843), .A2(KEYINPUT96), .A3(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT96), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n847), .B(KEYINPUT37), .C1(new_n839), .C2(new_n842), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT38), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT17), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n840), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n422), .A2(KEYINPUT17), .A3(new_n443), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n456), .A2(new_n462), .A3(new_n852), .A4(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n841), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n850), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n854), .A2(new_n855), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n846), .A2(new_n857), .A3(new_n848), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n849), .A2(new_n856), .B1(new_n858), .B2(new_n850), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT31), .ZN(new_n860));
  AOI211_X1 g0660(.A(new_n860), .B(new_n671), .C1(new_n707), .C2(new_n700), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n705), .B1(new_n704), .B2(new_n678), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n542), .A2(new_n582), .A3(new_n570), .A4(new_n576), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n864), .A2(new_n664), .ZN(new_n865));
  AND3_X1   g0665(.A1(new_n615), .A2(new_n626), .A3(new_n584), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n865), .B(new_n671), .C1(new_n627), .C2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n355), .A2(new_n678), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n634), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n365), .ZN(new_n871));
  OAI21_X1  g0671(.A(G169), .B1(new_n359), .B2(new_n360), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(KEYINPUT14), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n873), .A2(new_n362), .A3(new_n361), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n874), .B1(new_n308), .B2(new_n311), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n871), .B1(new_n875), .B2(new_n869), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n868), .A2(new_n876), .A3(new_n798), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n838), .B1(new_n859), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(KEYINPUT98), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT98), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n880), .B(new_n838), .C1(new_n859), .C2(new_n877), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT99), .ZN(new_n883));
  AND3_X1   g0683(.A1(new_n856), .A2(new_n848), .A3(new_n846), .ZN(new_n884));
  XNOR2_X1  g0684(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n843), .A2(new_n845), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n886), .B1(new_n857), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(KEYINPUT40), .B1(new_n884), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n883), .B1(new_n889), .B2(new_n877), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n857), .A2(new_n887), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n885), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n856), .A2(new_n848), .A3(new_n846), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n838), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n877), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n894), .A2(new_n895), .A3(KEYINPUT99), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n890), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n882), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n868), .A2(new_n464), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n898), .A2(new_n899), .ZN(new_n901));
  NOR3_X1   g0701(.A1(new_n900), .A2(new_n901), .A3(new_n711), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n892), .A2(new_n893), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT39), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n858), .A2(new_n850), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n893), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n906), .B1(new_n905), .B2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n365), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n671), .ZN(new_n911));
  OR2_X1    g0711(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n876), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n792), .B(KEYINPUT95), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n913), .B1(new_n799), .B2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n670), .ZN(new_n917));
  AOI22_X1  g0717(.A1(new_n916), .A2(new_n908), .B1(new_n632), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n912), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n464), .B1(new_n719), .B2(new_n720), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n643), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n919), .B(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n837), .B1(new_n903), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n922), .B2(new_n903), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n605), .A2(KEYINPUT35), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n605), .A2(KEYINPUT35), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n925), .A2(new_n926), .A3(G116), .A4(new_n220), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT36), .ZN(new_n928));
  OAI21_X1  g0728(.A(G77), .B1(new_n332), .B2(new_n248), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n247), .B1(new_n929), .B2(new_n217), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n930), .A2(G1), .A3(new_n723), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n924), .A2(new_n928), .A3(new_n931), .ZN(G367));
  OAI21_X1  g0732(.A(new_n776), .B1(new_n214), .B2(new_n388), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n933), .B1(new_n779), .B2(new_n242), .ZN(new_n934));
  AOI21_X1  g0734(.A(KEYINPUT46), .B1(new_n744), .B2(G116), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT105), .ZN(new_n936));
  OAI22_X1  g0736(.A1(new_n757), .A2(new_n824), .B1(new_n808), .B2(new_n734), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n747), .A2(new_n489), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n323), .B1(new_n738), .B2(G317), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n821), .B2(new_n740), .ZN(new_n940));
  NOR3_X1   g0740(.A1(new_n937), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(G283), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n751), .A2(new_n369), .B1(new_n733), .B2(new_n942), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n943), .B(KEYINPUT103), .Z(new_n944));
  NAND3_X1  g0744(.A1(new_n936), .A2(new_n941), .A3(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n744), .A2(KEYINPUT46), .A3(G116), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n946), .B(KEYINPUT104), .Z(new_n947));
  NOR2_X1   g0747(.A1(new_n751), .A2(new_n248), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n948), .B1(G143), .B2(new_n754), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n763), .B2(new_n757), .ZN(new_n950));
  OAI22_X1  g0750(.A1(new_n740), .A2(new_n806), .B1(new_n733), .B2(new_n202), .ZN(new_n951));
  AOI211_X1 g0751(.A(new_n428), .B(new_n951), .C1(G137), .C2(new_n738), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n748), .A2(G77), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n744), .A2(G58), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n945), .A2(new_n947), .B1(new_n950), .B2(new_n955), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT47), .ZN(new_n957));
  AOI211_X1 g0757(.A(new_n728), .B(new_n934), .C1(new_n957), .C2(new_n729), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n573), .A2(new_n671), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n570), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n577), .B2(new_n959), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT100), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n958), .B1(new_n963), .B2(new_n784), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n615), .A2(new_n626), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n678), .B1(new_n612), .B2(new_n614), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n655), .A2(new_n678), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n686), .A2(new_n970), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n971), .A2(KEYINPUT102), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(KEYINPUT102), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT45), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n972), .A2(KEYINPUT45), .A3(new_n973), .ZN(new_n977));
  INV_X1    g0777(.A(new_n970), .ZN(new_n978));
  NOR3_X1   g0778(.A1(new_n648), .A2(new_n650), .A3(new_n678), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n978), .B1(new_n979), .B2(new_n684), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT44), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n976), .A2(new_n977), .A3(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n682), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n684), .ZN(new_n986));
  INV_X1    g0786(.A(new_n683), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n986), .B1(new_n681), .B2(new_n987), .ZN(new_n988));
  MUX2_X1   g0788(.A(new_n676), .B(new_n787), .S(new_n988), .Z(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n721), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n981), .B1(new_n974), .B2(new_n975), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n992), .A2(new_n682), .A3(new_n977), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n985), .A2(new_n991), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n721), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n689), .B(KEYINPUT41), .Z(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n726), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n966), .A2(new_n647), .A3(new_n967), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n678), .B1(new_n999), .B2(new_n615), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n970), .A2(new_n684), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1000), .B1(new_n1001), .B2(KEYINPUT42), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(KEYINPUT42), .B2(new_n1001), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT43), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1003), .B1(new_n1004), .B2(new_n962), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n962), .A2(new_n1004), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT101), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1005), .B(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n682), .A2(new_n978), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n964), .B1(new_n998), .B2(new_n1012), .ZN(G387));
  NOR2_X1   g0813(.A1(new_n991), .A2(new_n690), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n721), .B2(new_n989), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n989), .A2(new_n726), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n323), .B1(new_n738), .B2(G326), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(G311), .A2(new_n756), .B1(new_n754), .B2(G322), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n1018), .A2(KEYINPUT107), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(KEYINPUT107), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n741), .A2(G317), .B1(new_n804), .B2(G303), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT48), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n744), .A2(G294), .B1(new_n752), .B2(G283), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT49), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1017), .B1(new_n485), .B2(new_n747), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(new_n1028), .B2(new_n1027), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n752), .A2(new_n379), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n1031), .B1(new_n757), .B2(new_n385), .C1(new_n763), .C2(new_n808), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n428), .B1(new_n738), .B2(G150), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1033), .B1(new_n202), .B2(new_n740), .C1(new_n248), .C2(new_n733), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n743), .A2(new_n294), .ZN(new_n1035));
  NOR4_X1   g0835(.A1(new_n1032), .A2(new_n1034), .A3(new_n938), .A4(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n729), .B1(new_n1030), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n691), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n777), .A2(new_n1038), .B1(new_n369), .B2(new_n688), .ZN(new_n1039));
  AND2_X1   g0839(.A1(new_n239), .A2(G45), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n336), .A2(new_n202), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT50), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n691), .B(new_n274), .C1(new_n248), .C2(new_n294), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n779), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT106), .Z(new_n1045));
  OAI21_X1  g0845(.A(new_n1039), .B1(new_n1040), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n728), .B1(new_n1046), .B2(new_n776), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1037), .B(new_n1047), .C1(new_n681), .C2(new_n784), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1015), .A2(new_n1016), .A3(new_n1048), .ZN(G393));
  NOR2_X1   g0849(.A1(new_n983), .A2(new_n984), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n682), .B1(new_n992), .B2(new_n977), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n990), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1052), .A2(new_n689), .A3(new_n994), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n985), .A2(new_n726), .A3(new_n993), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n779), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n776), .B1(new_n489), .B2(new_n214), .C1(new_n1055), .C2(new_n246), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(new_n727), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G116), .A2(new_n752), .B1(new_n756), .B2(G303), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n428), .B1(new_n733), .B2(new_n824), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(G322), .B2(new_n738), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n744), .A2(G283), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1058), .A2(new_n1060), .A3(new_n768), .A4(new_n1061), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(G317), .A2(new_n754), .B1(new_n741), .B2(G311), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT52), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(G150), .A2(new_n754), .B1(new_n741), .B2(G159), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT51), .ZN(new_n1066));
  INV_X1    g0866(.A(G143), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n323), .B1(new_n737), .B2(new_n1067), .C1(new_n385), .C2(new_n733), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G77), .A2(new_n752), .B1(new_n756), .B2(G50), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n744), .A2(G68), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1069), .A2(new_n1070), .A3(new_n818), .A4(new_n1071), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n1062), .A2(new_n1064), .B1(new_n1066), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1057), .B1(new_n1073), .B2(new_n729), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n970), .B2(new_n784), .ZN(new_n1075));
  AND2_X1   g0875(.A1(new_n1054), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1053), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT108), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1053), .A2(new_n1076), .A3(KEYINPUT108), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(new_n1080), .ZN(G390));
  NAND2_X1  g0881(.A1(new_n909), .A2(new_n773), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n738), .A2(G125), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n323), .B1(new_n747), .B2(new_n202), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT114), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1083), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(new_n1085), .B2(new_n1084), .ZN(new_n1087));
  XOR2_X1   g0887(.A(new_n1087), .B(KEYINPUT115), .Z(new_n1088));
  OAI22_X1  g0888(.A1(new_n757), .A2(new_n807), .B1(new_n814), .B2(new_n740), .ZN(new_n1089));
  INV_X1    g0889(.A(G128), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n808), .A2(new_n1090), .B1(new_n763), .B2(new_n751), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n743), .A2(new_n806), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT53), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(KEYINPUT54), .B(G143), .ZN(new_n1095));
  XOR2_X1   g0895(.A(new_n1095), .B(KEYINPUT113), .Z(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1092), .B(new_n1094), .C1(new_n733), .C2(new_n1097), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(G77), .A2(new_n752), .B1(new_n754), .B2(G283), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n369), .B2(new_n757), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n813), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(G97), .A2(new_n804), .B1(new_n738), .B2(G294), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n323), .B1(new_n741), .B2(G116), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1101), .A2(new_n767), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n1088), .A2(new_n1098), .B1(new_n1100), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n729), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n728), .B1(new_n385), .B2(new_n829), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1082), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n911), .ZN(new_n1109));
  OAI21_X1  g0909(.A(KEYINPUT110), .B1(new_n916), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n678), .B1(new_n653), .B2(new_n660), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n914), .B1(new_n1112), .B2(new_n798), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1111), .B(new_n911), .C1(new_n1113), .C2(new_n913), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1110), .A2(new_n909), .A3(new_n1114), .ZN(new_n1115));
  XOR2_X1   g0915(.A(new_n911), .B(KEYINPUT109), .Z(new_n1116));
  AOI21_X1  g0916(.A(new_n914), .B1(new_n717), .B2(new_n798), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1116), .B(new_n904), .C1(new_n1117), .C2(new_n913), .ZN(new_n1118));
  OR2_X1    g0918(.A1(new_n708), .A2(KEYINPUT31), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n867), .A2(new_n1119), .A3(new_n706), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n796), .A2(new_n711), .ZN(new_n1121));
  AND3_X1   g0921(.A1(new_n1120), .A2(new_n876), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  AND3_X1   g0923(.A1(new_n1115), .A2(new_n1118), .A3(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n868), .A2(new_n876), .A3(new_n1121), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(KEYINPUT111), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT111), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n868), .A2(new_n876), .A3(new_n1127), .A4(new_n1121), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(new_n1115), .B2(new_n1118), .ZN(new_n1130));
  OR2_X1    g0930(.A1(new_n1124), .A2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1108), .B1(new_n1131), .B2(new_n725), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1121), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n913), .B1(new_n710), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1126), .A2(new_n1128), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1113), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n876), .B1(new_n868), .B2(new_n1121), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1122), .A2(new_n1137), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n1135), .A2(new_n1136), .B1(new_n1138), .B2(new_n1117), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n868), .A2(new_n464), .A3(G330), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(KEYINPUT112), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT112), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n868), .A2(new_n464), .A3(new_n1142), .A4(G330), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1144), .A2(new_n643), .A3(new_n920), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1139), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n690), .B1(new_n1131), .B2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1124), .A2(new_n1130), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n1146), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1132), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(G378));
  AOI21_X1  g0952(.A(new_n711), .B1(new_n890), .B2(new_n896), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n882), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n402), .A2(new_n404), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n354), .A2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n403), .A2(new_n917), .ZN(new_n1157));
  OR2_X1    g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1160));
  AND3_X1   g0960(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1160), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1154), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT117), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1163), .A2(KEYINPUT116), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT116), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n882), .A2(new_n1153), .A3(new_n1165), .A4(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1164), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n882), .A2(new_n1153), .A3(new_n1169), .ZN(new_n1172));
  AND2_X1   g0972(.A1(new_n1172), .A2(KEYINPUT117), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n919), .B1(new_n1171), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1172), .A2(KEYINPUT117), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n919), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1175), .A2(new_n1164), .A3(new_n1176), .A4(new_n1170), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1174), .A2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1166), .A2(new_n773), .A3(new_n1168), .ZN(new_n1179));
  NOR3_X1   g0979(.A1(new_n729), .A2(G50), .A3(new_n773), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(new_n428), .B2(new_n273), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n740), .A2(new_n369), .B1(new_n733), .B2(new_n388), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n273), .B(new_n428), .C1(new_n737), .C2(new_n942), .ZN(new_n1184));
  NOR3_X1   g0984(.A1(new_n1035), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n754), .A2(G116), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n948), .B1(G97), .B2(new_n756), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n748), .A2(G58), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT58), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1182), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n740), .A2(new_n1090), .B1(new_n733), .B2(new_n807), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(G132), .B2(new_n756), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(G150), .A2(new_n752), .B1(new_n754), .B2(G125), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1193), .B(new_n1194), .C1(new_n1097), .C2(new_n743), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(KEYINPUT59), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n748), .A2(G159), .ZN(new_n1197));
  AOI211_X1 g0997(.A(G33), .B(G41), .C1(new_n738), .C2(G124), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1195), .A2(KEYINPUT59), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1191), .B1(new_n1190), .B2(new_n1189), .C1(new_n1199), .C2(new_n1200), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n728), .B(new_n1180), .C1(new_n1201), .C2(new_n729), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n1178), .A2(new_n726), .B1(new_n1179), .B2(new_n1202), .ZN(new_n1203));
  AND3_X1   g1003(.A1(new_n1144), .A2(new_n643), .A3(new_n920), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1150), .A2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1163), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(new_n882), .B2(new_n1153), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n882), .A2(new_n1153), .A3(new_n1169), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1207), .B1(new_n1208), .B2(new_n1165), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1176), .B1(new_n1209), .B2(new_n1175), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1177), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1205), .B(KEYINPUT57), .C1(new_n1210), .C2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(new_n689), .ZN(new_n1213));
  AOI21_X1  g1013(.A(KEYINPUT57), .B1(new_n1178), .B2(new_n1205), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1203), .B1(new_n1213), .B2(new_n1214), .ZN(G375));
  NAND2_X1  g1015(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1138), .A2(new_n1117), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1145), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1147), .A2(new_n997), .A3(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n913), .A2(new_n773), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n728), .B1(new_n248), .B2(new_n829), .ZN(new_n1222));
  XOR2_X1   g1022(.A(new_n1222), .B(KEYINPUT118), .Z(new_n1223));
  OAI221_X1 g1023(.A(new_n1188), .B1(new_n763), .B2(new_n743), .C1(new_n1097), .C2(new_n757), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(G50), .A2(new_n752), .B1(new_n754), .B2(G132), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n428), .B1(new_n738), .B2(G128), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n741), .A2(G137), .B1(new_n804), .B2(G150), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n741), .A2(G283), .B1(new_n804), .B2(G107), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n744), .A2(G97), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n323), .B1(new_n738), .B2(G303), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1229), .A2(new_n953), .A3(new_n1230), .A4(new_n1231), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n1031), .B1(new_n757), .B2(new_n485), .C1(new_n824), .C2(new_n808), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n1224), .A2(new_n1228), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1223), .B1(new_n1234), .B2(new_n729), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n1220), .A2(new_n726), .B1(new_n1221), .B2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1219), .A2(new_n1236), .ZN(G381));
  INV_X1    g1037(.A(KEYINPUT119), .ZN(new_n1238));
  OR2_X1    g1038(.A1(G375), .A2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(G375), .A2(new_n1238), .ZN(new_n1240));
  OR4_X1    g1040(.A1(G396), .A2(G393), .A3(G381), .A4(G384), .ZN(new_n1241));
  NOR3_X1   g1041(.A1(new_n1241), .A2(G390), .A3(G387), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1239), .A2(new_n1151), .A3(new_n1240), .A4(new_n1242), .ZN(G407));
  NAND3_X1  g1043(.A1(new_n1239), .A2(new_n1151), .A3(new_n1240), .ZN(new_n1244));
  INV_X1    g1044(.A(G343), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(G213), .ZN(new_n1246));
  XOR2_X1   g1046(.A(new_n1246), .B(KEYINPUT120), .Z(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  OAI211_X1 g1048(.A(G407), .B(G213), .C1(new_n1244), .C2(new_n1248), .ZN(G409));
  INV_X1    g1049(.A(KEYINPUT126), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n996), .B1(new_n994), .B2(new_n721), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1011), .B(new_n1010), .C1(new_n1251), .C2(new_n726), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n1053), .A2(new_n1076), .A3(KEYINPUT108), .ZN(new_n1253));
  AOI21_X1  g1053(.A(KEYINPUT108), .B1(new_n1053), .B2(new_n1076), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1252), .B(new_n964), .C1(new_n1253), .C2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(G387), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1256));
  XOR2_X1   g1056(.A(G393), .B(G396), .Z(new_n1257));
  NAND3_X1  g1057(.A1(new_n1255), .A2(new_n1256), .A3(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1257), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1250), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1257), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1264), .A2(KEYINPUT126), .A3(new_n1258), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1261), .A2(new_n1265), .ZN(new_n1266));
  OAI211_X1 g1066(.A(G378), .B(new_n1203), .C1(new_n1213), .C2(new_n1214), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1178), .A2(new_n726), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1179), .A2(new_n1202), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  AND3_X1   g1070(.A1(new_n1178), .A2(new_n997), .A3(new_n1205), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1151), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1267), .A2(new_n1272), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1145), .A2(new_n1216), .A3(KEYINPUT60), .A4(new_n1217), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(KEYINPUT121), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n690), .B1(new_n1220), .B2(new_n1204), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT60), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1218), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT121), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1139), .A2(new_n1279), .A3(KEYINPUT60), .A4(new_n1145), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1275), .A2(new_n1276), .A3(new_n1278), .A4(new_n1280), .ZN(new_n1281));
  AND3_X1   g1081(.A1(new_n1281), .A2(G384), .A3(new_n1236), .ZN(new_n1282));
  AOI21_X1  g1082(.A(G384), .B1(new_n1281), .B2(new_n1236), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1273), .A2(new_n1246), .A3(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT62), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1247), .B1(new_n1267), .B2(new_n1272), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1284), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1288), .A2(new_n1286), .ZN(new_n1289));
  AOI22_X1  g1089(.A1(new_n1285), .A2(new_n1286), .B1(new_n1287), .B2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT61), .ZN(new_n1291));
  AND2_X1   g1091(.A1(new_n1247), .A2(G2897), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1292), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT123), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  OAI211_X1 g1095(.A(KEYINPUT123), .B(new_n1292), .C1(new_n1282), .C2(new_n1283), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1281), .A2(new_n1236), .ZN(new_n1298));
  INV_X1    g1098(.A(G384), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1281), .A2(G384), .A3(new_n1236), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1245), .A2(G213), .A3(G2897), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1300), .A2(new_n1301), .A3(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT122), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1300), .A2(KEYINPUT122), .A3(new_n1301), .A4(new_n1302), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1297), .A2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT124), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1297), .A2(new_n1307), .A3(KEYINPUT124), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1291), .B1(new_n1312), .B2(new_n1287), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1266), .B1(new_n1290), .B2(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1264), .A2(new_n1291), .A3(new_n1258), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT63), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1288), .A2(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1315), .B1(new_n1287), .B2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1285), .A2(new_n1316), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1310), .A2(KEYINPUT125), .A3(new_n1311), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1273), .A2(new_n1246), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(KEYINPUT125), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1323));
  OAI211_X1 g1123(.A(new_n1318), .B(new_n1319), .C1(new_n1322), .C2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1314), .A2(new_n1324), .ZN(G405));
  NOR3_X1   g1125(.A1(new_n1259), .A2(new_n1260), .A3(new_n1250), .ZN(new_n1326));
  AOI21_X1  g1126(.A(KEYINPUT126), .B1(new_n1264), .B2(new_n1258), .ZN(new_n1327));
  OAI21_X1  g1127(.A(KEYINPUT127), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(G375), .A2(new_n1151), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1329), .A2(new_n1288), .A3(new_n1267), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1288), .B1(new_n1329), .B2(new_n1267), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT127), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1261), .A2(new_n1265), .A3(new_n1333), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1328), .A2(new_n1330), .A3(new_n1332), .A4(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1330), .ZN(new_n1336));
  OAI211_X1 g1136(.A(new_n1266), .B(KEYINPUT127), .C1(new_n1336), .C2(new_n1331), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1335), .A2(new_n1337), .ZN(G402));
endmodule


