

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U554 ( .A(KEYINPUT66), .B(n536), .Z(n643) );
  XOR2_X2 U555 ( .A(KEYINPUT93), .B(n751), .Z(n788) );
  OR2_X1 U556 ( .A1(n518), .A2(n803), .ZN(n804) );
  NOR2_X1 U557 ( .A1(n780), .A2(n779), .ZN(n800) );
  XNOR2_X1 U558 ( .A(n773), .B(n772), .ZN(n780) );
  NOR2_X1 U559 ( .A1(n788), .A2(n787), .ZN(n789) );
  NOR2_X1 U560 ( .A1(n800), .A2(n799), .ZN(n802) );
  XOR2_X1 U561 ( .A(n731), .B(KEYINPUT96), .Z(n517) );
  AND2_X1 U562 ( .A1(n796), .A2(n801), .ZN(n518) );
  XNOR2_X1 U563 ( .A(n743), .B(KEYINPUT29), .ZN(n744) );
  XNOR2_X1 U564 ( .A(n745), .B(n744), .ZN(n750) );
  NOR2_X1 U565 ( .A1(n750), .A2(n749), .ZN(n761) );
  INV_X1 U566 ( .A(KEYINPUT100), .ZN(n762) );
  INV_X1 U567 ( .A(KEYINPUT32), .ZN(n772) );
  NOR2_X1 U568 ( .A1(G164), .A2(G1384), .ZN(n716) );
  NAND2_X1 U569 ( .A1(n587), .A2(n586), .ZN(n923) );
  INV_X1 U570 ( .A(G2105), .ZN(n522) );
  AND2_X1 U571 ( .A1(n522), .A2(G2104), .ZN(n881) );
  NAND2_X1 U572 ( .A1(G102), .A2(n881), .ZN(n521) );
  NOR2_X1 U573 ( .A1(G2104), .A2(G2105), .ZN(n519) );
  XOR2_X2 U574 ( .A(KEYINPUT17), .B(n519), .Z(n882) );
  NAND2_X1 U575 ( .A1(G138), .A2(n882), .ZN(n520) );
  NAND2_X1 U576 ( .A1(n521), .A2(n520), .ZN(n526) );
  AND2_X1 U577 ( .A1(G2104), .A2(G2105), .ZN(n877) );
  NAND2_X1 U578 ( .A1(G114), .A2(n877), .ZN(n524) );
  NOR2_X1 U579 ( .A1(G2104), .A2(n522), .ZN(n878) );
  NAND2_X1 U580 ( .A1(G126), .A2(n878), .ZN(n523) );
  NAND2_X1 U581 ( .A1(n524), .A2(n523), .ZN(n525) );
  NOR2_X1 U582 ( .A1(n526), .A2(n525), .ZN(G164) );
  XNOR2_X1 U583 ( .A(KEYINPUT70), .B(KEYINPUT6), .ZN(n532) );
  INV_X1 U584 ( .A(G651), .ZN(n535) );
  NOR2_X1 U585 ( .A1(G543), .A2(n535), .ZN(n527) );
  XOR2_X1 U586 ( .A(KEYINPUT1), .B(n527), .Z(n639) );
  NAND2_X1 U587 ( .A1(G63), .A2(n639), .ZN(n530) );
  XOR2_X1 U588 ( .A(KEYINPUT0), .B(G543), .Z(n534) );
  NOR2_X1 U589 ( .A1(n534), .A2(G651), .ZN(n528) );
  XNOR2_X1 U590 ( .A(KEYINPUT64), .B(n528), .ZN(n637) );
  NAND2_X1 U591 ( .A1(G51), .A2(n637), .ZN(n529) );
  NAND2_X1 U592 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U593 ( .A(n532), .B(n531), .ZN(n541) );
  NOR2_X1 U594 ( .A1(G543), .A2(G651), .ZN(n640) );
  NAND2_X1 U595 ( .A1(n640), .A2(G89), .ZN(n533) );
  XNOR2_X1 U596 ( .A(n533), .B(KEYINPUT4), .ZN(n538) );
  OR2_X1 U597 ( .A1(n535), .A2(n534), .ZN(n536) );
  NAND2_X1 U598 ( .A1(G76), .A2(n643), .ZN(n537) );
  NAND2_X1 U599 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U600 ( .A(KEYINPUT5), .B(n539), .Z(n540) );
  NOR2_X1 U601 ( .A1(n541), .A2(n540), .ZN(n543) );
  XNOR2_X1 U602 ( .A(KEYINPUT7), .B(KEYINPUT71), .ZN(n542) );
  XNOR2_X1 U603 ( .A(n543), .B(n542), .ZN(G168) );
  XOR2_X1 U604 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U605 ( .A1(G65), .A2(n639), .ZN(n545) );
  NAND2_X1 U606 ( .A1(G91), .A2(n640), .ZN(n544) );
  NAND2_X1 U607 ( .A1(n545), .A2(n544), .ZN(n548) );
  NAND2_X1 U608 ( .A1(G78), .A2(n643), .ZN(n546) );
  XNOR2_X1 U609 ( .A(KEYINPUT67), .B(n546), .ZN(n547) );
  NOR2_X1 U610 ( .A1(n548), .A2(n547), .ZN(n550) );
  NAND2_X1 U611 ( .A1(G53), .A2(n637), .ZN(n549) );
  NAND2_X1 U612 ( .A1(n550), .A2(n549), .ZN(G299) );
  NAND2_X1 U613 ( .A1(G101), .A2(n881), .ZN(n551) );
  XOR2_X1 U614 ( .A(KEYINPUT23), .B(n551), .Z(n680) );
  NAND2_X1 U615 ( .A1(G137), .A2(n882), .ZN(n552) );
  XOR2_X1 U616 ( .A(KEYINPUT65), .B(n552), .Z(n684) );
  NAND2_X1 U617 ( .A1(G113), .A2(n877), .ZN(n554) );
  NAND2_X1 U618 ( .A1(G125), .A2(n878), .ZN(n553) );
  AND2_X1 U619 ( .A1(n554), .A2(n553), .ZN(n682) );
  AND2_X1 U620 ( .A1(n684), .A2(n682), .ZN(n555) );
  AND2_X1 U621 ( .A1(n680), .A2(n555), .ZN(G160) );
  AND2_X1 U622 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U623 ( .A1(G111), .A2(n877), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n556), .B(KEYINPUT74), .ZN(n560) );
  XOR2_X1 U625 ( .A(KEYINPUT18), .B(KEYINPUT73), .Z(n558) );
  NAND2_X1 U626 ( .A1(G123), .A2(n878), .ZN(n557) );
  XNOR2_X1 U627 ( .A(n558), .B(n557), .ZN(n559) );
  NAND2_X1 U628 ( .A1(n560), .A2(n559), .ZN(n564) );
  NAND2_X1 U629 ( .A1(G99), .A2(n881), .ZN(n562) );
  NAND2_X1 U630 ( .A1(G135), .A2(n882), .ZN(n561) );
  NAND2_X1 U631 ( .A1(n562), .A2(n561), .ZN(n563) );
  NOR2_X1 U632 ( .A1(n564), .A2(n563), .ZN(n1009) );
  XNOR2_X1 U633 ( .A(n1009), .B(G2096), .ZN(n565) );
  XNOR2_X1 U634 ( .A(n565), .B(KEYINPUT75), .ZN(n566) );
  OR2_X1 U635 ( .A1(G2100), .A2(n566), .ZN(G156) );
  INV_X1 U636 ( .A(G57), .ZN(G237) );
  INV_X1 U637 ( .A(G108), .ZN(G238) );
  INV_X1 U638 ( .A(G132), .ZN(G219) );
  INV_X1 U639 ( .A(G82), .ZN(G220) );
  NAND2_X1 U640 ( .A1(G64), .A2(n639), .ZN(n568) );
  NAND2_X1 U641 ( .A1(G52), .A2(n637), .ZN(n567) );
  NAND2_X1 U642 ( .A1(n568), .A2(n567), .ZN(n573) );
  NAND2_X1 U643 ( .A1(G90), .A2(n640), .ZN(n570) );
  NAND2_X1 U644 ( .A1(G77), .A2(n643), .ZN(n569) );
  NAND2_X1 U645 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U646 ( .A(KEYINPUT9), .B(n571), .Z(n572) );
  NOR2_X1 U647 ( .A1(n573), .A2(n572), .ZN(G171) );
  NAND2_X1 U648 ( .A1(G7), .A2(G661), .ZN(n574) );
  XNOR2_X1 U649 ( .A(n574), .B(KEYINPUT10), .ZN(n575) );
  XNOR2_X1 U650 ( .A(KEYINPUT68), .B(n575), .ZN(G223) );
  INV_X1 U651 ( .A(G567), .ZN(n675) );
  NOR2_X1 U652 ( .A1(n675), .A2(G223), .ZN(n576) );
  XOR2_X1 U653 ( .A(KEYINPUT11), .B(n576), .Z(n577) );
  XNOR2_X1 U654 ( .A(KEYINPUT69), .B(n577), .ZN(G234) );
  NAND2_X1 U655 ( .A1(G68), .A2(n643), .ZN(n580) );
  NAND2_X1 U656 ( .A1(n640), .A2(G81), .ZN(n578) );
  XNOR2_X1 U657 ( .A(n578), .B(KEYINPUT12), .ZN(n579) );
  NAND2_X1 U658 ( .A1(n580), .A2(n579), .ZN(n582) );
  INV_X1 U659 ( .A(KEYINPUT13), .ZN(n581) );
  XNOR2_X1 U660 ( .A(n582), .B(n581), .ZN(n585) );
  NAND2_X1 U661 ( .A1(G56), .A2(n639), .ZN(n583) );
  XOR2_X1 U662 ( .A(KEYINPUT14), .B(n583), .Z(n584) );
  NOR2_X1 U663 ( .A1(n585), .A2(n584), .ZN(n587) );
  NAND2_X1 U664 ( .A1(G43), .A2(n637), .ZN(n586) );
  INV_X1 U665 ( .A(G860), .ZN(n600) );
  OR2_X1 U666 ( .A1(n923), .A2(n600), .ZN(G153) );
  INV_X1 U667 ( .A(G171), .ZN(G301) );
  NAND2_X1 U668 ( .A1(G868), .A2(G301), .ZN(n596) );
  NAND2_X1 U669 ( .A1(G79), .A2(n643), .ZN(n589) );
  NAND2_X1 U670 ( .A1(G54), .A2(n637), .ZN(n588) );
  NAND2_X1 U671 ( .A1(n589), .A2(n588), .ZN(n593) );
  NAND2_X1 U672 ( .A1(G66), .A2(n639), .ZN(n591) );
  NAND2_X1 U673 ( .A1(G92), .A2(n640), .ZN(n590) );
  NAND2_X1 U674 ( .A1(n591), .A2(n590), .ZN(n592) );
  NOR2_X1 U675 ( .A1(n593), .A2(n592), .ZN(n594) );
  XOR2_X1 U676 ( .A(KEYINPUT15), .B(n594), .Z(n918) );
  OR2_X1 U677 ( .A1(n918), .A2(G868), .ZN(n595) );
  NAND2_X1 U678 ( .A1(n596), .A2(n595), .ZN(G284) );
  NOR2_X1 U679 ( .A1(G868), .A2(G299), .ZN(n597) );
  XNOR2_X1 U680 ( .A(n597), .B(KEYINPUT72), .ZN(n599) );
  INV_X1 U681 ( .A(G868), .ZN(n649) );
  NOR2_X1 U682 ( .A1(n649), .A2(G286), .ZN(n598) );
  NOR2_X1 U683 ( .A1(n599), .A2(n598), .ZN(G297) );
  NAND2_X1 U684 ( .A1(n600), .A2(G559), .ZN(n601) );
  NAND2_X1 U685 ( .A1(n601), .A2(n918), .ZN(n602) );
  XNOR2_X1 U686 ( .A(n602), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U687 ( .A1(G868), .A2(n923), .ZN(n605) );
  NAND2_X1 U688 ( .A1(G868), .A2(n918), .ZN(n603) );
  NOR2_X1 U689 ( .A1(G559), .A2(n603), .ZN(n604) );
  NOR2_X1 U690 ( .A1(n605), .A2(n604), .ZN(G282) );
  NAND2_X1 U691 ( .A1(n918), .A2(G559), .ZN(n659) );
  XNOR2_X1 U692 ( .A(n923), .B(n659), .ZN(n606) );
  NOR2_X1 U693 ( .A1(G860), .A2(n606), .ZN(n616) );
  NAND2_X1 U694 ( .A1(G67), .A2(n639), .ZN(n608) );
  NAND2_X1 U695 ( .A1(G55), .A2(n637), .ZN(n607) );
  NAND2_X1 U696 ( .A1(n608), .A2(n607), .ZN(n614) );
  NAND2_X1 U697 ( .A1(n640), .A2(G93), .ZN(n609) );
  XNOR2_X1 U698 ( .A(n609), .B(KEYINPUT76), .ZN(n611) );
  NAND2_X1 U699 ( .A1(G80), .A2(n643), .ZN(n610) );
  NAND2_X1 U700 ( .A1(n611), .A2(n610), .ZN(n612) );
  XOR2_X1 U701 ( .A(KEYINPUT77), .B(n612), .Z(n613) );
  NOR2_X1 U702 ( .A1(n614), .A2(n613), .ZN(n653) );
  XNOR2_X1 U703 ( .A(n653), .B(KEYINPUT78), .ZN(n615) );
  XNOR2_X1 U704 ( .A(n616), .B(n615), .ZN(G145) );
  NAND2_X1 U705 ( .A1(G88), .A2(n640), .ZN(n617) );
  XOR2_X1 U706 ( .A(KEYINPUT82), .B(n617), .Z(n622) );
  NAND2_X1 U707 ( .A1(G62), .A2(n639), .ZN(n619) );
  NAND2_X1 U708 ( .A1(G50), .A2(n637), .ZN(n618) );
  NAND2_X1 U709 ( .A1(n619), .A2(n618), .ZN(n620) );
  XOR2_X1 U710 ( .A(KEYINPUT81), .B(n620), .Z(n621) );
  NOR2_X1 U711 ( .A1(n622), .A2(n621), .ZN(n624) );
  NAND2_X1 U712 ( .A1(G75), .A2(n643), .ZN(n623) );
  NAND2_X1 U713 ( .A1(n624), .A2(n623), .ZN(G303) );
  INV_X1 U714 ( .A(G303), .ZN(G166) );
  NAND2_X1 U715 ( .A1(G651), .A2(G74), .ZN(n626) );
  NAND2_X1 U716 ( .A1(G49), .A2(n637), .ZN(n625) );
  NAND2_X1 U717 ( .A1(n626), .A2(n625), .ZN(n627) );
  XOR2_X1 U718 ( .A(KEYINPUT79), .B(n627), .Z(n628) );
  NOR2_X1 U719 ( .A1(n639), .A2(n628), .ZN(n630) );
  NAND2_X1 U720 ( .A1(n534), .A2(G87), .ZN(n629) );
  NAND2_X1 U721 ( .A1(n630), .A2(n629), .ZN(G288) );
  AND2_X1 U722 ( .A1(n639), .A2(G60), .ZN(n634) );
  NAND2_X1 U723 ( .A1(G85), .A2(n640), .ZN(n632) );
  NAND2_X1 U724 ( .A1(G47), .A2(n637), .ZN(n631) );
  NAND2_X1 U725 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U726 ( .A1(n634), .A2(n633), .ZN(n636) );
  NAND2_X1 U727 ( .A1(G72), .A2(n643), .ZN(n635) );
  NAND2_X1 U728 ( .A1(n636), .A2(n635), .ZN(G290) );
  NAND2_X1 U729 ( .A1(n637), .A2(G48), .ZN(n638) );
  XNOR2_X1 U730 ( .A(n638), .B(KEYINPUT80), .ZN(n648) );
  NAND2_X1 U731 ( .A1(G61), .A2(n639), .ZN(n642) );
  NAND2_X1 U732 ( .A1(G86), .A2(n640), .ZN(n641) );
  NAND2_X1 U733 ( .A1(n642), .A2(n641), .ZN(n646) );
  NAND2_X1 U734 ( .A1(n643), .A2(G73), .ZN(n644) );
  XOR2_X1 U735 ( .A(KEYINPUT2), .B(n644), .Z(n645) );
  NOR2_X1 U736 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U737 ( .A1(n648), .A2(n647), .ZN(G305) );
  NAND2_X1 U738 ( .A1(n649), .A2(n653), .ZN(n662) );
  INV_X1 U739 ( .A(G299), .ZN(n917) );
  XNOR2_X1 U740 ( .A(G166), .B(G288), .ZN(n656) );
  XNOR2_X1 U741 ( .A(KEYINPUT84), .B(KEYINPUT83), .ZN(n651) );
  XNOR2_X1 U742 ( .A(n923), .B(KEYINPUT19), .ZN(n650) );
  XNOR2_X1 U743 ( .A(n651), .B(n650), .ZN(n652) );
  XNOR2_X1 U744 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U745 ( .A(n654), .B(G290), .ZN(n655) );
  XNOR2_X1 U746 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U747 ( .A(n917), .B(n657), .ZN(n658) );
  XNOR2_X1 U748 ( .A(n658), .B(G305), .ZN(n905) );
  XNOR2_X1 U749 ( .A(n905), .B(n659), .ZN(n660) );
  NAND2_X1 U750 ( .A1(n660), .A2(G868), .ZN(n661) );
  NAND2_X1 U751 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U752 ( .A(n663), .B(KEYINPUT85), .ZN(G295) );
  NAND2_X1 U753 ( .A1(G2078), .A2(G2084), .ZN(n664) );
  XOR2_X1 U754 ( .A(KEYINPUT20), .B(n664), .Z(n665) );
  NAND2_X1 U755 ( .A1(G2090), .A2(n665), .ZN(n666) );
  XNOR2_X1 U756 ( .A(KEYINPUT21), .B(n666), .ZN(n667) );
  NAND2_X1 U757 ( .A1(n667), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U758 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U759 ( .A1(G220), .A2(G219), .ZN(n668) );
  XOR2_X1 U760 ( .A(KEYINPUT22), .B(n668), .Z(n669) );
  NOR2_X1 U761 ( .A1(G218), .A2(n669), .ZN(n670) );
  NAND2_X1 U762 ( .A1(G96), .A2(n670), .ZN(n840) );
  NAND2_X1 U763 ( .A1(G2106), .A2(n840), .ZN(n671) );
  XOR2_X1 U764 ( .A(KEYINPUT86), .B(n671), .Z(n677) );
  NAND2_X1 U765 ( .A1(G120), .A2(G69), .ZN(n672) );
  NOR2_X1 U766 ( .A1(G237), .A2(n672), .ZN(n673) );
  XNOR2_X1 U767 ( .A(n673), .B(KEYINPUT87), .ZN(n674) );
  NOR2_X1 U768 ( .A1(G238), .A2(n674), .ZN(n842) );
  NOR2_X1 U769 ( .A1(n842), .A2(n675), .ZN(n676) );
  NOR2_X1 U770 ( .A1(n677), .A2(n676), .ZN(G319) );
  INV_X1 U771 ( .A(G319), .ZN(n679) );
  NAND2_X1 U772 ( .A1(G483), .A2(G661), .ZN(n678) );
  NOR2_X1 U773 ( .A1(n679), .A2(n678), .ZN(n839) );
  NAND2_X1 U774 ( .A1(n839), .A2(G36), .ZN(G176) );
  XNOR2_X1 U775 ( .A(G1986), .B(G290), .ZN(n920) );
  AND2_X1 U776 ( .A1(G40), .A2(n680), .ZN(n681) );
  AND2_X1 U777 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U778 ( .A1(n684), .A2(n683), .ZN(n717) );
  NOR2_X1 U779 ( .A1(n716), .A2(n717), .ZN(n821) );
  NAND2_X1 U780 ( .A1(n920), .A2(n821), .ZN(n809) );
  NAND2_X1 U781 ( .A1(n881), .A2(G104), .ZN(n685) );
  XNOR2_X1 U782 ( .A(n685), .B(KEYINPUT88), .ZN(n687) );
  NAND2_X1 U783 ( .A1(G140), .A2(n882), .ZN(n686) );
  NAND2_X1 U784 ( .A1(n687), .A2(n686), .ZN(n689) );
  XOR2_X1 U785 ( .A(KEYINPUT34), .B(KEYINPUT89), .Z(n688) );
  XNOR2_X1 U786 ( .A(n689), .B(n688), .ZN(n695) );
  NAND2_X1 U787 ( .A1(n878), .A2(G128), .ZN(n690) );
  XNOR2_X1 U788 ( .A(n690), .B(KEYINPUT90), .ZN(n692) );
  NAND2_X1 U789 ( .A1(G116), .A2(n877), .ZN(n691) );
  NAND2_X1 U790 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U791 ( .A(KEYINPUT35), .B(n693), .Z(n694) );
  NOR2_X1 U792 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U793 ( .A(KEYINPUT36), .B(n696), .Z(n901) );
  XOR2_X1 U794 ( .A(KEYINPUT37), .B(G2067), .Z(n819) );
  NAND2_X1 U795 ( .A1(n901), .A2(n819), .ZN(n697) );
  XNOR2_X1 U796 ( .A(KEYINPUT91), .B(n697), .ZN(n1003) );
  NAND2_X1 U797 ( .A1(n821), .A2(n1003), .ZN(n817) );
  NAND2_X1 U798 ( .A1(G95), .A2(n881), .ZN(n699) );
  NAND2_X1 U799 ( .A1(G131), .A2(n882), .ZN(n698) );
  NAND2_X1 U800 ( .A1(n699), .A2(n698), .ZN(n703) );
  NAND2_X1 U801 ( .A1(G107), .A2(n877), .ZN(n701) );
  NAND2_X1 U802 ( .A1(G119), .A2(n878), .ZN(n700) );
  NAND2_X1 U803 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U804 ( .A1(n703), .A2(n702), .ZN(n890) );
  INV_X1 U805 ( .A(G1991), .ZN(n810) );
  NOR2_X1 U806 ( .A1(n890), .A2(n810), .ZN(n713) );
  NAND2_X1 U807 ( .A1(G141), .A2(n882), .ZN(n704) );
  XNOR2_X1 U808 ( .A(n704), .B(KEYINPUT92), .ZN(n711) );
  NAND2_X1 U809 ( .A1(G117), .A2(n877), .ZN(n706) );
  NAND2_X1 U810 ( .A1(G129), .A2(n878), .ZN(n705) );
  NAND2_X1 U811 ( .A1(n706), .A2(n705), .ZN(n709) );
  NAND2_X1 U812 ( .A1(n881), .A2(G105), .ZN(n707) );
  XOR2_X1 U813 ( .A(KEYINPUT38), .B(n707), .Z(n708) );
  NOR2_X1 U814 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U815 ( .A1(n711), .A2(n710), .ZN(n899) );
  AND2_X1 U816 ( .A1(n899), .A2(G1996), .ZN(n712) );
  NOR2_X1 U817 ( .A1(n713), .A2(n712), .ZN(n1013) );
  INV_X1 U818 ( .A(n821), .ZN(n714) );
  NOR2_X1 U819 ( .A1(n1013), .A2(n714), .ZN(n814) );
  INV_X1 U820 ( .A(n814), .ZN(n715) );
  NAND2_X1 U821 ( .A1(n817), .A2(n715), .ZN(n807) );
  INV_X1 U822 ( .A(n716), .ZN(n718) );
  NOR2_X2 U823 ( .A1(n718), .A2(n717), .ZN(n746) );
  INV_X1 U824 ( .A(n746), .ZN(n764) );
  NAND2_X1 U825 ( .A1(G1956), .A2(n764), .ZN(n722) );
  INV_X1 U826 ( .A(KEYINPUT27), .ZN(n720) );
  NAND2_X1 U827 ( .A1(n746), .A2(G2072), .ZN(n719) );
  XNOR2_X1 U828 ( .A(n720), .B(n719), .ZN(n721) );
  NAND2_X1 U829 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U830 ( .A(n723), .B(KEYINPUT94), .Z(n738) );
  NOR2_X1 U831 ( .A1(n917), .A2(n738), .ZN(n724) );
  XOR2_X1 U832 ( .A(n724), .B(KEYINPUT28), .Z(n742) );
  NAND2_X1 U833 ( .A1(n764), .A2(G1341), .ZN(n726) );
  INV_X1 U834 ( .A(n923), .ZN(n725) );
  NAND2_X1 U835 ( .A1(n726), .A2(n725), .ZN(n730) );
  INV_X1 U836 ( .A(G1996), .ZN(n946) );
  NOR2_X1 U837 ( .A1(n764), .A2(n946), .ZN(n728) );
  XOR2_X1 U838 ( .A(KEYINPUT26), .B(KEYINPUT95), .Z(n727) );
  XNOR2_X1 U839 ( .A(n728), .B(n727), .ZN(n729) );
  NOR2_X1 U840 ( .A1(n730), .A2(n729), .ZN(n732) );
  NOR2_X1 U841 ( .A1(n732), .A2(n918), .ZN(n731) );
  NAND2_X1 U842 ( .A1(n732), .A2(n918), .ZN(n736) );
  NOR2_X1 U843 ( .A1(n746), .A2(G1348), .ZN(n734) );
  NOR2_X1 U844 ( .A1(G2067), .A2(n764), .ZN(n733) );
  NOR2_X1 U845 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U846 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U847 ( .A1(n517), .A2(n737), .ZN(n740) );
  NAND2_X1 U848 ( .A1(n917), .A2(n738), .ZN(n739) );
  NAND2_X1 U849 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U850 ( .A1(n742), .A2(n741), .ZN(n745) );
  XOR2_X1 U851 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n743) );
  NAND2_X1 U852 ( .A1(G1961), .A2(n764), .ZN(n748) );
  XOR2_X1 U853 ( .A(G2078), .B(KEYINPUT25), .Z(n948) );
  NAND2_X1 U854 ( .A1(n746), .A2(n948), .ZN(n747) );
  NAND2_X1 U855 ( .A1(n748), .A2(n747), .ZN(n755) );
  NOR2_X1 U856 ( .A1(G301), .A2(n755), .ZN(n749) );
  NAND2_X1 U857 ( .A1(n764), .A2(G8), .ZN(n751) );
  NOR2_X1 U858 ( .A1(G1966), .A2(n788), .ZN(n778) );
  NOR2_X1 U859 ( .A1(G2084), .A2(n764), .ZN(n774) );
  NOR2_X1 U860 ( .A1(n778), .A2(n774), .ZN(n752) );
  NAND2_X1 U861 ( .A1(G8), .A2(n752), .ZN(n753) );
  XNOR2_X1 U862 ( .A(KEYINPUT30), .B(n753), .ZN(n754) );
  NOR2_X1 U863 ( .A1(n754), .A2(G168), .ZN(n758) );
  NAND2_X1 U864 ( .A1(G301), .A2(n755), .ZN(n756) );
  XNOR2_X1 U865 ( .A(n756), .B(KEYINPUT99), .ZN(n757) );
  NOR2_X1 U866 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U867 ( .A(n759), .B(KEYINPUT31), .ZN(n760) );
  NOR2_X1 U868 ( .A1(n761), .A2(n760), .ZN(n763) );
  XNOR2_X1 U869 ( .A(n763), .B(n762), .ZN(n776) );
  NAND2_X1 U870 ( .A1(n776), .A2(G286), .ZN(n770) );
  NOR2_X1 U871 ( .A1(G2090), .A2(n764), .ZN(n765) );
  XNOR2_X1 U872 ( .A(KEYINPUT101), .B(n765), .ZN(n768) );
  NOR2_X1 U873 ( .A1(G1971), .A2(n788), .ZN(n766) );
  NOR2_X1 U874 ( .A1(G166), .A2(n766), .ZN(n767) );
  NAND2_X1 U875 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U876 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U877 ( .A1(n771), .A2(G8), .ZN(n773) );
  NAND2_X1 U878 ( .A1(G8), .A2(n774), .ZN(n775) );
  NAND2_X1 U879 ( .A1(n776), .A2(n775), .ZN(n777) );
  NOR2_X1 U880 ( .A1(n778), .A2(n777), .ZN(n779) );
  INV_X1 U881 ( .A(n800), .ZN(n784) );
  NOR2_X1 U882 ( .A1(G1976), .A2(G288), .ZN(n785) );
  NOR2_X1 U883 ( .A1(G1971), .A2(G303), .ZN(n781) );
  NOR2_X1 U884 ( .A1(n785), .A2(n781), .ZN(n927) );
  INV_X1 U885 ( .A(KEYINPUT33), .ZN(n782) );
  AND2_X1 U886 ( .A1(n927), .A2(n782), .ZN(n783) );
  AND2_X1 U887 ( .A1(n784), .A2(n783), .ZN(n794) );
  AND2_X1 U888 ( .A1(n785), .A2(KEYINPUT33), .ZN(n786) );
  INV_X1 U889 ( .A(n788), .ZN(n801) );
  NAND2_X1 U890 ( .A1(n786), .A2(n801), .ZN(n792) );
  NAND2_X1 U891 ( .A1(G1976), .A2(G288), .ZN(n926) );
  INV_X1 U892 ( .A(n926), .ZN(n787) );
  NOR2_X1 U893 ( .A1(KEYINPUT33), .A2(n789), .ZN(n790) );
  XNOR2_X1 U894 ( .A(G1981), .B(G305), .ZN(n937) );
  NOR2_X1 U895 ( .A1(n790), .A2(n937), .ZN(n791) );
  NAND2_X1 U896 ( .A1(n792), .A2(n791), .ZN(n793) );
  NOR2_X1 U897 ( .A1(n794), .A2(n793), .ZN(n805) );
  NOR2_X1 U898 ( .A1(G1981), .A2(G305), .ZN(n795) );
  XNOR2_X1 U899 ( .A(n795), .B(KEYINPUT24), .ZN(n796) );
  NAND2_X1 U900 ( .A1(G8), .A2(G166), .ZN(n797) );
  NOR2_X1 U901 ( .A1(G2090), .A2(n797), .ZN(n798) );
  XNOR2_X1 U902 ( .A(n798), .B(KEYINPUT102), .ZN(n799) );
  NOR2_X1 U903 ( .A1(n802), .A2(n801), .ZN(n803) );
  NOR2_X1 U904 ( .A1(n805), .A2(n804), .ZN(n806) );
  NOR2_X1 U905 ( .A1(n807), .A2(n806), .ZN(n808) );
  NAND2_X1 U906 ( .A1(n809), .A2(n808), .ZN(n824) );
  NOR2_X1 U907 ( .A1(G1996), .A2(n899), .ZN(n1005) );
  AND2_X1 U908 ( .A1(n810), .A2(n890), .ZN(n1010) );
  NOR2_X1 U909 ( .A1(G1986), .A2(G290), .ZN(n811) );
  XOR2_X1 U910 ( .A(n811), .B(KEYINPUT103), .Z(n812) );
  NOR2_X1 U911 ( .A1(n1010), .A2(n812), .ZN(n813) );
  NOR2_X1 U912 ( .A1(n814), .A2(n813), .ZN(n815) );
  NOR2_X1 U913 ( .A1(n1005), .A2(n815), .ZN(n816) );
  XNOR2_X1 U914 ( .A(KEYINPUT39), .B(n816), .ZN(n818) );
  NAND2_X1 U915 ( .A1(n818), .A2(n817), .ZN(n820) );
  OR2_X1 U916 ( .A1(n901), .A2(n819), .ZN(n1000) );
  NAND2_X1 U917 ( .A1(n820), .A2(n1000), .ZN(n822) );
  NAND2_X1 U918 ( .A1(n822), .A2(n821), .ZN(n823) );
  NAND2_X1 U919 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U920 ( .A(n825), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U921 ( .A(G2454), .B(G2435), .ZN(n834) );
  XNOR2_X1 U922 ( .A(KEYINPUT104), .B(G2427), .ZN(n832) );
  XOR2_X1 U923 ( .A(G2430), .B(G2446), .Z(n827) );
  XNOR2_X1 U924 ( .A(G2443), .B(G2451), .ZN(n826) );
  XNOR2_X1 U925 ( .A(n827), .B(n826), .ZN(n828) );
  XOR2_X1 U926 ( .A(n828), .B(G2438), .Z(n830) );
  XNOR2_X1 U927 ( .A(G1348), .B(G1341), .ZN(n829) );
  XNOR2_X1 U928 ( .A(n830), .B(n829), .ZN(n831) );
  XNOR2_X1 U929 ( .A(n832), .B(n831), .ZN(n833) );
  XNOR2_X1 U930 ( .A(n834), .B(n833), .ZN(n835) );
  NAND2_X1 U931 ( .A1(n835), .A2(G14), .ZN(n910) );
  XNOR2_X1 U932 ( .A(KEYINPUT105), .B(n910), .ZN(G401) );
  INV_X1 U933 ( .A(G223), .ZN(n836) );
  NAND2_X1 U934 ( .A1(G2106), .A2(n836), .ZN(G217) );
  AND2_X1 U935 ( .A1(G15), .A2(G2), .ZN(n837) );
  NAND2_X1 U936 ( .A1(G661), .A2(n837), .ZN(G259) );
  NAND2_X1 U937 ( .A1(G3), .A2(G1), .ZN(n838) );
  NAND2_X1 U938 ( .A1(n839), .A2(n838), .ZN(G188) );
  XOR2_X1 U939 ( .A(G120), .B(KEYINPUT106), .Z(G236) );
  XNOR2_X1 U940 ( .A(G69), .B(KEYINPUT107), .ZN(G235) );
  INV_X1 U942 ( .A(G96), .ZN(G221) );
  INV_X1 U943 ( .A(n840), .ZN(n841) );
  NAND2_X1 U944 ( .A1(n842), .A2(n841), .ZN(G261) );
  INV_X1 U945 ( .A(G261), .ZN(G325) );
  XOR2_X1 U946 ( .A(G2100), .B(G2096), .Z(n844) );
  XNOR2_X1 U947 ( .A(KEYINPUT42), .B(G2678), .ZN(n843) );
  XNOR2_X1 U948 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U949 ( .A(KEYINPUT43), .B(G2090), .Z(n846) );
  XNOR2_X1 U950 ( .A(G2067), .B(G2072), .ZN(n845) );
  XNOR2_X1 U951 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U952 ( .A(n848), .B(n847), .Z(n850) );
  XNOR2_X1 U953 ( .A(G2078), .B(G2084), .ZN(n849) );
  XNOR2_X1 U954 ( .A(n850), .B(n849), .ZN(G227) );
  XOR2_X1 U955 ( .A(KEYINPUT109), .B(G1976), .Z(n852) );
  XNOR2_X1 U956 ( .A(G1966), .B(G1981), .ZN(n851) );
  XNOR2_X1 U957 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U958 ( .A(n853), .B(KEYINPUT41), .Z(n855) );
  XNOR2_X1 U959 ( .A(G1996), .B(G1991), .ZN(n854) );
  XNOR2_X1 U960 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U961 ( .A(G1971), .B(G1956), .Z(n857) );
  XNOR2_X1 U962 ( .A(G1986), .B(G1961), .ZN(n856) );
  XNOR2_X1 U963 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U964 ( .A(n859), .B(n858), .Z(n861) );
  XNOR2_X1 U965 ( .A(KEYINPUT108), .B(G2474), .ZN(n860) );
  XNOR2_X1 U966 ( .A(n861), .B(n860), .ZN(G229) );
  NAND2_X1 U967 ( .A1(G124), .A2(n878), .ZN(n862) );
  XNOR2_X1 U968 ( .A(n862), .B(KEYINPUT44), .ZN(n863) );
  XNOR2_X1 U969 ( .A(n863), .B(KEYINPUT110), .ZN(n865) );
  NAND2_X1 U970 ( .A1(G112), .A2(n877), .ZN(n864) );
  NAND2_X1 U971 ( .A1(n865), .A2(n864), .ZN(n869) );
  NAND2_X1 U972 ( .A1(G100), .A2(n881), .ZN(n867) );
  NAND2_X1 U973 ( .A1(G136), .A2(n882), .ZN(n866) );
  NAND2_X1 U974 ( .A1(n867), .A2(n866), .ZN(n868) );
  NOR2_X1 U975 ( .A1(n869), .A2(n868), .ZN(G162) );
  NAND2_X1 U976 ( .A1(G103), .A2(n881), .ZN(n871) );
  NAND2_X1 U977 ( .A1(G139), .A2(n882), .ZN(n870) );
  NAND2_X1 U978 ( .A1(n871), .A2(n870), .ZN(n876) );
  NAND2_X1 U979 ( .A1(G115), .A2(n877), .ZN(n873) );
  NAND2_X1 U980 ( .A1(G127), .A2(n878), .ZN(n872) );
  NAND2_X1 U981 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U982 ( .A(KEYINPUT47), .B(n874), .Z(n875) );
  NOR2_X1 U983 ( .A1(n876), .A2(n875), .ZN(n996) );
  XNOR2_X1 U984 ( .A(n996), .B(G162), .ZN(n889) );
  NAND2_X1 U985 ( .A1(G118), .A2(n877), .ZN(n880) );
  NAND2_X1 U986 ( .A1(G130), .A2(n878), .ZN(n879) );
  NAND2_X1 U987 ( .A1(n880), .A2(n879), .ZN(n887) );
  NAND2_X1 U988 ( .A1(G106), .A2(n881), .ZN(n884) );
  NAND2_X1 U989 ( .A1(G142), .A2(n882), .ZN(n883) );
  NAND2_X1 U990 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U991 ( .A(KEYINPUT45), .B(n885), .Z(n886) );
  NOR2_X1 U992 ( .A1(n887), .A2(n886), .ZN(n888) );
  XNOR2_X1 U993 ( .A(n889), .B(n888), .ZN(n893) );
  XNOR2_X1 U994 ( .A(G164), .B(n890), .ZN(n891) );
  XNOR2_X1 U995 ( .A(n891), .B(n1009), .ZN(n892) );
  XOR2_X1 U996 ( .A(n893), .B(n892), .Z(n898) );
  XOR2_X1 U997 ( .A(KEYINPUT112), .B(KEYINPUT48), .Z(n895) );
  XNOR2_X1 U998 ( .A(KEYINPUT113), .B(KEYINPUT46), .ZN(n894) );
  XNOR2_X1 U999 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U1000 ( .A(KEYINPUT111), .B(n896), .ZN(n897) );
  XNOR2_X1 U1001 ( .A(n898), .B(n897), .ZN(n900) );
  XNOR2_X1 U1002 ( .A(n900), .B(n899), .ZN(n903) );
  XNOR2_X1 U1003 ( .A(G160), .B(n901), .ZN(n902) );
  XNOR2_X1 U1004 ( .A(n903), .B(n902), .ZN(n904) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n904), .ZN(G395) );
  XNOR2_X1 U1006 ( .A(n905), .B(KEYINPUT114), .ZN(n907) );
  XNOR2_X1 U1007 ( .A(n918), .B(G286), .ZN(n906) );
  XNOR2_X1 U1008 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1009 ( .A(G171), .B(n908), .ZN(n909) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n909), .ZN(G397) );
  NAND2_X1 U1011 ( .A1(G319), .A2(n910), .ZN(n914) );
  NOR2_X1 U1012 ( .A1(G227), .A2(G229), .ZN(n911) );
  XOR2_X1 U1013 ( .A(KEYINPUT115), .B(n911), .Z(n912) );
  XNOR2_X1 U1014 ( .A(n912), .B(KEYINPUT49), .ZN(n913) );
  NOR2_X1 U1015 ( .A1(n914), .A2(n913), .ZN(n916) );
  NOR2_X1 U1016 ( .A1(G395), .A2(G397), .ZN(n915) );
  NAND2_X1 U1017 ( .A1(n916), .A2(n915), .ZN(G225) );
  INV_X1 U1018 ( .A(G225), .ZN(G308) );
  XNOR2_X1 U1019 ( .A(n917), .B(G1956), .ZN(n922) );
  XOR2_X1 U1020 ( .A(G1348), .B(n918), .Z(n919) );
  NOR2_X1 U1021 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1022 ( .A1(n922), .A2(n921), .ZN(n934) );
  XNOR2_X1 U1023 ( .A(G301), .B(G1961), .ZN(n925) );
  XNOR2_X1 U1024 ( .A(n923), .B(G1341), .ZN(n924) );
  NOR2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(n932) );
  AND2_X1 U1026 ( .A1(G303), .A2(G1971), .ZN(n929) );
  NAND2_X1 U1027 ( .A1(n927), .A2(n926), .ZN(n928) );
  NOR2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1029 ( .A(n930), .B(KEYINPUT120), .ZN(n931) );
  NAND2_X1 U1030 ( .A1(n932), .A2(n931), .ZN(n933) );
  NOR2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1032 ( .A(KEYINPUT121), .B(n935), .ZN(n940) );
  XOR2_X1 U1033 ( .A(G1966), .B(G168), .Z(n936) );
  NOR2_X1 U1034 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1035 ( .A(KEYINPUT57), .B(n938), .ZN(n939) );
  NOR2_X1 U1036 ( .A1(n940), .A2(n939), .ZN(n942) );
  XOR2_X1 U1037 ( .A(KEYINPUT56), .B(G16), .Z(n941) );
  NOR2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n943) );
  XOR2_X1 U1039 ( .A(KEYINPUT122), .B(n943), .Z(n994) );
  XNOR2_X1 U1040 ( .A(G2067), .B(G26), .ZN(n945) );
  XNOR2_X1 U1041 ( .A(G33), .B(G2072), .ZN(n944) );
  NOR2_X1 U1042 ( .A1(n945), .A2(n944), .ZN(n953) );
  XNOR2_X1 U1043 ( .A(G32), .B(n946), .ZN(n947) );
  NAND2_X1 U1044 ( .A1(n947), .A2(G28), .ZN(n951) );
  XNOR2_X1 U1045 ( .A(G27), .B(n948), .ZN(n949) );
  XNOR2_X1 U1046 ( .A(KEYINPUT118), .B(n949), .ZN(n950) );
  NOR2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1048 ( .A1(n953), .A2(n952), .ZN(n955) );
  XNOR2_X1 U1049 ( .A(G25), .B(G1991), .ZN(n954) );
  NOR2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n956) );
  XOR2_X1 U1051 ( .A(KEYINPUT53), .B(n956), .Z(n960) );
  XNOR2_X1 U1052 ( .A(KEYINPUT54), .B(KEYINPUT119), .ZN(n957) );
  XNOR2_X1 U1053 ( .A(n957), .B(G34), .ZN(n958) );
  XNOR2_X1 U1054 ( .A(G2084), .B(n958), .ZN(n959) );
  NAND2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n962) );
  XNOR2_X1 U1056 ( .A(G35), .B(G2090), .ZN(n961) );
  NOR2_X1 U1057 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1058 ( .A(KEYINPUT55), .B(n963), .Z(n964) );
  NOR2_X1 U1059 ( .A1(G29), .A2(n964), .ZN(n992) );
  XOR2_X1 U1060 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n987) );
  XNOR2_X1 U1061 ( .A(G1348), .B(KEYINPUT59), .ZN(n965) );
  XNOR2_X1 U1062 ( .A(n965), .B(G4), .ZN(n969) );
  XNOR2_X1 U1063 ( .A(G1341), .B(G19), .ZN(n967) );
  XNOR2_X1 U1064 ( .A(G1956), .B(G20), .ZN(n966) );
  NOR2_X1 U1065 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1066 ( .A1(n969), .A2(n968), .ZN(n972) );
  XOR2_X1 U1067 ( .A(KEYINPUT123), .B(G1981), .Z(n970) );
  XNOR2_X1 U1068 ( .A(G6), .B(n970), .ZN(n971) );
  NOR2_X1 U1069 ( .A1(n972), .A2(n971), .ZN(n973) );
  XOR2_X1 U1070 ( .A(KEYINPUT60), .B(n973), .Z(n975) );
  XNOR2_X1 U1071 ( .A(G1966), .B(G21), .ZN(n974) );
  NOR2_X1 U1072 ( .A1(n975), .A2(n974), .ZN(n985) );
  XNOR2_X1 U1073 ( .A(G1971), .B(G22), .ZN(n977) );
  XNOR2_X1 U1074 ( .A(G1976), .B(G23), .ZN(n976) );
  NOR2_X1 U1075 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1076 ( .A(KEYINPUT124), .B(n978), .Z(n980) );
  XNOR2_X1 U1077 ( .A(G1986), .B(G24), .ZN(n979) );
  NOR2_X1 U1078 ( .A1(n980), .A2(n979), .ZN(n981) );
  XOR2_X1 U1079 ( .A(KEYINPUT58), .B(n981), .Z(n983) );
  XNOR2_X1 U1080 ( .A(G1961), .B(G5), .ZN(n982) );
  NOR2_X1 U1081 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1082 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1083 ( .A(n987), .B(n986), .ZN(n988) );
  NOR2_X1 U1084 ( .A1(G16), .A2(n988), .ZN(n989) );
  XOR2_X1 U1085 ( .A(KEYINPUT126), .B(n989), .Z(n990) );
  NAND2_X1 U1086 ( .A1(G11), .A2(n990), .ZN(n991) );
  NOR2_X1 U1087 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1088 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1089 ( .A(n995), .B(KEYINPUT127), .ZN(n1024) );
  XOR2_X1 U1090 ( .A(G2072), .B(n996), .Z(n998) );
  XOR2_X1 U1091 ( .A(G164), .B(G2078), .Z(n997) );
  NOR2_X1 U1092 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1093 ( .A(n999), .B(KEYINPUT50), .ZN(n1001) );
  NAND2_X1 U1094 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NOR2_X1 U1095 ( .A1(n1003), .A2(n1002), .ZN(n1017) );
  XNOR2_X1 U1096 ( .A(G160), .B(G2084), .ZN(n1008) );
  XOR2_X1 U1097 ( .A(G2090), .B(G162), .Z(n1004) );
  NOR2_X1 U1098 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1099 ( .A(KEYINPUT51), .B(n1006), .Z(n1007) );
  NAND2_X1 U1100 ( .A1(n1008), .A2(n1007), .ZN(n1015) );
  NOR2_X1 U1101 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1102 ( .A(n1011), .B(KEYINPUT116), .ZN(n1012) );
  NAND2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1106 ( .A(KEYINPUT52), .B(n1018), .ZN(n1019) );
  XNOR2_X1 U1107 ( .A(KEYINPUT117), .B(n1019), .ZN(n1021) );
  INV_X1 U1108 ( .A(KEYINPUT55), .ZN(n1020) );
  NAND2_X1 U1109 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1110 ( .A1(n1022), .A2(G29), .ZN(n1023) );
  NAND2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XOR2_X1 U1112 ( .A(KEYINPUT62), .B(n1025), .Z(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
endmodule

