//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0 1 0 1 1 0 0 1 0 1 1 1 1 1 0 1 1 1 1 0 0 0 0 1 0 0 1 0 0 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:05 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n596,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n857, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G146), .ZN(new_n187));
  INV_X1    g001(.A(G143), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT1), .ZN(new_n190));
  OAI21_X1  g004(.A(G128), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n188), .A2(G146), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n192), .B1(new_n187), .B2(new_n188), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n191), .A2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n188), .A2(G146), .ZN(new_n196));
  INV_X1    g010(.A(G128), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(KEYINPUT1), .ZN(new_n198));
  OAI211_X1 g012(.A(new_n196), .B(new_n198), .C1(new_n187), .C2(new_n188), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n195), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G134), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT65), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT65), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G134), .ZN(new_n204));
  INV_X1    g018(.A(G137), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n202), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT11), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(KEYINPUT66), .ZN(new_n209));
  INV_X1    g023(.A(G131), .ZN(new_n210));
  NOR3_X1   g024(.A1(new_n207), .A2(new_n201), .A3(G137), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n202), .A2(new_n204), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n211), .B1(new_n212), .B2(G137), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT66), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n206), .A2(new_n214), .A3(new_n207), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n209), .A2(new_n210), .A3(new_n213), .A4(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n206), .B1(G134), .B2(new_n205), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G131), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n200), .A2(new_n216), .A3(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n221));
  AND3_X1   g035(.A1(new_n206), .A2(new_n214), .A3(new_n207), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n214), .B1(new_n206), .B2(new_n207), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n210), .B1(new_n224), .B2(new_n213), .ZN(new_n225));
  INV_X1    g039(.A(new_n216), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n221), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n209), .A2(new_n213), .A3(new_n215), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G131), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n229), .A2(KEYINPUT67), .A3(new_n216), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n189), .B1(new_n188), .B2(G146), .ZN(new_n232));
  AND2_X1   g046(.A1(KEYINPUT0), .A2(G128), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n193), .A2(new_n233), .ZN(new_n234));
  OR2_X1    g048(.A1(KEYINPUT0), .A2(G128), .ZN(new_n235));
  AOI22_X1  g049(.A1(new_n232), .A2(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n220), .B1(new_n231), .B2(new_n236), .ZN(new_n237));
  XOR2_X1   g051(.A(G116), .B(G119), .Z(new_n238));
  XNOR2_X1  g052(.A(KEYINPUT2), .B(G113), .ZN(new_n239));
  XNOR2_X1  g053(.A(new_n238), .B(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n237), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n237), .A2(new_n241), .ZN(new_n244));
  OAI21_X1  g058(.A(KEYINPUT28), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(KEYINPUT28), .B1(new_n237), .B2(new_n241), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G237), .ZN(new_n248));
  INV_X1    g062(.A(G953), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n248), .A2(new_n249), .A3(G210), .ZN(new_n250));
  INV_X1    g064(.A(G101), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n253));
  XOR2_X1   g067(.A(new_n252), .B(new_n253), .Z(new_n254));
  NAND4_X1  g068(.A1(new_n245), .A2(KEYINPUT29), .A3(new_n247), .A4(new_n254), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n255), .B(KEYINPUT71), .ZN(new_n256));
  XNOR2_X1  g070(.A(KEYINPUT72), .B(G902), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n229), .A2(new_n216), .ZN(new_n258));
  AND2_X1   g072(.A1(new_n258), .A2(new_n236), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n240), .B1(new_n259), .B2(new_n220), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT70), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI211_X1 g076(.A(KEYINPUT70), .B(new_n240), .C1(new_n259), .C2(new_n220), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n242), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n246), .B1(new_n264), .B2(KEYINPUT28), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(new_n254), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n229), .A2(KEYINPUT67), .A3(new_n216), .ZN(new_n267));
  AOI21_X1  g081(.A(KEYINPUT67), .B1(new_n229), .B2(new_n216), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n236), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n269), .A2(KEYINPUT30), .A3(new_n219), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT30), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n271), .B1(new_n259), .B2(new_n220), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n270), .A2(new_n240), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n254), .B1(new_n273), .B2(new_n242), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n274), .A2(KEYINPUT29), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n257), .B1(new_n266), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n256), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G472), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT32), .ZN(new_n279));
  INV_X1    g093(.A(new_n254), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n280), .B1(new_n237), .B2(new_n241), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT31), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n273), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n283), .B1(new_n265), .B2(new_n254), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n273), .A2(new_n281), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT68), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n273), .A2(new_n281), .A3(KEYINPUT68), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(KEYINPUT69), .B1(new_n290), .B2(KEYINPUT31), .ZN(new_n291));
  AND3_X1   g105(.A1(new_n273), .A2(new_n281), .A3(KEYINPUT68), .ZN(new_n292));
  AOI21_X1  g106(.A(KEYINPUT68), .B1(new_n273), .B2(new_n281), .ZN(new_n293));
  OAI211_X1 g107(.A(KEYINPUT69), .B(KEYINPUT31), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n285), .B1(new_n291), .B2(new_n295), .ZN(new_n296));
  NOR2_X1   g110(.A1(G472), .A2(G902), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n279), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(KEYINPUT31), .B1(new_n292), .B2(new_n293), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT69), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n284), .B1(new_n301), .B2(new_n294), .ZN(new_n302));
  INV_X1    g116(.A(new_n297), .ZN(new_n303));
  NOR3_X1   g117(.A1(new_n302), .A2(KEYINPUT32), .A3(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n278), .B1(new_n298), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT25), .ZN(new_n306));
  INV_X1    g120(.A(G119), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G128), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n197), .A2(G119), .ZN(new_n309));
  AND2_X1   g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  XOR2_X1   g124(.A(KEYINPUT24), .B(G110), .Z(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G110), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n308), .A2(KEYINPUT23), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n309), .A2(KEYINPUT74), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n314), .B(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G140), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G125), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT75), .B1(new_n318), .B2(KEYINPUT16), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT75), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT16), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n320), .A2(new_n321), .A3(new_n317), .A4(G125), .ZN(new_n322));
  INV_X1    g136(.A(G125), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G140), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n318), .A2(new_n324), .ZN(new_n325));
  OAI211_X1 g139(.A(new_n319), .B(new_n322), .C1(new_n325), .C2(new_n321), .ZN(new_n326));
  INV_X1    g140(.A(G146), .ZN(new_n327));
  AND2_X1   g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n326), .A2(new_n327), .ZN(new_n329));
  OAI221_X1 g143(.A(new_n312), .B1(new_n313), .B2(new_n316), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT76), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n330), .B(new_n331), .ZN(new_n332));
  XOR2_X1   g146(.A(KEYINPUT77), .B(G110), .Z(new_n333));
  NAND2_X1  g147(.A1(new_n316), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n334), .B1(new_n310), .B2(new_n311), .ZN(new_n335));
  INV_X1    g149(.A(new_n325), .ZN(new_n336));
  XOR2_X1   g150(.A(KEYINPUT64), .B(G146), .Z(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n335), .B(new_n338), .C1(new_n327), .C2(new_n326), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n332), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT78), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(KEYINPUT22), .B(G137), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n249), .A2(G221), .A3(G234), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n344), .B(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n347), .B1(new_n340), .B2(KEYINPUT78), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n341), .A2(new_n342), .A3(new_n347), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n257), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n306), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  AOI211_X1 g167(.A(KEYINPUT25), .B(new_n257), .C1(new_n349), .C2(new_n350), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  XOR2_X1   g169(.A(KEYINPUT73), .B(G217), .Z(new_n356));
  AOI21_X1  g170(.A(new_n356), .B1(new_n352), .B2(G234), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n357), .A2(G902), .ZN(new_n358));
  AOI22_X1  g172(.A1(new_n355), .A2(new_n357), .B1(new_n358), .B2(new_n351), .ZN(new_n359));
  INV_X1    g173(.A(G469), .ZN(new_n360));
  XNOR2_X1  g174(.A(KEYINPUT80), .B(G104), .ZN(new_n361));
  OAI21_X1  g175(.A(KEYINPUT3), .B1(new_n361), .B2(G107), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(G107), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT3), .ZN(new_n364));
  INV_X1    g178(.A(G107), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n364), .A2(new_n365), .A3(G104), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n362), .A2(new_n251), .A3(new_n363), .A4(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n361), .A2(G107), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n365), .A2(G104), .ZN(new_n369));
  OAI21_X1  g183(.A(G101), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n192), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n197), .B1(new_n373), .B2(KEYINPUT1), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n199), .B1(new_n232), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT10), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n362), .A2(new_n363), .A3(new_n366), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G101), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n380), .A2(KEYINPUT4), .A3(new_n367), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT4), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n379), .A2(new_n382), .A3(G101), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n381), .A2(new_n236), .A3(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n372), .A2(new_n200), .A3(KEYINPUT10), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n378), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n386), .A2(new_n231), .ZN(new_n387));
  XNOR2_X1  g201(.A(G110), .B(G140), .ZN(new_n388));
  INV_X1    g202(.A(G227), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n389), .A2(G953), .ZN(new_n390));
  XOR2_X1   g204(.A(new_n388), .B(new_n390), .Z(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n387), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n376), .B1(new_n200), .B2(new_n372), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n231), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT12), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n394), .A2(KEYINPUT12), .A3(new_n258), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n393), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n387), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n386), .A2(new_n231), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n391), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n360), .B(new_n352), .C1(new_n400), .C2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT81), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n393), .A2(new_n399), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n401), .A2(new_n402), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n407), .B1(new_n408), .B2(new_n391), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n409), .A2(KEYINPUT81), .A3(new_n360), .A4(new_n352), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n406), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n399), .A2(new_n401), .ZN(new_n412));
  AOI22_X1  g226(.A1(new_n412), .A2(new_n392), .B1(new_n393), .B2(new_n402), .ZN(new_n413));
  OAI21_X1  g227(.A(G469), .B1(new_n413), .B2(G902), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(KEYINPUT9), .B(G234), .ZN(new_n416));
  OAI21_X1  g230(.A(G221), .B1(new_n416), .B2(G902), .ZN(new_n417));
  XOR2_X1   g231(.A(new_n417), .B(KEYINPUT79), .Z(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(G214), .B1(G237), .B2(G902), .ZN(new_n421));
  XOR2_X1   g235(.A(new_n421), .B(KEYINPUT82), .Z(new_n422));
  NAND2_X1  g236(.A1(new_n236), .A2(G125), .ZN(new_n423));
  AOI22_X1  g237(.A1(new_n232), .A2(new_n198), .B1(new_n191), .B2(new_n194), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n423), .B1(G125), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(G224), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n426), .A2(G953), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n425), .B(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT6), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n381), .A2(new_n240), .A3(new_n383), .ZN(new_n431));
  OR2_X1    g245(.A1(new_n238), .A2(new_n239), .ZN(new_n432));
  INV_X1    g246(.A(G116), .ZN(new_n433));
  NOR3_X1   g247(.A1(new_n433), .A2(KEYINPUT5), .A3(G119), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n434), .B(KEYINPUT83), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT5), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n435), .B(G113), .C1(new_n436), .C2(new_n238), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n372), .A2(new_n432), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n431), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT84), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  XOR2_X1   g255(.A(G110), .B(G122), .Z(new_n442));
  NAND3_X1  g256(.A1(new_n431), .A2(KEYINPUT84), .A3(new_n438), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  OR2_X1    g258(.A1(new_n439), .A2(new_n442), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n430), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AND3_X1   g260(.A1(new_n431), .A2(KEYINPUT84), .A3(new_n438), .ZN(new_n447));
  AOI21_X1  g261(.A(KEYINPUT84), .B1(new_n431), .B2(new_n438), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(KEYINPUT6), .B1(new_n449), .B2(new_n442), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n429), .B1(new_n446), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(G902), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n371), .A2(KEYINPUT85), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n437), .A2(new_n432), .ZN(new_n454));
  XOR2_X1   g268(.A(new_n453), .B(new_n454), .Z(new_n455));
  XOR2_X1   g269(.A(new_n442), .B(KEYINPUT8), .Z(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  AND2_X1   g271(.A1(new_n428), .A2(KEYINPUT7), .ZN(new_n458));
  OR2_X1    g272(.A1(new_n425), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n425), .A2(KEYINPUT7), .A3(new_n428), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n457), .A2(new_n459), .A3(new_n445), .A4(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n451), .A2(new_n452), .A3(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(G210), .B1(G237), .B2(G902), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n451), .A2(new_n452), .A3(new_n463), .A4(new_n461), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n422), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OR2_X1    g281(.A1(KEYINPUT93), .A2(G952), .ZN(new_n468));
  NAND2_X1  g282(.A1(KEYINPUT93), .A2(G952), .ZN(new_n469));
  AOI21_X1  g283(.A(G953), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(G234), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n470), .B1(new_n471), .B2(new_n248), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n257), .B(G953), .C1(new_n471), .C2(new_n248), .ZN(new_n473));
  XOR2_X1   g287(.A(KEYINPUT21), .B(G898), .Z(new_n474));
  OAI21_X1  g288(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n467), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n328), .A2(new_n329), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT87), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n248), .A2(new_n249), .A3(G214), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n188), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n248), .A2(new_n249), .A3(G143), .A4(G214), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n478), .B1(new_n482), .B2(G131), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n482), .A2(new_n478), .A3(G131), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(KEYINPUT17), .A3(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n485), .ZN(new_n487));
  OAI22_X1  g301(.A1(new_n487), .A2(new_n483), .B1(G131), .B2(new_n482), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n477), .B(new_n486), .C1(new_n488), .C2(KEYINPUT17), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n480), .A2(new_n481), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT86), .ZN(new_n491));
  AND2_X1   g305(.A1(KEYINPUT18), .A2(G131), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n490), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(KEYINPUT86), .B1(new_n482), .B2(new_n492), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n325), .A2(G146), .ZN(new_n496));
  AOI22_X1  g310(.A1(new_n494), .A2(new_n495), .B1(new_n338), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n482), .A2(new_n492), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  XOR2_X1   g313(.A(KEYINPUT89), .B(G104), .Z(new_n500));
  XNOR2_X1  g314(.A(G113), .B(G122), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n500), .B(new_n501), .ZN(new_n502));
  XOR2_X1   g316(.A(new_n502), .B(KEYINPUT90), .Z(new_n503));
  NAND3_X1  g317(.A1(new_n489), .A2(new_n499), .A3(new_n503), .ZN(new_n504));
  XOR2_X1   g318(.A(new_n325), .B(KEYINPUT19), .Z(new_n505));
  AOI21_X1  g319(.A(new_n329), .B1(new_n337), .B2(new_n505), .ZN(new_n506));
  AOI22_X1  g320(.A1(new_n506), .A2(new_n488), .B1(new_n497), .B2(new_n498), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT88), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n502), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n506), .A2(new_n488), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n510), .A2(new_n508), .A3(new_n499), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n504), .B1(new_n509), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(G475), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(new_n514), .A3(new_n452), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT20), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n504), .ZN(new_n518));
  INV_X1    g332(.A(new_n502), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n519), .B1(new_n489), .B2(new_n499), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n452), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(G475), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n513), .A2(KEYINPUT20), .A3(new_n514), .A4(new_n452), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n517), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(KEYINPUT91), .B(KEYINPUT13), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n525), .A2(G128), .A3(new_n188), .ZN(new_n526));
  XNOR2_X1  g340(.A(G128), .B(G143), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n526), .B(G134), .C1(new_n528), .C2(new_n525), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n212), .A2(new_n527), .ZN(new_n530));
  XNOR2_X1  g344(.A(G116), .B(G122), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n531), .A2(new_n365), .ZN(new_n532));
  INV_X1    g346(.A(new_n531), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n533), .A2(G107), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n529), .B(new_n530), .C1(new_n532), .C2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(KEYINPUT92), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n212), .B(new_n527), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n433), .A2(KEYINPUT14), .A3(G122), .ZN(new_n538));
  OAI211_X1 g352(.A(G107), .B(new_n538), .C1(new_n533), .C2(KEYINPUT14), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT92), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n540), .B1(new_n533), .B2(G107), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n536), .A2(new_n537), .A3(new_n539), .A4(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n535), .A2(new_n542), .ZN(new_n543));
  NOR3_X1   g357(.A1(new_n356), .A2(G953), .A3(new_n416), .ZN(new_n544));
  XOR2_X1   g358(.A(new_n543), .B(new_n544), .Z(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n352), .ZN(new_n546));
  INV_X1    g360(.A(G478), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n547), .A2(KEYINPUT15), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n546), .B(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n524), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NOR3_X1   g365(.A1(new_n420), .A2(new_n476), .A3(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n305), .A2(new_n359), .A3(new_n552), .ZN(new_n553));
  XNOR2_X1  g367(.A(KEYINPUT94), .B(G101), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n553), .B(new_n554), .ZN(G3));
  OAI21_X1  g369(.A(G472), .B1(new_n302), .B2(new_n257), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n296), .A2(new_n297), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n418), .B1(new_n411), .B2(new_n414), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n546), .A2(new_n547), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n561), .B(KEYINPUT96), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT95), .ZN(new_n563));
  OR3_X1    g377(.A1(new_n545), .A2(new_n563), .A3(KEYINPUT33), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT33), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(KEYINPUT95), .ZN(new_n566));
  OR2_X1    g380(.A1(new_n565), .A2(KEYINPUT95), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n545), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n569), .A2(G478), .A3(new_n352), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n562), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n524), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n476), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n559), .A2(new_n359), .A3(new_n560), .A4(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(G104), .ZN(new_n575));
  XNOR2_X1  g389(.A(KEYINPUT97), .B(KEYINPUT34), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n575), .B(new_n576), .ZN(G6));
  NAND4_X1  g391(.A1(new_n556), .A2(new_n359), .A3(new_n557), .A4(new_n560), .ZN(new_n578));
  INV_X1    g392(.A(new_n524), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n549), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n467), .A2(new_n475), .A3(new_n581), .ZN(new_n582));
  OR2_X1    g396(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  XOR2_X1   g397(.A(KEYINPUT35), .B(G107), .Z(new_n584));
  XNOR2_X1  g398(.A(new_n583), .B(new_n584), .ZN(G9));
  NAND2_X1  g399(.A1(new_n355), .A2(new_n357), .ZN(new_n586));
  OR2_X1    g400(.A1(new_n347), .A2(KEYINPUT36), .ZN(new_n587));
  XOR2_X1   g401(.A(new_n340), .B(new_n587), .Z(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n358), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n591), .A2(new_n558), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n552), .ZN(new_n593));
  XOR2_X1   g407(.A(KEYINPUT37), .B(G110), .Z(new_n594));
  XNOR2_X1  g408(.A(new_n593), .B(new_n594), .ZN(G12));
  NAND4_X1  g409(.A1(new_n305), .A2(new_n560), .A3(new_n467), .A4(new_n590), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n472), .B1(new_n473), .B2(G900), .ZN(new_n597));
  XOR2_X1   g411(.A(new_n597), .B(KEYINPUT98), .Z(new_n598));
  NOR2_X1   g412(.A1(new_n580), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(new_n197), .ZN(G30));
  NAND2_X1  g416(.A1(new_n524), .A2(new_n549), .ZN(new_n603));
  NOR3_X1   g417(.A1(new_n590), .A2(new_n422), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(KEYINPUT100), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n465), .A2(new_n466), .ZN(new_n606));
  XNOR2_X1  g420(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n296), .A2(new_n279), .A3(new_n297), .ZN(new_n609));
  OAI21_X1  g423(.A(KEYINPUT32), .B1(new_n302), .B2(new_n303), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n290), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n243), .A2(new_n244), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n612), .B1(new_n280), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(G472), .B1(new_n615), .B2(G902), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n611), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g431(.A(new_n598), .B(KEYINPUT39), .Z(new_n618));
  NAND2_X1  g432(.A1(new_n560), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(new_n619), .B(KEYINPUT40), .Z(new_n620));
  NAND4_X1  g434(.A1(new_n605), .A2(new_n608), .A3(new_n617), .A4(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(G143), .ZN(G45));
  NOR2_X1   g436(.A1(new_n572), .A2(new_n598), .ZN(new_n623));
  AND2_X1   g437(.A1(new_n560), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n305), .A2(new_n467), .A3(new_n590), .A4(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(KEYINPUT101), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n591), .B1(new_n611), .B2(new_n278), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT101), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n627), .A2(new_n628), .A3(new_n467), .A4(new_n624), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(G146), .ZN(G48));
  AOI22_X1  g445(.A1(new_n609), .A2(new_n610), .B1(G472), .B2(new_n277), .ZN(new_n632));
  INV_X1    g446(.A(new_n359), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n409), .A2(new_n352), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(G469), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n411), .A2(new_n419), .A3(new_n635), .ZN(new_n636));
  NOR3_X1   g450(.A1(new_n632), .A2(new_n633), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n637), .A2(KEYINPUT102), .A3(new_n573), .ZN(new_n638));
  INV_X1    g452(.A(new_n636), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n305), .A2(new_n359), .A3(new_n573), .A4(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT102), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(KEYINPUT41), .B(G113), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G15));
  INV_X1    g459(.A(new_n582), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n637), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT103), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n637), .A2(KEYINPUT103), .A3(new_n646), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G116), .ZN(G18));
  INV_X1    g466(.A(new_n467), .ZN(new_n653));
  NOR4_X1   g467(.A1(new_n632), .A2(new_n591), .A3(new_n653), .A4(new_n551), .ZN(new_n654));
  INV_X1    g468(.A(new_n475), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n636), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G119), .ZN(G21));
  INV_X1    g472(.A(new_n422), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT104), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n603), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n524), .A2(KEYINPUT104), .A3(new_n549), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n606), .A2(new_n659), .A3(new_n661), .A4(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(KEYINPUT105), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT105), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n467), .A2(new_n665), .A3(new_n661), .A4(new_n662), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n245), .A2(new_n247), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n299), .B1(new_n668), .B2(new_n254), .ZN(new_n669));
  INV_X1    g483(.A(new_n283), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n297), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n656), .A2(new_n556), .A3(new_n359), .A4(new_n671), .ZN(new_n672));
  OR2_X1    g486(.A1(new_n667), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G122), .ZN(G24));
  NAND4_X1  g488(.A1(new_n590), .A2(new_n556), .A3(new_n623), .A4(new_n671), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n639), .A2(new_n467), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(new_n323), .ZN(G27));
  NAND3_X1  g492(.A1(new_n609), .A2(new_n610), .A3(KEYINPUT106), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  AOI21_X1  g494(.A(KEYINPUT106), .B1(new_n609), .B2(new_n610), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n633), .B1(new_n682), .B2(new_n278), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n465), .A2(new_n659), .A3(new_n466), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n683), .A2(KEYINPUT42), .A3(new_n624), .A4(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n632), .A2(new_n633), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n420), .A2(new_n684), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n687), .A2(new_n623), .A3(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT42), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n686), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT107), .B(G131), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G33));
  NAND3_X1  g508(.A1(new_n687), .A2(new_n599), .A3(new_n688), .ZN(new_n695));
  XOR2_X1   g509(.A(KEYINPUT108), .B(G134), .Z(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G36));
  OAI21_X1  g511(.A(G469), .B1(new_n413), .B2(KEYINPUT45), .ZN(new_n698));
  OR2_X1    g512(.A1(new_n698), .A2(KEYINPUT109), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n413), .A2(KEYINPUT45), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n698), .A2(KEYINPUT109), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(G469), .A2(G902), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OR2_X1    g518(.A1(new_n704), .A2(KEYINPUT46), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n702), .A2(KEYINPUT46), .A3(new_n703), .ZN(new_n706));
  OR2_X1    g520(.A1(new_n706), .A2(KEYINPUT110), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(KEYINPUT110), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n705), .A2(new_n411), .A3(new_n707), .A4(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n709), .A2(new_n419), .A3(new_n618), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n571), .A2(new_n579), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(KEYINPUT43), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n558), .A2(new_n713), .A3(new_n590), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n685), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n714), .A2(new_n715), .ZN(new_n717));
  OR3_X1    g531(.A1(new_n710), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G137), .ZN(G39));
  NOR2_X1   g533(.A1(KEYINPUT111), .A2(KEYINPUT47), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n720), .B1(new_n709), .B2(new_n419), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n305), .A2(new_n359), .A3(new_n684), .ZN(new_n723));
  XOR2_X1   g537(.A(KEYINPUT111), .B(KEYINPUT47), .Z(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n709), .A2(new_n419), .A3(new_n725), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n722), .A2(new_n623), .A3(new_n723), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G140), .ZN(G42));
  INV_X1    g542(.A(KEYINPUT115), .ZN(new_n729));
  INV_X1    g543(.A(new_n695), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n730), .B1(new_n686), .B2(new_n691), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n574), .A2(new_n553), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n593), .B1(new_n732), .B2(KEYINPUT112), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n733), .B1(new_n649), .B2(new_n650), .ZN(new_n734));
  OAI22_X1  g548(.A1(new_n667), .A2(new_n672), .B1(new_n578), .B2(new_n582), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n735), .B1(new_n654), .B2(new_n656), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n732), .A2(KEYINPUT112), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n643), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n598), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n627), .A2(new_n550), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n675), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n688), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n731), .A2(new_n734), .A3(new_n738), .A4(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT114), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT52), .ZN(new_n745));
  OR2_X1    g559(.A1(new_n675), .A2(new_n676), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n746), .B1(new_n596), .B2(new_n600), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n747), .B1(new_n629), .B2(new_n626), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n420), .B1(new_n664), .B2(new_n666), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n617), .A2(new_n749), .A3(new_n591), .A4(new_n739), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT113), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AOI211_X1 g566(.A(new_n598), .B(new_n420), .C1(new_n664), .C2(new_n666), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n753), .A2(KEYINPUT113), .A3(new_n591), .A4(new_n617), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n745), .B1(new_n748), .B2(new_n755), .ZN(new_n756));
  NOR4_X1   g570(.A1(new_n632), .A2(new_n591), .A3(new_n420), .A4(new_n653), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n677), .B1(new_n757), .B2(new_n599), .ZN(new_n758));
  AND4_X1   g572(.A1(new_n745), .A2(new_n755), .A3(new_n758), .A4(new_n630), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n744), .B1(new_n756), .B2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n755), .A2(new_n630), .A3(new_n758), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(KEYINPUT52), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n755), .A2(new_n630), .A3(new_n758), .A4(new_n745), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(KEYINPUT114), .A3(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n743), .B1(new_n760), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n765), .A2(KEYINPUT53), .ZN(new_n766));
  AND4_X1   g580(.A1(new_n731), .A2(new_n734), .A3(new_n738), .A4(new_n742), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n756), .A2(new_n759), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n767), .A2(KEYINPUT53), .A3(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  OAI211_X1 g584(.A(new_n729), .B(KEYINPUT54), .C1(new_n766), .C2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(KEYINPUT116), .B(KEYINPUT51), .ZN(new_n772));
  INV_X1    g586(.A(new_n608), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT118), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n639), .A2(new_n774), .A3(new_n422), .ZN(new_n775));
  OAI21_X1  g589(.A(KEYINPUT118), .B1(new_n636), .B2(new_n659), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n773), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT119), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n556), .A2(new_n671), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n780), .A2(new_n359), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n712), .A2(new_n472), .ZN(new_n782));
  OR2_X1    g596(.A1(new_n777), .A2(new_n778), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n779), .A2(new_n781), .A3(new_n782), .A4(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT50), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n636), .A2(new_n684), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n780), .A2(new_n782), .A3(new_n590), .A4(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n617), .ZN(new_n789));
  INV_X1    g603(.A(new_n472), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n789), .A2(new_n359), .A3(new_n790), .A4(new_n787), .ZN(new_n791));
  OR3_X1    g605(.A1(new_n791), .A2(new_n524), .A3(new_n571), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n786), .A2(new_n788), .A3(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n781), .A2(new_n782), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n795), .A2(new_n684), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT117), .ZN(new_n797));
  INV_X1    g611(.A(new_n726), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n797), .B1(new_n798), .B2(new_n721), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n722), .A2(KEYINPUT117), .A3(new_n726), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n411), .A2(new_n635), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n802), .A2(new_n419), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n796), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n772), .B1(new_n794), .B2(new_n804), .ZN(new_n805));
  OAI221_X1 g619(.A(new_n470), .B1(new_n795), .B2(new_n676), .C1(new_n572), .C2(new_n791), .ZN(new_n806));
  XOR2_X1   g620(.A(new_n806), .B(KEYINPUT120), .Z(new_n807));
  AOI21_X1  g621(.A(new_n803), .B1(new_n722), .B2(new_n726), .ZN(new_n808));
  INV_X1    g622(.A(new_n796), .ZN(new_n809));
  OAI21_X1  g623(.A(KEYINPUT51), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n807), .B1(new_n793), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n683), .A2(new_n782), .A3(new_n787), .ZN(new_n812));
  XOR2_X1   g626(.A(new_n812), .B(KEYINPUT48), .Z(new_n813));
  NOR3_X1   g627(.A1(new_n805), .A2(new_n811), .A3(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n767), .A2(new_n815), .A3(new_n768), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n816), .B1(new_n765), .B2(new_n815), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT54), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT115), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n762), .A2(KEYINPUT114), .A3(new_n763), .ZN(new_n820));
  AOI21_X1  g634(.A(KEYINPUT114), .B1(new_n762), .B2(new_n763), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n767), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(new_n815), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n818), .B1(new_n823), .B2(new_n769), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n771), .B(new_n814), .C1(new_n819), .C2(new_n824), .ZN(new_n825));
  OR2_X1    g639(.A1(G952), .A2(G953), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n359), .B1(KEYINPUT49), .B2(new_n802), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n828), .B1(KEYINPUT49), .B2(new_n802), .ZN(new_n829));
  NOR4_X1   g643(.A1(new_n608), .A2(new_n418), .A3(new_n422), .A4(new_n711), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n829), .A2(new_n789), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n827), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT121), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n827), .A2(KEYINPUT121), .A3(new_n831), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(G75));
  OR2_X1    g650(.A1(new_n446), .A2(new_n450), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(new_n429), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n838), .B(KEYINPUT122), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n839), .B(KEYINPUT55), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT56), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n822), .A2(KEYINPUT53), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n842), .A2(new_n257), .A3(new_n816), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n841), .B1(new_n843), .B2(new_n463), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT123), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT123), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n846), .B(new_n841), .C1(new_n843), .C2(new_n463), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n840), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n249), .A2(G952), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n847), .A2(new_n840), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(G51));
  XNOR2_X1  g665(.A(new_n817), .B(KEYINPUT54), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n703), .B(KEYINPUT57), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n409), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  OR2_X1    g668(.A1(new_n843), .A2(new_n702), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n849), .B1(new_n854), .B2(new_n855), .ZN(G54));
  INV_X1    g670(.A(new_n817), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n857), .A2(KEYINPUT58), .A3(G475), .A4(new_n257), .ZN(new_n858));
  XOR2_X1   g672(.A(new_n858), .B(new_n513), .Z(new_n859));
  NOR2_X1   g673(.A1(new_n859), .A2(new_n849), .ZN(G60));
  NAND2_X1  g674(.A1(G478), .A2(G902), .ZN(new_n861));
  XOR2_X1   g675(.A(new_n861), .B(KEYINPUT59), .Z(new_n862));
  AOI211_X1 g676(.A(new_n862), .B(new_n852), .C1(new_n564), .C2(new_n568), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n771), .B1(new_n819), .B2(new_n824), .ZN(new_n864));
  INV_X1    g678(.A(new_n862), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n569), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n863), .A2(new_n866), .A3(new_n849), .ZN(G63));
  INV_X1    g681(.A(KEYINPUT124), .ZN(new_n868));
  NAND2_X1  g682(.A1(G217), .A2(G902), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(KEYINPUT60), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n842), .A2(new_n816), .A3(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(new_n588), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n868), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n857), .A2(KEYINPUT124), .A3(new_n588), .A4(new_n871), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n849), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n872), .A2(new_n350), .A3(new_n349), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT61), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n879), .B(new_n880), .ZN(G66));
  INV_X1    g695(.A(new_n474), .ZN(new_n882));
  OAI21_X1  g696(.A(G953), .B1(new_n882), .B2(new_n426), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n738), .A2(new_n734), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n883), .B1(new_n885), .B2(G953), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT125), .ZN(new_n887));
  INV_X1    g701(.A(G898), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n837), .B1(new_n888), .B2(G953), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n887), .B(new_n889), .ZN(G69));
  AND2_X1   g704(.A1(new_n270), .A2(new_n272), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n891), .B(new_n505), .Z(new_n892));
  OAI21_X1  g706(.A(G900), .B1(new_n892), .B2(new_n389), .ZN(new_n893));
  AOI211_X1 g707(.A(new_n249), .B(new_n893), .C1(new_n389), .C2(new_n892), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n718), .A2(new_n748), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT126), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n710), .A2(new_n667), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(new_n683), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n898), .A2(new_n731), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n896), .A2(new_n727), .A3(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(new_n892), .ZN(new_n901));
  AOI21_X1  g715(.A(G953), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n748), .A2(new_n621), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n903), .B(KEYINPUT62), .Z(new_n904));
  AOI211_X1 g718(.A(new_n684), .B(new_n619), .C1(new_n572), .C2(new_n580), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(new_n687), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n904), .A2(new_n718), .A3(new_n727), .A4(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n892), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n894), .B1(new_n902), .B2(new_n908), .ZN(G72));
  NAND2_X1  g723(.A1(new_n273), .A2(new_n242), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n896), .A2(new_n727), .A3(new_n885), .A4(new_n899), .ZN(new_n911));
  NAND2_X1  g725(.A1(G472), .A2(G902), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(KEYINPUT63), .Z(new_n913));
  AOI21_X1  g727(.A(new_n910), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n849), .B1(new_n914), .B2(new_n280), .ZN(new_n915));
  OAI221_X1 g729(.A(new_n913), .B1(new_n612), .B2(new_n274), .C1(new_n766), .C2(new_n770), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n913), .B1(new_n907), .B2(new_n884), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n917), .A2(new_n254), .A3(new_n910), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n915), .A2(new_n916), .A3(new_n918), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT127), .ZN(G57));
endmodule


