//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 1 0 0 0 1 0 0 1 1 1 1 0 0 1 0 0 1 0 0 0 1 0 0 1 0 1 0 0 1 1 1 0 0 0 1 1 0 1 0 1 0 1 0 1 0 1 0 1 0 1 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:13 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n762, new_n763, new_n764,
    new_n765, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1002, new_n1003, new_n1004, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(G113), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(KEYINPUT2), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT2), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G113), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(G116), .B(G119), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n192), .B(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT1), .ZN(new_n196));
  INV_X1    g010(.A(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G143), .ZN(new_n198));
  INV_X1    g012(.A(G143), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G146), .ZN(new_n200));
  AND4_X1   g014(.A1(new_n196), .A2(new_n198), .A3(new_n200), .A4(G128), .ZN(new_n201));
  OAI21_X1  g015(.A(KEYINPUT1), .B1(new_n199), .B2(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT68), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT68), .ZN(new_n204));
  OAI211_X1 g018(.A(new_n204), .B(KEYINPUT1), .C1(new_n199), .C2(G146), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n203), .A2(G128), .A3(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(G143), .B(G146), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n201), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G137), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G134), .ZN(new_n211));
  INV_X1    g025(.A(G134), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G137), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G131), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT11), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n216), .B1(new_n212), .B2(G137), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n210), .A2(KEYINPUT11), .A3(G134), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n218), .A3(new_n213), .ZN(new_n219));
  XNOR2_X1  g033(.A(KEYINPUT66), .B(G131), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n215), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n209), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT72), .ZN(new_n223));
  NAND2_X1  g037(.A1(KEYINPUT0), .A2(G128), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n198), .A2(new_n200), .A3(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT71), .ZN(new_n226));
  INV_X1    g040(.A(new_n224), .ZN(new_n227));
  NOR2_X1   g041(.A1(KEYINPUT0), .A2(G128), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n225), .B(new_n226), .C1(new_n229), .C2(new_n207), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n199), .A2(G146), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n197), .A2(G143), .ZN(new_n233));
  OAI22_X1  g047(.A1(new_n232), .A2(new_n233), .B1(new_n227), .B2(new_n228), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n226), .B1(new_n234), .B2(new_n225), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n231), .A2(new_n235), .ZN(new_n236));
  AND2_X1   g050(.A1(new_n219), .A2(KEYINPUT67), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n217), .A2(new_n218), .A3(new_n238), .A4(new_n213), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G131), .ZN(new_n240));
  OAI22_X1  g054(.A1(new_n237), .A2(new_n240), .B1(new_n220), .B2(new_n219), .ZN(new_n241));
  AOI22_X1  g055(.A1(new_n222), .A2(new_n223), .B1(new_n236), .B2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(KEYINPUT72), .B1(new_n209), .B2(new_n221), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n195), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n236), .A2(new_n241), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n205), .A2(G128), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n204), .B1(new_n198), .B2(KEYINPUT1), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n208), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n201), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  AND3_X1   g064(.A1(new_n217), .A2(new_n218), .A3(new_n213), .ZN(new_n251));
  XOR2_X1   g065(.A(KEYINPUT66), .B(G131), .Z(new_n252));
  AOI22_X1  g066(.A1(new_n251), .A2(new_n252), .B1(G131), .B2(new_n214), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n250), .A2(new_n223), .A3(new_n253), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n245), .A2(new_n195), .A3(new_n243), .A4(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  OAI21_X1  g070(.A(KEYINPUT28), .B1(new_n244), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT75), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n245), .A2(new_n243), .A3(new_n254), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(new_n194), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(new_n255), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n262), .A2(KEYINPUT75), .A3(KEYINPUT28), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT28), .ZN(new_n265));
  AND2_X1   g079(.A1(new_n239), .A2(G131), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n219), .A2(KEYINPUT67), .ZN(new_n267));
  AOI22_X1  g081(.A1(new_n266), .A2(new_n267), .B1(new_n252), .B2(new_n251), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n225), .B1(new_n229), .B2(new_n207), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT71), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(new_n230), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n195), .B1(new_n209), .B2(new_n221), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n265), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NOR2_X1   g088(.A1(G237), .A2(G953), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G210), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n276), .B(KEYINPUT27), .ZN(new_n277));
  XNOR2_X1  g091(.A(KEYINPUT26), .B(G101), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n277), .B(new_n278), .ZN(new_n279));
  AND3_X1   g093(.A1(new_n274), .A2(KEYINPUT29), .A3(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(G902), .B1(new_n264), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n274), .A2(new_n279), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT69), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n283), .B1(new_n209), .B2(new_n221), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n250), .A2(KEYINPUT69), .A3(new_n253), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n225), .B(KEYINPUT65), .C1(new_n229), .C2(new_n207), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT65), .B1(new_n234), .B2(new_n225), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI22_X1  g103(.A1(new_n284), .A2(new_n285), .B1(new_n241), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n255), .B1(new_n290), .B2(new_n195), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n282), .B1(new_n291), .B2(KEYINPUT28), .ZN(new_n292));
  AOI21_X1  g106(.A(KEYINPUT29), .B1(new_n292), .B2(KEYINPUT74), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT74), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n291), .A2(KEYINPUT28), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n294), .B1(new_n295), .B2(new_n282), .ZN(new_n296));
  INV_X1    g110(.A(new_n279), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n245), .A2(KEYINPUT30), .A3(new_n243), .A4(new_n254), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(new_n194), .ZN(new_n299));
  XOR2_X1   g113(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n300));
  OAI21_X1  g114(.A(KEYINPUT70), .B1(new_n290), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n289), .A2(new_n241), .ZN(new_n302));
  NOR3_X1   g116(.A1(new_n209), .A2(new_n283), .A3(new_n221), .ZN(new_n303));
  AOI21_X1  g117(.A(KEYINPUT69), .B1(new_n250), .B2(new_n253), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT70), .ZN(new_n306));
  INV_X1    g120(.A(new_n300), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n299), .B1(new_n301), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n297), .B1(new_n309), .B2(new_n256), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n293), .A2(new_n296), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n187), .B1(new_n281), .B2(new_n311), .ZN(new_n312));
  NOR2_X1   g126(.A1(G472), .A2(G902), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT32), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n299), .ZN(new_n318));
  NOR3_X1   g132(.A1(new_n290), .A2(KEYINPUT70), .A3(new_n300), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n306), .B1(new_n305), .B2(new_n307), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT73), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n255), .A2(new_n279), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n321), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT73), .B1(new_n309), .B2(new_n323), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n325), .A2(new_n326), .A3(KEYINPUT31), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n291), .A2(KEYINPUT28), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n279), .B1(new_n328), .B2(new_n274), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT31), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n301), .A2(new_n308), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n323), .B1(new_n331), .B2(new_n318), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n329), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n317), .B1(new_n327), .B2(new_n333), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n312), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n327), .A2(new_n333), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n313), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n315), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(G214), .B1(G237), .B2(G902), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G104), .ZN(new_n342));
  OAI21_X1  g156(.A(KEYINPUT3), .B1(new_n342), .B2(G107), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT3), .ZN(new_n344));
  INV_X1    g158(.A(G107), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n344), .A2(new_n345), .A3(G104), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n342), .A2(G107), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n343), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(G101), .ZN(new_n349));
  INV_X1    g163(.A(G101), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n343), .A2(new_n346), .A3(new_n350), .A4(new_n347), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n349), .A2(KEYINPUT4), .A3(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT4), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n348), .A2(new_n353), .A3(G101), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n352), .A2(new_n194), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n192), .A2(new_n193), .ZN(new_n356));
  INV_X1    g170(.A(G119), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G116), .ZN(new_n358));
  INV_X1    g172(.A(G116), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G119), .ZN(new_n360));
  AND3_X1   g174(.A1(new_n358), .A2(new_n360), .A3(KEYINPUT5), .ZN(new_n361));
  OAI21_X1  g175(.A(G113), .B1(new_n358), .B2(KEYINPUT5), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n356), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT79), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n364), .A2(new_n345), .A3(G104), .ZN(new_n365));
  OAI21_X1  g179(.A(KEYINPUT79), .B1(new_n342), .B2(G107), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n345), .A2(G104), .ZN(new_n367));
  OAI211_X1 g181(.A(G101), .B(new_n365), .C1(new_n366), .C2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n351), .ZN(new_n369));
  OR2_X1    g183(.A1(new_n363), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n355), .A2(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(G110), .B(G122), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n355), .A2(new_n370), .A3(new_n372), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n374), .A2(KEYINPUT6), .A3(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT6), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n371), .A2(new_n377), .A3(new_n373), .ZN(new_n378));
  INV_X1    g192(.A(G125), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n248), .A2(new_n249), .A3(new_n379), .ZN(new_n380));
  OAI211_X1 g194(.A(new_n225), .B(G125), .C1(new_n229), .C2(new_n207), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G224), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n383), .A2(G953), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n382), .B(new_n384), .ZN(new_n385));
  AND3_X1   g199(.A1(new_n376), .A2(new_n378), .A3(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(G902), .ZN(new_n387));
  OAI21_X1  g201(.A(KEYINPUT7), .B1(new_n383), .B2(G953), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  AND2_X1   g203(.A1(new_n381), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n380), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT84), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n390), .A2(new_n380), .A3(KEYINPUT84), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n389), .B1(new_n380), .B2(new_n381), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(KEYINPUT83), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n372), .B(KEYINPUT8), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n363), .A2(new_n369), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n358), .A2(new_n360), .A3(KEYINPUT5), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n401), .B(G113), .C1(KEYINPUT5), .C2(new_n358), .ZN(new_n402));
  AOI22_X1  g216(.A1(new_n402), .A2(new_n356), .B1(new_n351), .B2(new_n368), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n399), .B1(new_n400), .B2(new_n403), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n375), .B(new_n404), .C1(KEYINPUT83), .C2(new_n396), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n387), .B1(new_n398), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(KEYINPUT85), .B1(new_n386), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n375), .A2(new_n404), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n396), .A2(KEYINPUT83), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI22_X1  g224(.A1(new_n393), .A2(new_n394), .B1(KEYINPUT83), .B2(new_n396), .ZN(new_n411));
  AOI21_X1  g225(.A(G902), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT85), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n376), .A2(new_n378), .A3(new_n385), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(G210), .B1(G237), .B2(G902), .ZN(new_n416));
  XOR2_X1   g230(.A(new_n416), .B(KEYINPUT86), .Z(new_n417));
  NAND3_X1  g231(.A1(new_n407), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n412), .A2(new_n414), .A3(new_n416), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n341), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(G140), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(G125), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n379), .A2(G140), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n422), .A2(new_n423), .A3(KEYINPUT16), .ZN(new_n424));
  OR3_X1    g238(.A1(new_n379), .A2(KEYINPUT16), .A3(G140), .ZN(new_n425));
  AND3_X1   g239(.A1(new_n424), .A2(G146), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(G146), .B1(new_n424), .B2(new_n425), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n275), .A2(G143), .A3(G214), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(G143), .B1(new_n275), .B2(G214), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n220), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT17), .ZN(new_n433));
  INV_X1    g247(.A(G237), .ZN(new_n434));
  INV_X1    g248(.A(G953), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n434), .A2(new_n435), .A3(G214), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n199), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n252), .A2(new_n437), .A3(new_n429), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n432), .A2(new_n433), .A3(new_n438), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n428), .B(new_n439), .C1(new_n433), .C2(new_n432), .ZN(new_n440));
  OAI211_X1 g254(.A(KEYINPUT18), .B(G131), .C1(new_n430), .C2(new_n431), .ZN(new_n441));
  NAND2_X1  g255(.A1(KEYINPUT18), .A2(G131), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n437), .A2(new_n429), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n422), .A2(new_n423), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(G146), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n422), .A2(new_n423), .A3(new_n197), .ZN(new_n446));
  AND3_X1   g260(.A1(new_n445), .A2(new_n446), .A3(KEYINPUT87), .ZN(new_n447));
  AOI21_X1  g261(.A(KEYINPUT87), .B1(new_n445), .B2(new_n446), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n441), .B(new_n443), .C1(new_n447), .C2(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(G113), .B(G122), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n450), .B(new_n342), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n440), .A2(new_n449), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n451), .B1(new_n440), .B2(new_n449), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n387), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(G475), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT20), .ZN(new_n456));
  AND3_X1   g270(.A1(new_n422), .A2(new_n423), .A3(KEYINPUT19), .ZN(new_n457));
  AOI21_X1  g271(.A(KEYINPUT19), .B1(new_n422), .B2(new_n423), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(KEYINPUT88), .B1(new_n459), .B2(G146), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n424), .A2(new_n425), .A3(G146), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n432), .A2(new_n438), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT88), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n463), .B(new_n197), .C1(new_n457), .C2(new_n458), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n460), .A2(new_n461), .A3(new_n462), .A4(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n449), .ZN(new_n466));
  INV_X1    g280(.A(new_n451), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n440), .A2(new_n449), .A3(new_n451), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g284(.A1(G475), .A2(G902), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n456), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n451), .B1(new_n465), .B2(new_n449), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n456), .B(new_n471), .C1(new_n452), .C2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n455), .B1(new_n472), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n435), .A2(G952), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n477), .B1(G234), .B2(G237), .ZN(new_n478));
  XNOR2_X1  g292(.A(KEYINPUT21), .B(G898), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n479), .B(KEYINPUT96), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  AOI211_X1 g295(.A(new_n387), .B(new_n435), .C1(G234), .C2(G237), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n478), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n476), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(G128), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(G143), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n199), .A2(G128), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n486), .A2(new_n487), .A3(new_n212), .ZN(new_n488));
  XOR2_X1   g302(.A(new_n488), .B(KEYINPUT91), .Z(new_n489));
  INV_X1    g303(.A(KEYINPUT90), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n199), .A2(G128), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT13), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n490), .B(new_n487), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n485), .A2(G143), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n494), .B1(KEYINPUT13), .B2(new_n486), .ZN(new_n495));
  OAI21_X1  g309(.A(KEYINPUT90), .B1(new_n487), .B2(new_n492), .ZN(new_n496));
  OAI211_X1 g310(.A(G134), .B(new_n493), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT89), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n498), .B1(new_n359), .B2(G122), .ZN(new_n499));
  INV_X1    g313(.A(G122), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n500), .A2(KEYINPUT89), .A3(G116), .ZN(new_n501));
  AOI22_X1  g315(.A1(new_n499), .A2(new_n501), .B1(new_n359), .B2(G122), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n502), .A2(new_n345), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n502), .A2(new_n345), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n489), .B(new_n497), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n499), .A2(new_n501), .ZN(new_n506));
  OR3_X1    g320(.A1(new_n500), .A2(KEYINPUT14), .A3(G116), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(KEYINPUT14), .B1(new_n500), .B2(G116), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(KEYINPUT92), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT92), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n511), .B(KEYINPUT14), .C1(new_n500), .C2(G116), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(G107), .B1(new_n508), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(G134), .B1(new_n491), .B2(new_n494), .ZN(new_n515));
  AOI22_X1  g329(.A1(new_n345), .A2(new_n502), .B1(new_n515), .B2(new_n488), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT93), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n514), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n517), .B1(new_n514), .B2(new_n516), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n505), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  XNOR2_X1  g334(.A(KEYINPUT9), .B(G234), .ZN(new_n521));
  INV_X1    g335(.A(G217), .ZN(new_n522));
  NOR3_X1   g336(.A1(new_n521), .A2(new_n522), .A3(G953), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n505), .B(new_n523), .C1(new_n518), .C2(new_n519), .ZN(new_n526));
  AOI21_X1  g340(.A(G902), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT94), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI211_X1 g343(.A(KEYINPUT94), .B(G902), .C1(new_n525), .C2(new_n526), .ZN(new_n530));
  INV_X1    g344(.A(G478), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n531), .A2(KEYINPUT15), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NOR3_X1   g347(.A1(new_n529), .A2(new_n530), .A3(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT95), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n525), .A2(new_n526), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n387), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n537), .A2(new_n532), .ZN(new_n538));
  NOR3_X1   g352(.A1(new_n534), .A2(new_n535), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n537), .A2(KEYINPUT94), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n527), .A2(new_n528), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n540), .A2(new_n532), .A3(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n538), .ZN(new_n543));
  AOI21_X1  g357(.A(KEYINPUT95), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n420), .B(new_n484), .C1(new_n539), .C2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT78), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT23), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n548), .B1(new_n357), .B2(G128), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n357), .A2(G128), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n485), .A2(KEYINPUT23), .A3(G119), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(G119), .B(G128), .ZN(new_n553));
  INV_X1    g367(.A(G110), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(KEYINPUT24), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT24), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(G110), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  OAI22_X1  g372(.A1(new_n552), .A2(G110), .B1(new_n553), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n559), .A2(new_n461), .A3(new_n446), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n424), .A2(new_n425), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(new_n197), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n461), .ZN(new_n563));
  AOI22_X1  g377(.A1(new_n552), .A2(G110), .B1(new_n553), .B2(new_n558), .ZN(new_n564));
  AOI21_X1  g378(.A(KEYINPUT76), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n564), .B(KEYINPUT76), .C1(new_n426), .C2(new_n427), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n560), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(KEYINPUT22), .B(G137), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n435), .A2(G221), .A3(G234), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n569), .B(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n560), .B(new_n571), .C1(new_n565), .C2(new_n567), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n573), .A2(new_n387), .A3(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT25), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n573), .A2(KEYINPUT25), .A3(new_n387), .A4(new_n574), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n577), .A2(KEYINPUT77), .A3(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT77), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n575), .A2(new_n580), .A3(new_n576), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n522), .B1(G234), .B2(new_n387), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n547), .B1(new_n579), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n577), .A2(KEYINPUT77), .A3(new_n578), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n585), .A2(KEYINPUT78), .A3(new_n582), .A4(new_n581), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n582), .A2(G902), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n573), .A2(new_n574), .A3(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n584), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(G221), .B1(new_n521), .B2(G902), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n248), .A2(new_n369), .A3(new_n249), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n207), .B1(G128), .B2(new_n202), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n351), .B(new_n368), .C1(new_n594), .C2(new_n201), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n596), .A2(KEYINPUT12), .A3(new_n241), .ZN(new_n597));
  AOI21_X1  g411(.A(KEYINPUT12), .B1(new_n596), .B2(new_n241), .ZN(new_n598));
  OAI21_X1  g412(.A(KEYINPUT81), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n596), .A2(new_n241), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT12), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT81), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n596), .A2(KEYINPUT12), .A3(new_n241), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT10), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n595), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n352), .A2(new_n270), .A3(new_n230), .A4(new_n354), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n369), .A2(new_n606), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n250), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n607), .A2(new_n608), .A3(new_n610), .A4(new_n268), .ZN(new_n611));
  XNOR2_X1  g425(.A(G110), .B(G140), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n435), .A2(G227), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  AND2_X1   g429(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n599), .A2(new_n605), .A3(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT82), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n599), .A2(new_n605), .A3(new_n616), .A4(KEYINPUT82), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n608), .A2(new_n607), .A3(new_n610), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n241), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n611), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n614), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(KEYINPUT80), .B(G469), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n626), .A2(new_n387), .A3(new_n628), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n611), .B1(new_n597), .B2(new_n598), .ZN(new_n630));
  AOI22_X1  g444(.A1(new_n630), .A2(new_n614), .B1(new_n616), .B2(new_n623), .ZN(new_n631));
  OAI21_X1  g445(.A(G469), .B1(new_n631), .B2(G902), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n592), .B1(new_n629), .B2(new_n632), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n339), .A2(new_n546), .A3(new_n590), .A4(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(G101), .ZN(G3));
  NAND2_X1  g449(.A1(new_n336), .A2(new_n387), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(G472), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n337), .ZN(new_n638));
  AOI22_X1  g452(.A1(new_n619), .A2(new_n620), .B1(new_n614), .B2(new_n624), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n639), .A2(G902), .A3(new_n627), .ZN(new_n640));
  INV_X1    g454(.A(new_n632), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n591), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n470), .A2(new_n471), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(KEYINPUT20), .ZN(new_n645));
  AOI22_X1  g459(.A1(new_n645), .A2(new_n474), .B1(G475), .B2(new_n454), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n540), .A2(new_n531), .A3(new_n541), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n531), .A2(G902), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n536), .A2(KEYINPUT97), .A3(KEYINPUT33), .ZN(new_n649));
  NOR2_X1   g463(.A1(KEYINPUT97), .A2(KEYINPUT33), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT97), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT33), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AOI211_X1 g467(.A(new_n650), .B(new_n653), .C1(new_n525), .C2(new_n526), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n648), .B1(new_n649), .B2(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n646), .B1(new_n647), .B2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n416), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n657), .B1(new_n386), .B2(new_n406), .ZN(new_n658));
  AOI211_X1 g472(.A(new_n341), .B(new_n483), .C1(new_n658), .C2(new_n419), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n660), .A2(new_n589), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n643), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(new_n342), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT98), .B(KEYINPUT34), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G6));
  OAI21_X1  g479(.A(new_n535), .B1(new_n534), .B2(new_n538), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n542), .A2(new_n543), .A3(KEYINPUT95), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n666), .A2(new_n659), .A3(new_n667), .A4(new_n646), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n668), .A2(new_n589), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n643), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT35), .B(G107), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G9));
  AOI21_X1  g486(.A(new_n314), .B1(new_n327), .B2(new_n333), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n673), .B1(new_n636), .B2(G472), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n572), .A2(KEYINPUT36), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT99), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(new_n568), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n587), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n584), .A2(new_n586), .A3(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n546), .A2(new_n674), .A3(new_n633), .A4(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT37), .B(G110), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G12));
  AOI21_X1  g496(.A(new_n341), .B1(new_n658), .B2(new_n419), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n684), .A2(new_n642), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n666), .A2(new_n667), .ZN(new_n686));
  INV_X1    g500(.A(G900), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n482), .A2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n478), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n646), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n686), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n685), .A2(new_n339), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G128), .ZN(G30));
  XNOR2_X1  g508(.A(new_n690), .B(KEYINPUT39), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n642), .A2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  OR2_X1    g512(.A1(new_n698), .A2(KEYINPUT40), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(KEYINPUT40), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n418), .A2(new_n419), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT38), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n686), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n704), .A2(new_n340), .A3(new_n476), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n703), .A2(new_n705), .A3(new_n679), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n262), .A2(new_n297), .ZN(new_n707));
  AND3_X1   g521(.A1(new_n325), .A2(new_n326), .A3(new_n707), .ZN(new_n708));
  OAI21_X1  g522(.A(G472), .B1(new_n708), .B2(G902), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n336), .A2(new_n316), .ZN(new_n710));
  OAI211_X1 g524(.A(new_n709), .B(new_n710), .C1(KEYINPUT32), .C2(new_n673), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n699), .A2(new_n700), .A3(new_n706), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G143), .ZN(G45));
  NAND2_X1  g527(.A1(new_n656), .A2(new_n690), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n293), .A2(new_n296), .A3(new_n310), .ZN(new_n716));
  AOI21_X1  g530(.A(KEYINPUT75), .B1(new_n262), .B2(KEYINPUT28), .ZN(new_n717));
  AOI211_X1 g531(.A(new_n258), .B(new_n265), .C1(new_n261), .C2(new_n255), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n280), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n387), .ZN(new_n720));
  OAI21_X1  g534(.A(G472), .B1(new_n716), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n710), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n673), .A2(KEYINPUT32), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n715), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n633), .A2(new_n683), .A3(new_n679), .ZN(new_n725));
  OAI21_X1  g539(.A(KEYINPUT100), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n714), .B1(new_n335), .B2(new_n338), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT100), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n727), .A2(new_n728), .A3(new_n685), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G146), .ZN(G48));
  OAI21_X1  g545(.A(G469), .B1(new_n639), .B2(G902), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n629), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n733), .A2(new_n592), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n339), .A2(new_n734), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n735), .A2(new_n589), .A3(new_n660), .ZN(new_n736));
  XOR2_X1   g550(.A(KEYINPUT41), .B(G113), .Z(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(G15));
  NAND3_X1  g552(.A1(new_n339), .A2(new_n669), .A3(new_n734), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G116), .ZN(G18));
  NAND4_X1  g554(.A1(new_n629), .A2(new_n732), .A3(new_n591), .A4(new_n683), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n484), .B1(new_n539), .B2(new_n544), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n339), .A2(new_n742), .A3(new_n744), .A4(new_n679), .ZN(new_n745));
  XOR2_X1   g559(.A(KEYINPUT101), .B(G119), .Z(new_n746));
  XNOR2_X1  g560(.A(new_n745), .B(new_n746), .ZN(G21));
  OAI21_X1  g561(.A(new_n274), .B1(new_n717), .B2(new_n718), .ZN(new_n748));
  AOI22_X1  g562(.A1(new_n748), .A2(new_n297), .B1(new_n330), .B2(new_n332), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n327), .ZN(new_n750));
  XOR2_X1   g564(.A(new_n313), .B(KEYINPUT102), .Z(new_n751));
  AOI22_X1  g565(.A1(new_n636), .A2(G472), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  AND2_X1   g566(.A1(new_n375), .A2(new_n404), .ZN(new_n753));
  INV_X1    g567(.A(new_n409), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n411), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  AND4_X1   g569(.A1(new_n387), .A2(new_n414), .A3(new_n755), .A4(new_n416), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n416), .B1(new_n412), .B2(new_n414), .ZN(new_n757));
  OAI211_X1 g571(.A(new_n476), .B(new_n340), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  NOR4_X1   g572(.A1(new_n539), .A2(new_n544), .A3(new_n758), .A4(new_n483), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n752), .A2(new_n759), .A3(new_n734), .A4(new_n590), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G122), .ZN(G24));
  NAND2_X1  g575(.A1(new_n750), .A2(new_n751), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n637), .A2(new_n679), .A3(new_n762), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n741), .A2(new_n714), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G125), .ZN(G27));
  OAI21_X1  g580(.A(KEYINPUT104), .B1(new_n701), .B2(new_n341), .ZN(new_n767));
  INV_X1    g581(.A(G469), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n630), .A2(new_n614), .ZN(new_n769));
  INV_X1    g583(.A(new_n623), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n611), .A2(new_n615), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT103), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(KEYINPUT103), .B1(new_n616), .B2(new_n623), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n769), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n768), .B1(new_n775), .B2(new_n387), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n629), .A2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT104), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n418), .A2(new_n779), .A3(new_n340), .A4(new_n419), .ZN(new_n780));
  AND4_X1   g594(.A1(new_n591), .A2(new_n767), .A3(new_n778), .A4(new_n780), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n781), .A2(new_n339), .A3(new_n590), .A4(new_n715), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT42), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n767), .A2(new_n591), .A3(new_n780), .ZN(new_n785));
  AOI21_X1  g599(.A(G902), .B1(new_n621), .B2(new_n625), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n776), .B1(new_n786), .B2(new_n628), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n785), .A2(new_n714), .A3(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n723), .A2(new_n312), .ZN(new_n789));
  OR2_X1    g603(.A1(new_n334), .A2(KEYINPUT105), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n334), .A2(KEYINPUT105), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n789), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n788), .A2(new_n792), .A3(KEYINPUT42), .A4(new_n590), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n784), .A2(new_n793), .ZN(new_n794));
  XOR2_X1   g608(.A(KEYINPUT106), .B(G131), .Z(new_n795));
  XNOR2_X1  g609(.A(new_n794), .B(new_n795), .ZN(G33));
  NAND4_X1  g610(.A1(new_n781), .A2(new_n339), .A3(new_n590), .A4(new_n692), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G134), .ZN(G36));
  INV_X1    g612(.A(KEYINPUT107), .ZN(new_n799));
  NAND2_X1  g613(.A1(G469), .A2(G902), .ZN(new_n800));
  OAI211_X1 g614(.A(KEYINPUT45), .B(new_n769), .C1(new_n773), .C2(new_n774), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g616(.A(G469), .B1(new_n631), .B2(KEYINPUT45), .ZN(new_n803));
  OAI211_X1 g617(.A(KEYINPUT46), .B(new_n800), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n799), .B1(new_n804), .B2(new_n629), .ZN(new_n805));
  OR2_X1    g619(.A1(new_n802), .A2(new_n803), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT46), .B1(new_n806), .B2(new_n800), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n804), .A2(new_n799), .A3(new_n629), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n810), .A2(new_n591), .A3(new_n695), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n767), .A2(new_n780), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n638), .A2(new_n679), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(KEYINPUT109), .ZN(new_n815));
  AOI21_X1  g629(.A(KEYINPUT43), .B1(new_n646), .B2(KEYINPUT108), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n647), .A2(new_n655), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n816), .B1(new_n818), .B2(new_n476), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n817), .B(new_n646), .C1(KEYINPUT108), .C2(KEYINPUT43), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT109), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n638), .A2(new_n822), .A3(new_n679), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n815), .A2(new_n821), .A3(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT44), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n813), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT110), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n827), .B1(new_n824), .B2(new_n825), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n824), .A2(new_n827), .A3(new_n825), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(G137), .ZN(G39));
  XNOR2_X1  g646(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n809), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n835), .A2(new_n805), .A3(new_n807), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n834), .B1(new_n836), .B2(new_n592), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n810), .A2(new_n591), .A3(new_n833), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NOR4_X1   g653(.A1(new_n339), .A2(new_n812), .A3(new_n590), .A4(new_n714), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(G140), .ZN(G42));
  NAND4_X1  g656(.A1(new_n817), .A2(new_n591), .A3(new_n340), .A4(new_n646), .ZN(new_n843));
  AOI211_X1 g657(.A(new_n843), .B(new_n702), .C1(KEYINPUT49), .C2(new_n733), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n733), .A2(KEYINPUT49), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(KEYINPUT112), .ZN(new_n846));
  INV_X1    g660(.A(new_n711), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n590), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n844), .A2(new_n846), .A3(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT54), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT52), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT113), .ZN(new_n853));
  INV_X1    g667(.A(new_n758), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n854), .A2(new_n666), .A3(new_n667), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n592), .B1(new_n689), .B2(new_n688), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n584), .A2(new_n586), .A3(new_n678), .A4(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  AND4_X1   g672(.A1(new_n853), .A2(new_n858), .A3(new_n711), .A4(new_n778), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n855), .A2(new_n857), .A3(new_n787), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n853), .B1(new_n860), .B2(new_n711), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n693), .B(new_n765), .C1(new_n859), .C2(new_n861), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n724), .A2(KEYINPUT100), .A3(new_n725), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n728), .B1(new_n727), .B2(new_n685), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n852), .B1(new_n862), .B2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n861), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n860), .A2(new_n853), .A3(new_n711), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n765), .A2(new_n693), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n869), .A2(new_n870), .A3(new_n730), .A4(KEYINPUT52), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n866), .A2(new_n871), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n339), .B(new_n734), .C1(new_n669), .C2(new_n661), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n873), .A2(new_n634), .A3(new_n680), .ZN(new_n874));
  INV_X1    g688(.A(new_n483), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n476), .B1(new_n542), .B2(new_n543), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n875), .B1(new_n656), .B2(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n877), .A2(new_n589), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n878), .A2(new_n674), .A3(new_n633), .A4(new_n420), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n745), .A2(new_n879), .A3(new_n760), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n874), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n763), .A2(new_n781), .A3(new_n715), .ZN(new_n882));
  INV_X1    g696(.A(new_n812), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n629), .A2(new_n632), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n691), .A2(new_n538), .A3(new_n534), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n884), .A2(new_n885), .A3(new_n679), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n339), .A2(new_n883), .A3(new_n886), .A4(new_n591), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n797), .A2(new_n882), .A3(new_n887), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n881), .A2(new_n794), .A3(new_n888), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n872), .A2(KEYINPUT53), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(KEYINPUT53), .B1(new_n872), .B2(new_n889), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n851), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n872), .A2(new_n889), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT53), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n872), .A2(new_n889), .A3(KEYINPUT53), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n895), .A2(KEYINPUT54), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n892), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n629), .A2(new_n732), .A3(new_n478), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n785), .A2(new_n899), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n900), .A2(new_n821), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n790), .A2(new_n791), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n589), .B1(new_n902), .B2(new_n789), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT48), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n904), .B(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n849), .A2(new_n656), .A3(new_n900), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n435), .A2(G952), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n689), .B1(new_n819), .B2(new_n820), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n909), .A2(new_n590), .A3(new_n752), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n907), .B(new_n908), .C1(new_n741), .C2(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n906), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n817), .A2(new_n476), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n900), .A2(new_n590), .A3(new_n847), .A4(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n900), .A2(new_n763), .A3(new_n821), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT50), .ZN(new_n917));
  NOR4_X1   g731(.A1(new_n702), .A2(new_n592), .A3(new_n340), .A4(new_n733), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n917), .B1(new_n919), .B2(new_n910), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n752), .A2(new_n590), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n918), .A2(new_n921), .A3(KEYINPUT50), .A4(new_n909), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n916), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n733), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n591), .B1(new_n924), .B2(KEYINPUT114), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n925), .B1(KEYINPUT114), .B2(new_n924), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n837), .A2(new_n838), .A3(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n910), .A2(new_n812), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT51), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n923), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n930), .B1(new_n923), .B2(new_n929), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n912), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(KEYINPUT115), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT115), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n912), .B(new_n935), .C1(new_n931), .C2(new_n932), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n898), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(G952), .A2(G953), .ZN(new_n938));
  OAI211_X1 g752(.A(KEYINPUT116), .B(new_n850), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT116), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n934), .A2(new_n936), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n938), .B1(new_n941), .B2(new_n898), .ZN(new_n942));
  INV_X1    g756(.A(new_n850), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n940), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n939), .A2(new_n944), .ZN(G75));
  NOR2_X1   g759(.A1(new_n435), .A2(G952), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(G902), .B1(new_n890), .B2(new_n891), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(KEYINPUT56), .B1(new_n949), .B2(G210), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n376), .A2(new_n378), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(new_n385), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT55), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n947), .B1(new_n950), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n948), .A2(KEYINPUT117), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT117), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n956), .B(G902), .C1(new_n890), .C2(new_n891), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n955), .A2(new_n417), .A3(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT56), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n953), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT118), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n958), .A2(KEYINPUT118), .A3(new_n960), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n954), .B1(new_n963), .B2(new_n964), .ZN(G51));
  XNOR2_X1  g779(.A(new_n800), .B(KEYINPUT57), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n626), .B1(new_n898), .B2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n806), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n955), .A2(new_n968), .A3(new_n957), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n946), .B1(new_n967), .B2(new_n969), .ZN(G54));
  AND2_X1   g784(.A1(KEYINPUT58), .A2(G475), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n955), .A2(new_n957), .A3(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n972), .A2(new_n469), .A3(new_n468), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n955), .A2(new_n470), .A3(new_n957), .A4(new_n971), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n973), .A2(new_n947), .A3(new_n974), .ZN(G60));
  NAND2_X1  g789(.A1(G478), .A2(G902), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(KEYINPUT119), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT59), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n892), .A2(new_n897), .A3(new_n978), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n649), .A2(new_n654), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n980), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n892), .A2(new_n897), .A3(new_n982), .A4(new_n978), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n981), .A2(new_n947), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(KEYINPUT120), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT120), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n981), .A2(new_n986), .A3(new_n947), .A4(new_n983), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n985), .A2(new_n987), .ZN(G63));
  NAND2_X1  g802(.A1(new_n895), .A2(new_n896), .ZN(new_n989));
  NAND2_X1  g803(.A1(G217), .A2(G902), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(KEYINPUT121), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(KEYINPUT60), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n573), .A2(new_n574), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n946), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(KEYINPUT61), .B1(new_n995), .B2(KEYINPUT122), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n989), .A2(new_n677), .A3(new_n992), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  OAI211_X1 g813(.A(new_n995), .B(new_n997), .C1(KEYINPUT122), .C2(KEYINPUT61), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n999), .A2(new_n1000), .ZN(G66));
  OAI21_X1  g815(.A(G953), .B1(new_n481), .B2(new_n383), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n1002), .B1(new_n881), .B2(G953), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n951), .B1(G898), .B2(new_n435), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1003), .B(new_n1004), .ZN(G69));
  NAND2_X1  g819(.A1(new_n331), .A2(new_n298), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1006), .B(new_n459), .ZN(new_n1007));
  NAND2_X1  g821(.A1(G900), .A2(G953), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n903), .A2(new_n704), .A3(new_n854), .ZN(new_n1009));
  OR2_X1    g823(.A1(new_n1009), .A2(new_n811), .ZN(new_n1010));
  AND4_X1   g824(.A1(new_n794), .A2(new_n1010), .A3(new_n797), .A4(new_n841), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n870), .A2(new_n730), .ZN(new_n1012));
  INV_X1    g826(.A(KEYINPUT123), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n1012), .B(new_n1013), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n1011), .A2(new_n831), .A3(new_n1014), .ZN(new_n1015));
  OAI211_X1 g829(.A(new_n1007), .B(new_n1008), .C1(new_n1015), .C2(G953), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(KEYINPUT125), .ZN(new_n1017));
  INV_X1    g831(.A(new_n1017), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n435), .B1(G227), .B2(G900), .ZN(new_n1019));
  INV_X1    g833(.A(new_n1019), .ZN(new_n1020));
  INV_X1    g834(.A(KEYINPUT62), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1021), .B1(new_n1014), .B2(new_n712), .ZN(new_n1022));
  INV_X1    g836(.A(KEYINPUT124), .ZN(new_n1023));
  XNOR2_X1  g837(.A(new_n1022), .B(new_n1023), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1014), .A2(new_n1021), .A3(new_n712), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n339), .A2(new_n590), .ZN(new_n1026));
  OAI211_X1 g840(.A(new_n697), .B(new_n883), .C1(new_n656), .C2(new_n876), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n841), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1028), .B1(new_n829), .B2(new_n830), .ZN(new_n1029));
  AND2_X1   g843(.A1(new_n1025), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g844(.A(G953), .B1(new_n1024), .B2(new_n1030), .ZN(new_n1031));
  OAI211_X1 g845(.A(new_n1018), .B(new_n1020), .C1(new_n1031), .C2(new_n1007), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1014), .A2(new_n712), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1023), .B1(new_n1033), .B2(KEYINPUT62), .ZN(new_n1034));
  AOI211_X1 g848(.A(KEYINPUT124), .B(new_n1021), .C1(new_n1014), .C2(new_n712), .ZN(new_n1035));
  OAI21_X1  g849(.A(new_n1030), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n1007), .B1(new_n1036), .B2(new_n435), .ZN(new_n1037));
  OAI21_X1  g851(.A(new_n1019), .B1(new_n1037), .B2(new_n1017), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1032), .A2(new_n1038), .ZN(G72));
  XNOR2_X1  g853(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1040));
  NAND2_X1  g854(.A1(G472), .A2(G902), .ZN(new_n1041));
  XNOR2_X1  g855(.A(new_n1040), .B(new_n1041), .ZN(new_n1042));
  INV_X1    g856(.A(new_n881), .ZN(new_n1043));
  OAI21_X1  g857(.A(new_n1042), .B1(new_n1015), .B2(new_n1043), .ZN(new_n1044));
  NOR3_X1   g858(.A1(new_n309), .A2(new_n256), .A3(new_n279), .ZN(new_n1045));
  AOI21_X1  g859(.A(new_n946), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g860(.A(KEYINPUT127), .ZN(new_n1047));
  NAND3_X1  g861(.A1(new_n325), .A2(new_n326), .A3(new_n310), .ZN(new_n1048));
  AND2_X1   g862(.A1(new_n1048), .A2(new_n1042), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n1047), .B1(new_n989), .B2(new_n1049), .ZN(new_n1050));
  AND3_X1   g864(.A1(new_n989), .A2(new_n1047), .A3(new_n1049), .ZN(new_n1051));
  OAI21_X1  g865(.A(new_n1046), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g866(.A(new_n279), .B1(new_n309), .B2(new_n256), .ZN(new_n1053));
  OAI211_X1 g867(.A(new_n1030), .B(new_n881), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1054));
  AOI21_X1  g868(.A(new_n1053), .B1(new_n1054), .B2(new_n1042), .ZN(new_n1055));
  NOR2_X1   g869(.A1(new_n1052), .A2(new_n1055), .ZN(G57));
endmodule


