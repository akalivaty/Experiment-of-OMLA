

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742;

  XNOR2_X1 U373 ( .A(n470), .B(n469), .ZN(n508) );
  XNOR2_X1 U374 ( .A(n724), .B(KEYINPUT75), .ZN(n479) );
  XNOR2_X1 U375 ( .A(n503), .B(n411), .ZN(n726) );
  XNOR2_X1 U376 ( .A(n400), .B(n408), .ZN(n503) );
  XNOR2_X1 U377 ( .A(n399), .B(n406), .ZN(n724) );
  XNOR2_X1 U378 ( .A(n407), .B(G110), .ZN(n399) );
  XNOR2_X1 U379 ( .A(G113), .B(KEYINPUT74), .ZN(n409) );
  BUF_X2 U380 ( .A(n640), .Z(n648) );
  NOR2_X1 U381 ( .A1(G237), .A2(G953), .ZN(n433) );
  INV_X1 U382 ( .A(n585), .ZN(n511) );
  XNOR2_X2 U383 ( .A(G101), .B(KEYINPUT79), .ZN(n407) );
  XNOR2_X2 U384 ( .A(n549), .B(n548), .ZN(n628) );
  AND2_X1 U385 ( .A1(n677), .A2(n676), .ZN(n683) );
  XNOR2_X1 U386 ( .A(KEYINPUT84), .B(G143), .ZN(n415) );
  NAND2_X1 U387 ( .A1(n719), .A2(n372), .ZN(n373) );
  AND2_X1 U388 ( .A1(n367), .A2(n358), .ZN(n738) );
  NOR2_X1 U389 ( .A1(n535), .A2(n630), .ZN(n536) );
  XNOR2_X1 U390 ( .A(n507), .B(KEYINPUT32), .ZN(n381) );
  XNOR2_X1 U391 ( .A(n553), .B(n552), .ZN(n711) );
  AND2_X1 U392 ( .A1(n561), .A2(n560), .ZN(n567) );
  XNOR2_X1 U393 ( .A(n497), .B(n496), .ZN(n677) );
  OR2_X1 U394 ( .A1(n608), .A2(n451), .ZN(n453) );
  XNOR2_X1 U395 ( .A(n415), .B(n414), .ZN(n456) );
  BUF_X1 U396 ( .A(n726), .Z(n351) );
  OR2_X1 U397 ( .A1(n649), .A2(G902), .ZN(n481) );
  XNOR2_X1 U398 ( .A(n474), .B(n473), .ZN(n504) );
  XNOR2_X1 U399 ( .A(G119), .B(G116), .ZN(n408) );
  XNOR2_X1 U400 ( .A(n409), .B(KEYINPUT3), .ZN(n400) );
  NOR2_X1 U401 ( .A1(n608), .A2(n412), .ZN(n376) );
  INV_X1 U402 ( .A(G224), .ZN(n412) );
  XNOR2_X1 U403 ( .A(n390), .B(n389), .ZN(n541) );
  INV_X1 U404 ( .A(KEYINPUT98), .ZN(n389) );
  NAND2_X1 U405 ( .A1(n426), .A2(G902), .ZN(n390) );
  INV_X1 U406 ( .A(G237), .ZN(n420) );
  XNOR2_X1 U407 ( .A(KEYINPUT66), .B(KEYINPUT4), .ZN(n472) );
  XNOR2_X1 U408 ( .A(G146), .B(G125), .ZN(n438) );
  OR2_X1 U409 ( .A1(n555), .A2(n677), .ZN(n583) );
  INV_X1 U410 ( .A(G900), .ZN(n388) );
  XNOR2_X1 U411 ( .A(n368), .B(G101), .ZN(n500) );
  INV_X1 U412 ( .A(KEYINPUT5), .ZN(n368) );
  XNOR2_X1 U413 ( .A(G146), .B(G137), .ZN(n499) );
  XNOR2_X1 U414 ( .A(n597), .B(n361), .ZN(n367) );
  XNOR2_X1 U415 ( .A(n456), .B(G134), .ZN(n474) );
  XNOR2_X1 U416 ( .A(n418), .B(n378), .ZN(n377) );
  XNOR2_X1 U417 ( .A(n479), .B(n726), .ZN(n379) );
  NAND2_X1 U418 ( .A1(n521), .A2(n355), .ZN(n513) );
  INV_X1 U419 ( .A(G953), .ZN(n718) );
  XNOR2_X1 U420 ( .A(n547), .B(n546), .ZN(n392) );
  NOR2_X1 U421 ( .A1(n575), .A2(n554), .ZN(n545) );
  OR2_X1 U422 ( .A1(n635), .A2(G902), .ZN(n505) );
  INV_X1 U423 ( .A(n663), .ZN(n383) );
  NOR2_X1 U424 ( .A1(n593), .A2(n592), .ZN(n594) );
  XOR2_X1 U425 ( .A(KEYINPUT8), .B(KEYINPUT70), .Z(n452) );
  INV_X1 U426 ( .A(G128), .ZN(n414) );
  XNOR2_X1 U427 ( .A(KEYINPUT72), .B(G131), .ZN(n471) );
  XNOR2_X1 U428 ( .A(G143), .B(G113), .ZN(n431) );
  XOR2_X1 U429 ( .A(G104), .B(G140), .Z(n432) );
  XNOR2_X1 U430 ( .A(n374), .B(n413), .ZN(n378) );
  XNOR2_X1 U431 ( .A(n376), .B(n375), .ZN(n374) );
  INV_X1 U432 ( .A(n472), .ZN(n375) );
  XNOR2_X1 U433 ( .A(n391), .B(n359), .ZN(n426) );
  XNOR2_X1 U434 ( .A(KEYINPUT14), .B(KEYINPUT97), .ZN(n391) );
  XNOR2_X1 U435 ( .A(G107), .B(G104), .ZN(n406) );
  XNOR2_X1 U436 ( .A(KEYINPUT71), .B(KEYINPUT10), .ZN(n437) );
  XNOR2_X1 U437 ( .A(G122), .B(KEYINPUT106), .ZN(n447) );
  XOR2_X1 U438 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n448) );
  INV_X1 U439 ( .A(KEYINPUT15), .ZN(n419) );
  NAND2_X1 U440 ( .A1(n719), .A2(n602), .ZN(n603) );
  AND2_X1 U441 ( .A1(n738), .A2(KEYINPUT90), .ZN(n372) );
  NAND2_X1 U442 ( .A1(n551), .A2(n694), .ZN(n553) );
  NAND2_X1 U443 ( .A1(n398), .A2(n712), .ZN(n397) );
  XNOR2_X1 U444 ( .A(n387), .B(n386), .ZN(n569) );
  INV_X1 U445 ( .A(KEYINPUT85), .ZN(n386) );
  NAND2_X1 U446 ( .A1(n385), .A2(n542), .ZN(n387) );
  NAND2_X1 U447 ( .A1(n540), .A2(n364), .ZN(n575) );
  XNOR2_X1 U448 ( .A(n366), .B(n365), .ZN(n364) );
  INV_X1 U449 ( .A(KEYINPUT30), .ZN(n365) );
  INV_X1 U450 ( .A(KEYINPUT19), .ZN(n424) );
  XNOR2_X1 U451 ( .A(n445), .B(G475), .ZN(n570) );
  XNOR2_X1 U452 ( .A(n504), .B(n362), .ZN(n635) );
  XNOR2_X1 U453 ( .A(KEYINPUT16), .B(G122), .ZN(n410) );
  XNOR2_X1 U454 ( .A(KEYINPUT31), .B(KEYINPUT102), .ZN(n525) );
  XNOR2_X1 U455 ( .A(n393), .B(KEYINPUT107), .ZN(n630) );
  XNOR2_X1 U456 ( .A(n532), .B(KEYINPUT93), .ZN(n394) );
  XNOR2_X1 U457 ( .A(n381), .B(n633), .ZN(G21) );
  AND2_X1 U458 ( .A1(n603), .A2(n462), .ZN(n352) );
  AND2_X1 U459 ( .A1(n610), .A2(n644), .ZN(G63) );
  XOR2_X1 U460 ( .A(G140), .B(G137), .Z(n354) );
  AND2_X1 U461 ( .A1(n511), .A2(n683), .ZN(n355) );
  AND2_X1 U462 ( .A1(n508), .A2(n598), .ZN(n356) );
  AND2_X1 U463 ( .A1(n541), .A2(n608), .ZN(n357) );
  AND2_X1 U464 ( .A1(n673), .A2(n624), .ZN(n358) );
  AND2_X1 U465 ( .A1(G234), .A2(G237), .ZN(n359) );
  XOR2_X1 U466 ( .A(KEYINPUT65), .B(KEYINPUT45), .Z(n360) );
  XOR2_X1 U467 ( .A(n596), .B(KEYINPUT73), .Z(n361) );
  XNOR2_X1 U468 ( .A(n504), .B(n354), .ZN(n731) );
  XNOR2_X1 U469 ( .A(n363), .B(n503), .ZN(n362) );
  XNOR2_X1 U470 ( .A(n501), .B(n502), .ZN(n363) );
  NAND2_X1 U471 ( .A1(n681), .A2(n539), .ZN(n366) );
  NAND2_X1 U472 ( .A1(n369), .A2(n518), .ZN(n520) );
  NAND2_X1 U473 ( .A1(n371), .A2(n402), .ZN(n369) );
  INV_X1 U474 ( .A(n370), .ZN(n402) );
  NAND2_X1 U475 ( .A1(n380), .A2(n629), .ZN(n370) );
  INV_X1 U476 ( .A(n632), .ZN(n371) );
  XNOR2_X2 U477 ( .A(n517), .B(KEYINPUT35), .ZN(n632) );
  XNOR2_X2 U478 ( .A(n538), .B(n360), .ZN(n719) );
  NAND2_X1 U479 ( .A1(n604), .A2(n352), .ZN(n395) );
  XNOR2_X2 U480 ( .A(n373), .B(KEYINPUT2), .ZN(n604) );
  NAND2_X1 U481 ( .A1(n508), .A2(n585), .ZN(n532) );
  XNOR2_X2 U482 ( .A(KEYINPUT64), .B(G953), .ZN(n608) );
  XNOR2_X1 U483 ( .A(n379), .B(n377), .ZN(n611) );
  INV_X1 U484 ( .A(n381), .ZN(n380) );
  NAND2_X1 U485 ( .A1(n383), .A2(n382), .ZN(n580) );
  INV_X1 U486 ( .A(n692), .ZN(n382) );
  XNOR2_X2 U487 ( .A(n384), .B(n568), .ZN(n663) );
  NAND2_X1 U488 ( .A1(n567), .A2(n566), .ZN(n384) );
  NAND2_X1 U489 ( .A1(n357), .A2(n388), .ZN(n385) );
  INV_X1 U490 ( .A(n569), .ZN(n554) );
  NAND2_X1 U491 ( .A1(n392), .A2(n666), .ZN(n549) );
  NAND2_X1 U492 ( .A1(n392), .A2(n668), .ZN(n673) );
  XNOR2_X2 U493 ( .A(n560), .B(KEYINPUT1), .ZN(n521) );
  XNOR2_X2 U494 ( .A(n481), .B(G469), .ZN(n560) );
  NAND2_X1 U495 ( .A1(n394), .A2(n534), .ZN(n393) );
  XNOR2_X2 U496 ( .A(n395), .B(KEYINPUT67), .ZN(n640) );
  NAND2_X1 U497 ( .A1(n396), .A2(n404), .ZN(n517) );
  XNOR2_X1 U498 ( .A(n397), .B(n515), .ZN(n396) );
  INV_X1 U499 ( .A(n527), .ZN(n398) );
  NAND2_X1 U500 ( .A1(n604), .A2(n603), .ZN(n675) );
  NAND2_X1 U501 ( .A1(n401), .A2(n402), .ZN(n519) );
  NOR2_X1 U502 ( .A1(n632), .A2(n518), .ZN(n401) );
  NOR2_X1 U503 ( .A1(n506), .A2(n511), .ZN(n403) );
  AND2_X1 U504 ( .A1(n570), .A2(n516), .ZN(n404) );
  AND2_X1 U505 ( .A1(n697), .A2(n676), .ZN(n405) );
  XNOR2_X1 U506 ( .A(n434), .B(G122), .ZN(n435) );
  XNOR2_X1 U507 ( .A(n436), .B(n435), .ZN(n442) );
  INV_X1 U508 ( .A(KEYINPUT34), .ZN(n515) );
  INV_X1 U509 ( .A(n619), .ZN(n620) );
  XNOR2_X1 U510 ( .A(n526), .B(n525), .ZN(n669) );
  XNOR2_X1 U511 ( .A(n410), .B(KEYINPUT77), .ZN(n411) );
  XNOR2_X1 U512 ( .A(n438), .B(KEYINPUT17), .ZN(n413) );
  INV_X1 U513 ( .A(n456), .ZN(n417) );
  XOR2_X1 U514 ( .A(KEYINPUT18), .B(KEYINPUT96), .Z(n416) );
  XNOR2_X1 U515 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U516 ( .A(n419), .B(G902), .ZN(n462) );
  OR2_X2 U517 ( .A1(n611), .A2(n462), .ZN(n422) );
  INV_X1 U518 ( .A(G902), .ZN(n493) );
  NAND2_X1 U519 ( .A1(n493), .A2(n420), .ZN(n423) );
  NAND2_X1 U520 ( .A1(n423), .A2(G210), .ZN(n421) );
  XNOR2_X2 U521 ( .A(n422), .B(n421), .ZN(n543) );
  AND2_X1 U522 ( .A1(n423), .A2(G214), .ZN(n695) );
  NOR2_X2 U523 ( .A1(n543), .A2(n695), .ZN(n425) );
  XNOR2_X1 U524 ( .A(n425), .B(n424), .ZN(n565) );
  NOR2_X1 U525 ( .A1(G898), .A2(n718), .ZN(n727) );
  NAND2_X1 U526 ( .A1(n541), .A2(n727), .ZN(n427) );
  AND2_X1 U527 ( .A1(G952), .A2(n426), .ZN(n706) );
  NAND2_X1 U528 ( .A1(n706), .A2(n718), .ZN(n542) );
  NAND2_X1 U529 ( .A1(n427), .A2(n542), .ZN(n428) );
  NAND2_X1 U530 ( .A1(n565), .A2(n428), .ZN(n430) );
  INV_X1 U531 ( .A(KEYINPUT0), .ZN(n429) );
  XNOR2_X2 U532 ( .A(n430), .B(n429), .ZN(n523) );
  XNOR2_X1 U533 ( .A(KEYINPUT13), .B(KEYINPUT104), .ZN(n444) );
  XNOR2_X1 U534 ( .A(n432), .B(n431), .ZN(n436) );
  XNOR2_X1 U535 ( .A(n433), .B(KEYINPUT80), .ZN(n498) );
  NAND2_X1 U536 ( .A1(n498), .A2(G214), .ZN(n434) );
  XNOR2_X1 U537 ( .A(n438), .B(n437), .ZN(n732) );
  XOR2_X1 U538 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n439) );
  XNOR2_X1 U539 ( .A(n471), .B(n439), .ZN(n440) );
  XNOR2_X1 U540 ( .A(n732), .B(n440), .ZN(n441) );
  XNOR2_X1 U541 ( .A(n442), .B(n441), .ZN(n641) );
  NOR2_X1 U542 ( .A1(G902), .A2(n641), .ZN(n443) );
  XNOR2_X1 U543 ( .A(n444), .B(n443), .ZN(n445) );
  INV_X1 U544 ( .A(n570), .ZN(n461) );
  XNOR2_X1 U545 ( .A(G116), .B(G107), .ZN(n446) );
  XNOR2_X1 U546 ( .A(n446), .B(KEYINPUT105), .ZN(n450) );
  XNOR2_X1 U547 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U548 ( .A(n450), .B(n449), .Z(n455) );
  INV_X1 U549 ( .A(G234), .ZN(n451) );
  XNOR2_X1 U550 ( .A(n453), .B(n452), .ZN(n482) );
  NAND2_X1 U551 ( .A1(n482), .A2(G217), .ZN(n454) );
  XNOR2_X1 U552 ( .A(n455), .B(n454), .ZN(n458) );
  INV_X1 U553 ( .A(n474), .ZN(n457) );
  XNOR2_X1 U554 ( .A(n458), .B(n457), .ZN(n606) );
  NAND2_X1 U555 ( .A1(n606), .A2(n493), .ZN(n460) );
  INV_X1 U556 ( .A(G478), .ZN(n459) );
  XNOR2_X1 U557 ( .A(n460), .B(n459), .ZN(n571) );
  AND2_X1 U558 ( .A1(n461), .A2(n571), .ZN(n697) );
  INV_X1 U559 ( .A(n462), .ZN(n605) );
  NAND2_X1 U560 ( .A1(n605), .A2(G234), .ZN(n463) );
  XNOR2_X1 U561 ( .A(n463), .B(KEYINPUT20), .ZN(n494) );
  INV_X1 U562 ( .A(n494), .ZN(n465) );
  INV_X1 U563 ( .A(G221), .ZN(n464) );
  OR2_X1 U564 ( .A1(n465), .A2(n464), .ZN(n467) );
  INV_X1 U565 ( .A(KEYINPUT21), .ZN(n466) );
  XNOR2_X1 U566 ( .A(n467), .B(n466), .ZN(n676) );
  NAND2_X1 U567 ( .A1(n523), .A2(n405), .ZN(n470) );
  INV_X1 U568 ( .A(KEYINPUT68), .ZN(n468) );
  XNOR2_X1 U569 ( .A(n468), .B(KEYINPUT22), .ZN(n469) );
  XNOR2_X1 U570 ( .A(n472), .B(n471), .ZN(n473) );
  INV_X1 U571 ( .A(G227), .ZN(n733) );
  OR2_X1 U572 ( .A1(n608), .A2(n733), .ZN(n477) );
  XNOR2_X1 U573 ( .A(G146), .B(KEYINPUT81), .ZN(n475) );
  XNOR2_X1 U574 ( .A(n475), .B(KEYINPUT82), .ZN(n476) );
  XNOR2_X1 U575 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U576 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U577 ( .A(n731), .B(n480), .ZN(n649) );
  NAND2_X1 U578 ( .A1(n482), .A2(G221), .ZN(n487) );
  XNOR2_X1 U579 ( .A(G128), .B(G110), .ZN(n484) );
  XNOR2_X1 U580 ( .A(G119), .B(KEYINPUT24), .ZN(n483) );
  XNOR2_X1 U581 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U582 ( .A(n485), .B(n354), .ZN(n486) );
  XNOR2_X1 U583 ( .A(n487), .B(n486), .ZN(n492) );
  XNOR2_X1 U584 ( .A(KEYINPUT100), .B(KEYINPUT101), .ZN(n489) );
  XNOR2_X1 U585 ( .A(KEYINPUT23), .B(KEYINPUT88), .ZN(n488) );
  XNOR2_X1 U586 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U587 ( .A(n732), .B(n490), .ZN(n491) );
  XNOR2_X1 U588 ( .A(n492), .B(n491), .ZN(n619) );
  NAND2_X1 U589 ( .A1(n619), .A2(n493), .ZN(n497) );
  AND2_X1 U590 ( .A1(n494), .A2(G217), .ZN(n495) );
  XNOR2_X1 U591 ( .A(n495), .B(KEYINPUT25), .ZN(n496) );
  INV_X1 U592 ( .A(n677), .ZN(n533) );
  NAND2_X1 U593 ( .A1(n521), .A2(n533), .ZN(n506) );
  NAND2_X1 U594 ( .A1(G210), .A2(n498), .ZN(n502) );
  XNOR2_X1 U595 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X2 U596 ( .A(n505), .B(G472), .ZN(n681) );
  XNOR2_X1 U597 ( .A(n681), .B(KEYINPUT6), .ZN(n585) );
  AND2_X1 U598 ( .A1(n508), .A2(n403), .ZN(n507) );
  XNOR2_X1 U599 ( .A(n356), .B(KEYINPUT108), .ZN(n510) );
  NOR2_X1 U600 ( .A1(n681), .A2(n677), .ZN(n509) );
  NAND2_X1 U601 ( .A1(n510), .A2(n509), .ZN(n629) );
  XNOR2_X1 U602 ( .A(KEYINPUT109), .B(KEYINPUT33), .ZN(n512) );
  XNOR2_X1 U603 ( .A(n513), .B(n512), .ZN(n514) );
  INV_X1 U604 ( .A(n514), .ZN(n712) );
  XNOR2_X1 U605 ( .A(n523), .B(KEYINPUT99), .ZN(n527) );
  INV_X1 U606 ( .A(n571), .ZN(n516) );
  INV_X1 U607 ( .A(KEYINPUT44), .ZN(n518) );
  NAND2_X1 U608 ( .A1(n520), .A2(n519), .ZN(n537) );
  INV_X1 U609 ( .A(n521), .ZN(n598) );
  NAND2_X1 U610 ( .A1(n681), .A2(n683), .ZN(n522) );
  NOR2_X1 U611 ( .A1(n598), .A2(n522), .ZN(n687) );
  BUF_X1 U612 ( .A(n523), .Z(n524) );
  NAND2_X1 U613 ( .A1(n687), .A2(n524), .ZN(n526) );
  AND2_X1 U614 ( .A1(n560), .A2(n683), .ZN(n540) );
  INV_X1 U615 ( .A(n681), .ZN(n528) );
  NAND2_X1 U616 ( .A1(n540), .A2(n528), .ZN(n529) );
  NOR2_X1 U617 ( .A1(n527), .A2(n529), .ZN(n658) );
  OR2_X1 U618 ( .A1(n669), .A2(n658), .ZN(n530) );
  XNOR2_X1 U619 ( .A(n530), .B(KEYINPUT103), .ZN(n531) );
  NOR2_X1 U620 ( .A1(n570), .A2(n571), .ZN(n668) );
  AND2_X1 U621 ( .A1(n570), .A2(n571), .ZN(n666) );
  NOR2_X1 U622 ( .A1(n668), .A2(n666), .ZN(n692) );
  NOR2_X1 U623 ( .A1(n531), .A2(n692), .ZN(n535) );
  NOR2_X1 U624 ( .A1(n521), .A2(n533), .ZN(n534) );
  NAND2_X1 U625 ( .A1(n537), .A2(n536), .ZN(n538) );
  INV_X1 U626 ( .A(n695), .ZN(n539) );
  BUF_X1 U627 ( .A(n543), .Z(n573) );
  XNOR2_X1 U628 ( .A(KEYINPUT78), .B(KEYINPUT38), .ZN(n544) );
  XNOR2_X1 U629 ( .A(n573), .B(n544), .ZN(n694) );
  NAND2_X1 U630 ( .A1(n545), .A2(n694), .ZN(n547) );
  XNOR2_X1 U631 ( .A(KEYINPUT76), .B(KEYINPUT39), .ZN(n546) );
  XOR2_X1 U632 ( .A(KEYINPUT111), .B(KEYINPUT40), .Z(n548) );
  INV_X1 U633 ( .A(n697), .ZN(n550) );
  NOR2_X1 U634 ( .A1(n550), .A2(n695), .ZN(n551) );
  XNOR2_X1 U635 ( .A(KEYINPUT112), .B(KEYINPUT41), .ZN(n552) );
  NAND2_X1 U636 ( .A1(n569), .A2(n676), .ZN(n555) );
  INV_X1 U637 ( .A(n583), .ZN(n556) );
  NAND2_X1 U638 ( .A1(n556), .A2(n681), .ZN(n559) );
  INV_X1 U639 ( .A(KEYINPUT110), .ZN(n557) );
  XNOR2_X1 U640 ( .A(n557), .B(KEYINPUT28), .ZN(n558) );
  XNOR2_X1 U641 ( .A(n559), .B(n558), .ZN(n561) );
  NAND2_X1 U642 ( .A1(n711), .A2(n567), .ZN(n562) );
  XNOR2_X1 U643 ( .A(n562), .B(KEYINPUT42), .ZN(n631) );
  NAND2_X1 U644 ( .A1(n628), .A2(n631), .ZN(n564) );
  XOR2_X1 U645 ( .A(KEYINPUT92), .B(KEYINPUT46), .Z(n563) );
  XNOR2_X1 U646 ( .A(n564), .B(n563), .ZN(n595) );
  BUF_X1 U647 ( .A(n565), .Z(n566) );
  INV_X1 U648 ( .A(KEYINPUT83), .ZN(n568) );
  NAND2_X1 U649 ( .A1(n580), .A2(KEYINPUT47), .ZN(n578) );
  NAND2_X1 U650 ( .A1(n570), .A2(n569), .ZN(n572) );
  NOR2_X1 U651 ( .A1(n572), .A2(n571), .ZN(n574) );
  INV_X1 U652 ( .A(n573), .ZN(n587) );
  NAND2_X1 U653 ( .A1(n574), .A2(n587), .ZN(n576) );
  NOR2_X1 U654 ( .A1(n576), .A2(n575), .ZN(n623) );
  XNOR2_X1 U655 ( .A(n623), .B(KEYINPUT87), .ZN(n577) );
  NAND2_X1 U656 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U657 ( .A(n579), .B(KEYINPUT86), .ZN(n593) );
  INV_X1 U658 ( .A(n580), .ZN(n582) );
  XNOR2_X1 U659 ( .A(KEYINPUT47), .B(KEYINPUT69), .ZN(n581) );
  NAND2_X1 U660 ( .A1(n582), .A2(n581), .ZN(n591) );
  NOR2_X1 U661 ( .A1(n583), .A2(n695), .ZN(n584) );
  NAND2_X1 U662 ( .A1(n666), .A2(n584), .ZN(n586) );
  NOR2_X1 U663 ( .A1(n586), .A2(n585), .ZN(n599) );
  NAND2_X1 U664 ( .A1(n599), .A2(n587), .ZN(n589) );
  XOR2_X1 U665 ( .A(KEYINPUT94), .B(KEYINPUT36), .Z(n588) );
  XNOR2_X1 U666 ( .A(n589), .B(n588), .ZN(n590) );
  NAND2_X1 U667 ( .A1(n590), .A2(n521), .ZN(n671) );
  NAND2_X1 U668 ( .A1(n591), .A2(n671), .ZN(n592) );
  NAND2_X1 U669 ( .A1(n595), .A2(n594), .ZN(n597) );
  XNOR2_X1 U670 ( .A(KEYINPUT91), .B(KEYINPUT48), .ZN(n596) );
  NAND2_X1 U671 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U672 ( .A(n600), .B(KEYINPUT43), .ZN(n601) );
  NAND2_X1 U673 ( .A1(n601), .A2(n573), .ZN(n624) );
  NOR2_X1 U674 ( .A1(n738), .A2(KEYINPUT90), .ZN(n602) );
  NAND2_X1 U675 ( .A1(n648), .A2(G478), .ZN(n607) );
  XNOR2_X1 U676 ( .A(n607), .B(n606), .ZN(n610) );
  INV_X1 U677 ( .A(n608), .ZN(n740) );
  NOR2_X1 U678 ( .A1(n740), .A2(G952), .ZN(n609) );
  XNOR2_X1 U679 ( .A(n609), .B(KEYINPUT95), .ZN(n644) );
  INV_X1 U680 ( .A(n644), .ZN(n655) );
  NAND2_X1 U681 ( .A1(n640), .A2(G210), .ZN(n615) );
  BUF_X1 U682 ( .A(n611), .Z(n612) );
  XNOR2_X1 U683 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n613) );
  XNOR2_X1 U684 ( .A(n612), .B(n613), .ZN(n614) );
  XNOR2_X1 U685 ( .A(n615), .B(n614), .ZN(n616) );
  NAND2_X1 U686 ( .A1(n616), .A2(n644), .ZN(n618) );
  INV_X1 U687 ( .A(KEYINPUT56), .ZN(n617) );
  XNOR2_X1 U688 ( .A(n618), .B(n617), .ZN(G51) );
  NAND2_X1 U689 ( .A1(n648), .A2(G217), .ZN(n621) );
  XNOR2_X1 U690 ( .A(n621), .B(n620), .ZN(n622) );
  NOR2_X1 U691 ( .A1(n622), .A2(n655), .ZN(G66) );
  XOR2_X1 U692 ( .A(G143), .B(n623), .Z(G45) );
  XNOR2_X1 U693 ( .A(n624), .B(G140), .ZN(G42) );
  XOR2_X1 U694 ( .A(G128), .B(KEYINPUT29), .Z(n627) );
  INV_X1 U695 ( .A(n668), .ZN(n625) );
  NOR2_X1 U696 ( .A1(n663), .A2(n625), .ZN(n626) );
  XOR2_X1 U697 ( .A(n627), .B(n626), .Z(G30) );
  XNOR2_X1 U698 ( .A(n628), .B(G131), .ZN(G33) );
  XNOR2_X1 U699 ( .A(n629), .B(G110), .ZN(G12) );
  XOR2_X1 U700 ( .A(n630), .B(G101), .Z(G3) );
  XNOR2_X1 U701 ( .A(n631), .B(G137), .ZN(G39) );
  XOR2_X1 U702 ( .A(n632), .B(G122), .Z(G24) );
  XNOR2_X1 U703 ( .A(G119), .B(KEYINPUT127), .ZN(n633) );
  NAND2_X1 U704 ( .A1(n640), .A2(G472), .ZN(n637) );
  XNOR2_X1 U705 ( .A(KEYINPUT113), .B(KEYINPUT62), .ZN(n634) );
  XNOR2_X1 U706 ( .A(n635), .B(n634), .ZN(n636) );
  XNOR2_X1 U707 ( .A(n637), .B(n636), .ZN(n638) );
  NAND2_X1 U708 ( .A1(n638), .A2(n644), .ZN(n639) );
  XNOR2_X1 U709 ( .A(n639), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U710 ( .A1(n640), .A2(G475), .ZN(n643) );
  XNOR2_X1 U711 ( .A(n641), .B(KEYINPUT59), .ZN(n642) );
  XNOR2_X1 U712 ( .A(n643), .B(n642), .ZN(n645) );
  NAND2_X1 U713 ( .A1(n645), .A2(n644), .ZN(n647) );
  XOR2_X1 U714 ( .A(KEYINPUT124), .B(KEYINPUT60), .Z(n646) );
  XNOR2_X1 U715 ( .A(n647), .B(n646), .ZN(G60) );
  NAND2_X1 U716 ( .A1(n648), .A2(G469), .ZN(n654) );
  XOR2_X1 U717 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n651) );
  XNOR2_X1 U718 ( .A(KEYINPUT123), .B(KEYINPUT122), .ZN(n650) );
  XOR2_X1 U719 ( .A(n651), .B(n650), .Z(n652) );
  XNOR2_X1 U720 ( .A(n649), .B(n652), .ZN(n653) );
  XNOR2_X1 U721 ( .A(n654), .B(n653), .ZN(n656) );
  NOR2_X1 U722 ( .A1(n656), .A2(n655), .ZN(G54) );
  NAND2_X1 U723 ( .A1(n666), .A2(n658), .ZN(n657) );
  XNOR2_X1 U724 ( .A(G104), .B(n657), .ZN(G6) );
  XOR2_X1 U725 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n660) );
  NAND2_X1 U726 ( .A1(n658), .A2(n668), .ZN(n659) );
  XNOR2_X1 U727 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U728 ( .A(G107), .B(n661), .ZN(G9) );
  INV_X1 U729 ( .A(n666), .ZN(n662) );
  NOR2_X1 U730 ( .A1(n663), .A2(n662), .ZN(n664) );
  XOR2_X1 U731 ( .A(KEYINPUT114), .B(n664), .Z(n665) );
  XNOR2_X1 U732 ( .A(G146), .B(n665), .ZN(G48) );
  NAND2_X1 U733 ( .A1(n669), .A2(n666), .ZN(n667) );
  XNOR2_X1 U734 ( .A(n667), .B(G113), .ZN(G15) );
  NAND2_X1 U735 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U736 ( .A(n670), .B(G116), .ZN(G18) );
  XOR2_X1 U737 ( .A(G125), .B(n671), .Z(n672) );
  XNOR2_X1 U738 ( .A(n672), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U739 ( .A(G134), .B(n673), .Z(n674) );
  XNOR2_X1 U740 ( .A(n674), .B(KEYINPUT115), .ZN(G36) );
  XNOR2_X1 U741 ( .A(KEYINPUT121), .B(KEYINPUT53), .ZN(n717) );
  XNOR2_X1 U742 ( .A(n675), .B(KEYINPUT89), .ZN(n710) );
  NOR2_X1 U743 ( .A1(n677), .A2(n676), .ZN(n678) );
  XOR2_X1 U744 ( .A(KEYINPUT116), .B(n678), .Z(n679) );
  XNOR2_X1 U745 ( .A(n679), .B(KEYINPUT49), .ZN(n680) );
  NOR2_X1 U746 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U747 ( .A(KEYINPUT117), .B(n682), .ZN(n686) );
  NOR2_X1 U748 ( .A1(n521), .A2(n683), .ZN(n684) );
  XNOR2_X1 U749 ( .A(n684), .B(KEYINPUT50), .ZN(n685) );
  NOR2_X1 U750 ( .A1(n686), .A2(n685), .ZN(n688) );
  NOR2_X1 U751 ( .A1(n688), .A2(n687), .ZN(n690) );
  XNOR2_X1 U752 ( .A(KEYINPUT118), .B(KEYINPUT51), .ZN(n689) );
  XNOR2_X1 U753 ( .A(n690), .B(n689), .ZN(n691) );
  NAND2_X1 U754 ( .A1(n691), .A2(n711), .ZN(n704) );
  NOR2_X1 U755 ( .A1(n692), .A2(n695), .ZN(n693) );
  NAND2_X1 U756 ( .A1(n693), .A2(n694), .ZN(n700) );
  INV_X1 U757 ( .A(n694), .ZN(n696) );
  NAND2_X1 U758 ( .A1(n696), .A2(n695), .ZN(n698) );
  NAND2_X1 U759 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U760 ( .A1(n700), .A2(n699), .ZN(n701) );
  XOR2_X1 U761 ( .A(KEYINPUT119), .B(n701), .Z(n702) );
  NAND2_X1 U762 ( .A1(n702), .A2(n712), .ZN(n703) );
  NAND2_X1 U763 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U764 ( .A(n705), .B(KEYINPUT52), .ZN(n707) );
  NAND2_X1 U765 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U766 ( .A1(n708), .A2(n718), .ZN(n709) );
  NOR2_X1 U767 ( .A1(n710), .A2(n709), .ZN(n715) );
  NAND2_X1 U768 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U769 ( .A(n713), .B(KEYINPUT120), .ZN(n714) );
  NAND2_X1 U770 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U771 ( .A(n717), .B(n716), .ZN(G75) );
  NAND2_X1 U772 ( .A1(n719), .A2(n718), .ZN(n723) );
  NAND2_X1 U773 ( .A1(G953), .A2(G224), .ZN(n720) );
  XNOR2_X1 U774 ( .A(KEYINPUT61), .B(n720), .ZN(n721) );
  NAND2_X1 U775 ( .A1(n721), .A2(G898), .ZN(n722) );
  NAND2_X1 U776 ( .A1(n723), .A2(n722), .ZN(n730) );
  XOR2_X1 U777 ( .A(KEYINPUT125), .B(n724), .Z(n725) );
  XNOR2_X1 U778 ( .A(n351), .B(n725), .ZN(n728) );
  NOR2_X1 U779 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U780 ( .A(n730), .B(n729), .ZN(G69) );
  XOR2_X1 U781 ( .A(n732), .B(n731), .Z(n736) );
  XNOR2_X1 U782 ( .A(n736), .B(n733), .ZN(n734) );
  NAND2_X1 U783 ( .A1(n734), .A2(G900), .ZN(n735) );
  NAND2_X1 U784 ( .A1(n735), .A2(G953), .ZN(n742) );
  XNOR2_X1 U785 ( .A(n736), .B(KEYINPUT126), .ZN(n737) );
  XNOR2_X1 U786 ( .A(n738), .B(n737), .ZN(n739) );
  NAND2_X1 U787 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U788 ( .A1(n742), .A2(n741), .ZN(G72) );
endmodule

