//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 0 1 1 1 1 0 1 0 1 0 0 0 1 1 0 1 1 0 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1 1 0 1 0 1 1 0 0 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n768, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n856,
    new_n857, new_n858, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992;
  INV_X1    g000(.A(G190gat), .ZN(new_n202));
  AND2_X1   g001(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT28), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n206), .A2(KEYINPUT66), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n206), .A2(KEYINPUT66), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n207), .B(new_n202), .C1(new_n204), .C2(new_n203), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT67), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT26), .ZN(new_n216));
  NAND2_X1  g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT26), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n214), .A2(KEYINPUT67), .A3(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n216), .A2(new_n217), .A3(new_n219), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n212), .A2(new_n213), .A3(new_n220), .ZN(new_n221));
  XOR2_X1   g020(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n222));
  NAND2_X1  g021(.A1(new_n214), .A2(KEYINPUT23), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT24), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n224), .A2(G183gat), .A3(G190gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n223), .A2(new_n225), .A3(new_n217), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT23), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n227), .B1(G169gat), .B2(G176gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n213), .A2(KEYINPUT24), .ZN(new_n229));
  NOR2_X1   g028(.A1(G183gat), .A2(G190gat), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n228), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n222), .B1(new_n226), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT65), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n213), .A2(new_n233), .A3(new_n224), .ZN(new_n234));
  INV_X1    g033(.A(new_n230), .ZN(new_n235));
  OAI211_X1 g034(.A(G183gat), .B(G190gat), .C1(KEYINPUT65), .C2(KEYINPUT24), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n234), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n217), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n238), .B1(KEYINPUT23), .B2(new_n214), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n237), .A2(new_n239), .A3(KEYINPUT25), .A4(new_n228), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n232), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n221), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(G120gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(G113gat), .ZN(new_n244));
  INV_X1    g043(.A(G113gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(G120gat), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT1), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(G127gat), .ZN(new_n249));
  INV_X1    g048(.A(G134gat), .ZN(new_n250));
  OR2_X1    g049(.A1(new_n250), .A2(KEYINPUT68), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(KEYINPUT68), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n249), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  OR2_X1    g052(.A1(KEYINPUT69), .A2(G127gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(KEYINPUT69), .A2(G127gat), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n250), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n248), .B1(new_n253), .B2(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(G127gat), .B(G134gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n247), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT70), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT70), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n247), .A2(new_n261), .A3(new_n258), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n257), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n242), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT71), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n263), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n267), .A2(new_n241), .A3(new_n221), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n242), .A2(KEYINPUT71), .A3(new_n263), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n266), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(G227gat), .ZN(new_n271));
  INV_X1    g070(.A(G233gat), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT34), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n270), .A2(new_n273), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n275), .B1(new_n276), .B2(KEYINPUT32), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT32), .ZN(new_n278));
  AOI211_X1 g077(.A(new_n278), .B(KEYINPUT34), .C1(new_n270), .C2(new_n273), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n274), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  AND3_X1   g079(.A1(new_n242), .A2(KEYINPUT71), .A3(new_n263), .ZN(new_n281));
  AOI21_X1  g080(.A(KEYINPUT71), .B1(new_n242), .B2(new_n263), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n242), .A2(new_n263), .ZN(new_n283));
  NOR3_X1   g082(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n273), .ZN(new_n285));
  OAI21_X1  g084(.A(KEYINPUT32), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT34), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n276), .A2(KEYINPUT32), .A3(new_n275), .ZN(new_n288));
  INV_X1    g087(.A(new_n274), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT33), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(G15gat), .B(G43gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n293), .B(G71gat), .ZN(new_n294));
  INV_X1    g093(.A(G99gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n294), .B(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  AND3_X1   g097(.A1(new_n280), .A2(new_n290), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n298), .B1(new_n280), .B2(new_n290), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n301), .A2(KEYINPUT36), .ZN(new_n302));
  NOR3_X1   g101(.A1(new_n277), .A2(new_n279), .A3(new_n274), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n289), .B1(new_n287), .B2(new_n288), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n297), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n280), .A2(new_n290), .A3(new_n298), .ZN(new_n306));
  AND3_X1   g105(.A1(new_n305), .A2(KEYINPUT36), .A3(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(G141gat), .B(G148gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(G155gat), .A2(G162gat), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT2), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n308), .B1(new_n309), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT78), .ZN(new_n315));
  INV_X1    g114(.A(new_n309), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n316), .A2(new_n310), .ZN(new_n317));
  XOR2_X1   g116(.A(KEYINPUT77), .B(KEYINPUT2), .Z(new_n318));
  OAI211_X1 g117(.A(new_n315), .B(new_n317), .C1(new_n318), .C2(new_n308), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  XOR2_X1   g119(.A(G141gat), .B(G148gat), .Z(new_n321));
  XNOR2_X1  g120(.A(KEYINPUT77), .B(KEYINPUT2), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n315), .B1(new_n323), .B2(new_n317), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n314), .B1(new_n320), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(KEYINPUT4), .B1(new_n325), .B2(new_n263), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n317), .B1(new_n318), .B2(new_n308), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT78), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n313), .B1(new_n328), .B2(new_n319), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT4), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n267), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n326), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(G225gat), .A2(G233gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n333), .B(KEYINPUT79), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n325), .A2(KEYINPUT3), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT3), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n329), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n336), .A2(new_n263), .A3(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n332), .A2(new_n335), .A3(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT5), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n325), .B(new_n263), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(new_n334), .ZN(new_n344));
  AND2_X1   g143(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n342), .B1(new_n345), .B2(new_n341), .ZN(new_n346));
  XNOR2_X1  g145(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n347));
  XNOR2_X1  g146(.A(G1gat), .B(G29gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n347), .B(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G57gat), .B(G85gat), .ZN(new_n350));
  XOR2_X1   g149(.A(new_n349), .B(new_n350), .Z(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT6), .B1(new_n346), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n353), .B1(new_n352), .B2(new_n346), .ZN(new_n354));
  INV_X1    g153(.A(new_n342), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n341), .B1(new_n340), .B2(new_n344), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n357), .A2(KEYINPUT6), .A3(new_n351), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT76), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT29), .B1(new_n221), .B2(new_n241), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT75), .ZN(new_n361));
  AND2_X1   g160(.A1(G226gat), .A2(G233gat), .ZN(new_n362));
  NOR3_X1   g161(.A1(new_n360), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT29), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n362), .B1(new_n242), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT75), .B1(new_n242), .B2(new_n362), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n363), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(KEYINPUT73), .B(G218gat), .ZN(new_n369));
  AOI21_X1  g168(.A(KEYINPUT22), .B1(new_n369), .B2(G211gat), .ZN(new_n370));
  INV_X1    g169(.A(G197gat), .ZN(new_n371));
  AND2_X1   g170(.A1(KEYINPUT72), .A2(G204gat), .ZN(new_n372));
  NOR2_X1   g171(.A1(KEYINPUT72), .A2(G204gat), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT72), .ZN(new_n375));
  INV_X1    g174(.A(G204gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(KEYINPUT72), .A2(G204gat), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n377), .A2(G197gat), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n374), .A2(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(G211gat), .B1(new_n370), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(G218gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT73), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT73), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(G218gat), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n383), .A2(new_n385), .A3(G211gat), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT22), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(G211gat), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n388), .A2(new_n389), .A3(new_n379), .A4(new_n374), .ZN(new_n390));
  AND3_X1   g189(.A1(new_n381), .A2(G218gat), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(G218gat), .B1(new_n381), .B2(new_n390), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n359), .B1(new_n368), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n242), .A2(new_n362), .ZN(new_n395));
  OR2_X1    g194(.A1(new_n395), .A2(KEYINPUT74), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n395), .B(KEYINPUT74), .C1(new_n362), .C2(new_n360), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n396), .A2(new_n397), .A3(new_n393), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n395), .B(new_n361), .C1(new_n362), .C2(new_n360), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n365), .A2(KEYINPUT75), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n381), .A2(new_n390), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(new_n382), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n381), .A2(G218gat), .A3(new_n390), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n401), .A2(KEYINPUT76), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n394), .A2(new_n398), .A3(new_n406), .ZN(new_n407));
  XOR2_X1   g206(.A(G8gat), .B(G36gat), .Z(new_n408));
  XNOR2_X1  g207(.A(new_n408), .B(G64gat), .ZN(new_n409));
  INV_X1    g208(.A(G92gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n411), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n394), .A2(new_n398), .A3(new_n406), .A4(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n412), .A2(KEYINPUT30), .A3(new_n414), .ZN(new_n415));
  OR3_X1    g214(.A1(new_n407), .A2(KEYINPUT30), .A3(new_n411), .ZN(new_n416));
  AOI22_X1  g215(.A1(new_n354), .A2(new_n358), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(G22gat), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n364), .B1(new_n391), .B2(new_n392), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n329), .B1(new_n419), .B2(new_n337), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT29), .B1(new_n329), .B2(new_n337), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n405), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(G228gat), .ZN(new_n423));
  OAI22_X1  g222(.A1(new_n420), .A2(new_n422), .B1(new_n423), .B2(new_n272), .ZN(new_n424));
  INV_X1    g223(.A(new_n421), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(new_n393), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n423), .A2(new_n272), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT3), .B1(new_n405), .B2(new_n364), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n426), .B(new_n427), .C1(new_n428), .C2(new_n329), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n418), .B1(new_n424), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n424), .A2(new_n429), .A3(new_n418), .ZN(new_n432));
  XOR2_X1   g231(.A(G78gat), .B(G106gat), .Z(new_n433));
  XNOR2_X1  g232(.A(new_n433), .B(KEYINPUT31), .ZN(new_n434));
  INV_X1    g233(.A(G50gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n434), .B(new_n435), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n436), .A2(KEYINPUT81), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n432), .A2(new_n437), .ZN(new_n438));
  AND2_X1   g237(.A1(new_n432), .A2(KEYINPUT82), .ZN(new_n439));
  INV_X1    g238(.A(new_n436), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n431), .B(new_n438), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n438), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n440), .B1(new_n432), .B2(KEYINPUT82), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n430), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  OAI22_X1  g244(.A1(new_n302), .A2(new_n307), .B1(new_n417), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT86), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT76), .B1(new_n401), .B2(new_n405), .ZN(new_n449));
  AOI211_X1 g248(.A(new_n359), .B(new_n393), .C1(new_n399), .C2(new_n400), .ZN(new_n450));
  INV_X1    g249(.A(new_n398), .ZN(new_n451));
  NOR3_X1   g250(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT37), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n448), .B(new_n411), .C1(new_n452), .C2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n452), .A2(new_n453), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n407), .A2(KEYINPUT37), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n448), .B1(new_n457), .B2(new_n411), .ZN(new_n458));
  OAI21_X1  g257(.A(KEYINPUT38), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  OAI211_X1 g258(.A(KEYINPUT84), .B(new_n342), .C1(new_n345), .C2(new_n341), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT84), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n461), .B1(new_n355), .B2(new_n356), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n460), .A2(new_n462), .A3(new_n351), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n353), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n357), .A2(KEYINPUT6), .A3(new_n351), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT38), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n453), .B1(new_n401), .B2(new_n393), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n396), .A2(new_n397), .A3(new_n405), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n413), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n466), .B(new_n469), .C1(new_n407), .C2(KEYINPUT37), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n464), .A2(new_n465), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n459), .A2(new_n471), .A3(new_n414), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n335), .B1(new_n332), .B2(new_n339), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT39), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n352), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n343), .A2(new_n334), .ZN(new_n477));
  NOR3_X1   g276(.A1(new_n473), .A2(new_n477), .A3(new_n474), .ZN(new_n478));
  OAI21_X1  g277(.A(KEYINPUT83), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT40), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OAI211_X1 g280(.A(KEYINPUT83), .B(KEYINPUT40), .C1(new_n476), .C2(new_n478), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n483), .A2(new_n415), .A3(new_n416), .A4(new_n463), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT85), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n415), .A2(new_n416), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n487), .A2(KEYINPUT85), .A3(new_n463), .A4(new_n483), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n472), .A2(new_n445), .A3(new_n486), .A4(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT87), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n490), .B1(new_n299), .B2(new_n300), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n305), .A2(KEYINPUT87), .A3(new_n306), .ZN(new_n492));
  AND3_X1   g291(.A1(new_n491), .A2(new_n445), .A3(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT35), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n415), .A2(new_n416), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n464), .A2(new_n465), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n493), .A2(new_n494), .A3(new_n495), .A4(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n417), .A2(new_n445), .A3(new_n301), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT35), .ZN(new_n499));
  AOI22_X1  g298(.A1(new_n447), .A2(new_n489), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G15gat), .B(G22gat), .ZN(new_n501));
  OR2_X1    g300(.A1(new_n501), .A2(G1gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT90), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT16), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n501), .B1(new_n504), .B2(G1gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n503), .A2(new_n506), .A3(G8gat), .ZN(new_n507));
  INV_X1    g306(.A(G8gat), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n502), .B(new_n505), .C1(KEYINPUT90), .C2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT94), .ZN(new_n511));
  XNOR2_X1  g310(.A(G57gat), .B(G64gat), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  XOR2_X1   g313(.A(G71gat), .B(G78gat), .Z(new_n515));
  OR2_X1    g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n515), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n510), .B1(KEYINPUT21), .B2(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n519), .B(KEYINPUT96), .ZN(new_n520));
  NAND2_X1  g319(.A1(G231gat), .A2(G233gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n520), .B(new_n521), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n518), .A2(KEYINPUT21), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n522), .B(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G183gat), .B(G211gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(KEYINPUT95), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n526), .B(KEYINPUT19), .ZN(new_n527));
  XOR2_X1   g326(.A(G127gat), .B(G155gat), .Z(new_n528));
  XNOR2_X1  g327(.A(new_n528), .B(KEYINPUT20), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n527), .B(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n524), .B(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  XOR2_X1   g331(.A(G43gat), .B(G50gat), .Z(new_n533));
  INV_X1    g332(.A(KEYINPUT89), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(G29gat), .ZN(new_n536));
  INV_X1    g335(.A(G36gat), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n536), .A2(new_n537), .A3(KEYINPUT14), .ZN(new_n538));
  OAI21_X1  g337(.A(KEYINPUT14), .B1(new_n536), .B2(new_n537), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n539), .B1(G29gat), .B2(G36gat), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n535), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n533), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n542), .B1(new_n540), .B2(new_n538), .ZN(new_n543));
  OAI21_X1  g342(.A(KEYINPUT15), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT17), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n535), .A2(new_n538), .A3(new_n540), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT15), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n544), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n540), .A2(new_n538), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(new_n533), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n547), .B1(new_n551), .B2(new_n546), .ZN(new_n552));
  INV_X1    g351(.A(new_n550), .ZN(new_n553));
  AOI21_X1  g352(.A(KEYINPUT15), .B1(new_n553), .B2(new_n535), .ZN(new_n554));
  OAI21_X1  g353(.A(KEYINPUT17), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(G99gat), .A2(G106gat), .ZN(new_n556));
  INV_X1    g355(.A(G85gat), .ZN(new_n557));
  AOI22_X1  g356(.A1(KEYINPUT8), .A2(new_n556), .B1(new_n557), .B2(new_n410), .ZN(new_n558));
  NAND2_X1  g357(.A1(KEYINPUT98), .A2(KEYINPUT7), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n559), .B1(new_n557), .B2(new_n410), .ZN(new_n560));
  NAND4_X1  g359(.A1(KEYINPUT98), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n558), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(G99gat), .B(G106gat), .Z(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n549), .A2(new_n555), .A3(new_n564), .ZN(new_n565));
  AND2_X1   g364(.A1(new_n562), .A2(new_n563), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n562), .A2(new_n563), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n544), .A2(new_n568), .A3(new_n548), .ZN(new_n569));
  NAND3_X1  g368(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n565), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(KEYINPUT99), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT99), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n565), .A2(new_n573), .A3(new_n569), .A4(new_n570), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n572), .A2(new_n202), .A3(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n202), .B1(new_n572), .B2(new_n574), .ZN(new_n577));
  NOR3_X1   g376(.A1(new_n576), .A2(new_n577), .A3(new_n382), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n572), .A2(new_n574), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(G190gat), .ZN(new_n580));
  AOI21_X1  g379(.A(G218gat), .B1(new_n580), .B2(new_n575), .ZN(new_n581));
  OAI21_X1  g380(.A(KEYINPUT100), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(KEYINPUT97), .B(G134gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(G162gat), .ZN(new_n584));
  AOI21_X1  g383(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n382), .B1(new_n576), .B2(new_n577), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n580), .A2(G218gat), .A3(new_n575), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT100), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n582), .A2(new_n587), .A3(new_n591), .ZN(new_n592));
  OAI211_X1 g391(.A(KEYINPUT100), .B(new_n586), .C1(new_n578), .C2(new_n581), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n532), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n518), .A2(new_n568), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n564), .A2(new_n517), .A3(new_n516), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(G230gat), .A2(G233gat), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n602), .B(KEYINPUT102), .Z(new_n603));
  INV_X1    g402(.A(KEYINPUT10), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n597), .A2(new_n598), .A3(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT101), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n518), .A2(new_n568), .A3(KEYINPUT10), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n597), .A2(new_n598), .A3(KEYINPUT101), .A4(new_n604), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(new_n600), .ZN(new_n611));
  XNOR2_X1  g410(.A(G120gat), .B(G148gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT103), .ZN(new_n613));
  INV_X1    g412(.A(G176gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(new_n376), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n603), .A2(new_n611), .A3(new_n617), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n611), .A2(new_n602), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n616), .B(KEYINPUT104), .Z(new_n620));
  OAI21_X1  g419(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT105), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n618), .B(KEYINPUT105), .C1(new_n619), .C2(new_n620), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n596), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n510), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n549), .A2(new_n555), .A3(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n510), .A2(new_n544), .A3(new_n548), .ZN(new_n630));
  NAND2_X1  g429(.A1(G229gat), .A2(G233gat), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT18), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n635));
  XNOR2_X1  g434(.A(G113gat), .B(G141gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G169gat), .B(G197gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n639), .B(KEYINPUT12), .Z(new_n640));
  XNOR2_X1  g439(.A(new_n631), .B(KEYINPUT13), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n630), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n510), .B1(new_n544), .B2(new_n548), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n642), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n629), .A2(KEYINPUT18), .A3(new_n630), .A4(new_n631), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n634), .A2(new_n640), .A3(new_n645), .A4(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(KEYINPUT92), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n646), .A2(new_n645), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT92), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n650), .A2(new_n651), .A3(new_n640), .A4(new_n634), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n649), .A2(KEYINPUT91), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT91), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n646), .A2(new_n645), .A3(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n654), .A2(new_n634), .A3(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n640), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n653), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT93), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n653), .A2(new_n659), .A3(KEYINPUT93), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n500), .A2(new_n627), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n354), .A2(new_n358), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g468(.A1(new_n665), .A2(new_n487), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  OR2_X1    g470(.A1(new_n671), .A2(KEYINPUT106), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n508), .A2(KEYINPUT42), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n671), .A2(KEYINPUT106), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(KEYINPUT16), .B(G8gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(KEYINPUT107), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n671), .A2(KEYINPUT42), .A3(new_n677), .ZN(new_n678));
  OAI211_X1 g477(.A(new_n675), .B(new_n678), .C1(KEYINPUT42), .C2(new_n677), .ZN(G1325gat));
  NAND2_X1  g478(.A1(new_n491), .A2(new_n492), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(G15gat), .B1(new_n665), .B2(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n302), .A2(new_n307), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n683), .A2(KEYINPUT108), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n683), .A2(KEYINPUT108), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(G15gat), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n688), .B(KEYINPUT109), .Z(new_n689));
  AOI21_X1  g488(.A(new_n682), .B1(new_n689), .B2(new_n665), .ZN(G1326gat));
  INV_X1    g489(.A(new_n445), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n665), .A2(KEYINPUT110), .A3(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT110), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n489), .A2(new_n447), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n497), .A2(new_n499), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n532), .A2(new_n595), .A3(new_n625), .ZN(new_n697));
  INV_X1    g496(.A(new_n664), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n693), .B1(new_n699), .B2(new_n445), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n692), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(KEYINPUT43), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT43), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n692), .A2(new_n700), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(G22gat), .ZN(G1327gat));
  NOR2_X1   g505(.A1(new_n531), .A2(new_n625), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NOR4_X1   g507(.A1(new_n500), .A2(new_n594), .A3(new_n664), .A4(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n709), .A2(new_n536), .A3(new_n667), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT45), .ZN(new_n711));
  OAI21_X1  g510(.A(KEYINPUT44), .B1(new_n500), .B2(new_n594), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n713));
  INV_X1    g512(.A(new_n414), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n411), .B1(new_n452), .B2(new_n453), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(KEYINPUT86), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n716), .A2(new_n455), .A3(new_n454), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n714), .B1(new_n717), .B2(KEYINPUT38), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n691), .B1(new_n718), .B2(new_n471), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n488), .A2(new_n486), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n446), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n491), .A2(new_n492), .A3(new_n445), .A4(new_n495), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n722), .A2(KEYINPUT35), .ZN(new_n723));
  AOI22_X1  g522(.A1(new_n723), .A2(new_n496), .B1(KEYINPUT35), .B2(new_n498), .ZN(new_n724));
  OAI211_X1 g523(.A(new_n713), .B(new_n595), .C1(new_n721), .C2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n712), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  AND3_X1   g526(.A1(new_n653), .A2(new_n659), .A3(KEYINPUT111), .ZN(new_n728));
  AOI21_X1  g527(.A(KEYINPUT111), .B1(new_n653), .B2(new_n659), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR4_X1   g529(.A1(new_n727), .A2(new_n666), .A3(new_n730), .A4(new_n708), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n711), .B1(new_n536), .B2(new_n731), .ZN(G1328gat));
  NAND3_X1  g531(.A1(new_n709), .A2(new_n537), .A3(new_n487), .ZN(new_n733));
  XOR2_X1   g532(.A(new_n733), .B(KEYINPUT46), .Z(new_n734));
  NOR4_X1   g533(.A1(new_n727), .A2(new_n495), .A3(new_n730), .A4(new_n708), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n734), .B1(new_n537), .B2(new_n735), .ZN(G1329gat));
  INV_X1    g535(.A(G43gat), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n709), .A2(new_n737), .A3(new_n681), .ZN(new_n738));
  INV_X1    g537(.A(new_n730), .ZN(new_n739));
  AND4_X1   g538(.A1(new_n683), .A2(new_n726), .A3(new_n739), .A4(new_n707), .ZN(new_n740));
  OAI211_X1 g539(.A(KEYINPUT47), .B(new_n738), .C1(new_n740), .C2(new_n737), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n726), .A2(new_n687), .A3(new_n739), .A4(new_n707), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(G43gat), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n743), .A2(new_n738), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n741), .B1(new_n744), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g544(.A1(new_n726), .A2(new_n691), .A3(new_n739), .A4(new_n707), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(G50gat), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT112), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT48), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n709), .A2(new_n435), .A3(new_n691), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n747), .B(new_n750), .C1(new_n748), .C2(KEYINPUT48), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(G1331gat));
  NOR2_X1   g553(.A1(new_n739), .A2(new_n626), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n696), .A2(new_n596), .A3(new_n755), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n756), .A2(new_n666), .ZN(new_n757));
  XOR2_X1   g556(.A(new_n757), .B(G57gat), .Z(G1332gat));
  NOR2_X1   g557(.A1(new_n756), .A2(new_n495), .ZN(new_n759));
  NOR2_X1   g558(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n760));
  AND2_X1   g559(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n762), .B1(new_n759), .B2(new_n760), .ZN(G1333gat));
  OAI21_X1  g562(.A(G71gat), .B1(new_n756), .B2(new_n686), .ZN(new_n764));
  OR2_X1    g563(.A1(new_n680), .A2(G71gat), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n764), .B1(new_n756), .B2(new_n765), .ZN(new_n766));
  XOR2_X1   g565(.A(new_n766), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g566(.A1(new_n756), .A2(new_n445), .ZN(new_n768));
  XOR2_X1   g567(.A(new_n768), .B(G78gat), .Z(G1335gat));
  INV_X1    g568(.A(KEYINPUT51), .ZN(new_n770));
  OAI211_X1 g569(.A(new_n595), .B(new_n730), .C1(new_n721), .C2(new_n724), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n770), .B1(new_n771), .B2(new_n531), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n594), .B1(new_n694), .B2(new_n695), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n773), .A2(KEYINPUT51), .A3(new_n532), .A4(new_n730), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n626), .A2(new_n666), .A3(G85gat), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(KEYINPUT113), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n726), .A2(new_n532), .A3(new_n755), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n779), .A2(new_n667), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n778), .B1(new_n780), .B2(new_n557), .ZN(G1336gat));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n782), .A2(KEYINPUT114), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n775), .A2(new_n625), .A3(new_n487), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n410), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n495), .A2(new_n410), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n726), .A2(new_n532), .A3(new_n755), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n782), .A2(KEYINPUT114), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n784), .B1(new_n786), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n626), .B1(new_n772), .B2(new_n774), .ZN(new_n793));
  AOI21_X1  g592(.A(G92gat), .B1(new_n793), .B2(new_n487), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n794), .A2(new_n783), .A3(new_n790), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n792), .A2(new_n795), .ZN(G1337gat));
  AOI21_X1  g595(.A(G99gat), .B1(new_n793), .B2(new_n681), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n686), .A2(new_n295), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n797), .B1(new_n779), .B2(new_n798), .ZN(G1338gat));
  NAND4_X1  g598(.A1(new_n726), .A2(new_n532), .A3(new_n691), .A4(new_n755), .ZN(new_n800));
  XNOR2_X1  g599(.A(KEYINPUT115), .B(G106gat), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n445), .A2(G106gat), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n775), .A2(new_n625), .A3(new_n803), .ZN(new_n804));
  AOI211_X1 g603(.A(KEYINPUT116), .B(KEYINPUT53), .C1(new_n802), .C2(new_n804), .ZN(new_n805));
  OR2_X1    g604(.A1(KEYINPUT116), .A2(KEYINPUT53), .ZN(new_n806));
  NAND2_X1  g605(.A1(KEYINPUT116), .A2(KEYINPUT53), .ZN(new_n807));
  AND4_X1   g606(.A1(new_n806), .A2(new_n802), .A3(new_n807), .A4(new_n804), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n805), .A2(new_n808), .ZN(G1339gat));
  NOR2_X1   g608(.A1(new_n487), .A2(new_n666), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n607), .A2(new_n601), .A3(new_n608), .A4(new_n609), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n611), .A2(KEYINPUT54), .A3(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT54), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n610), .A2(new_n815), .A3(new_n600), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n616), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n814), .A2(new_n817), .A3(KEYINPUT55), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n816), .A2(new_n616), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n819), .B1(new_n820), .B2(new_n813), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n618), .B1(new_n818), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n629), .A2(new_n630), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n823), .A2(G229gat), .A3(G233gat), .ZN(new_n824));
  OR3_X1    g623(.A1(new_n643), .A2(new_n644), .A3(new_n642), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n639), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AOI211_X1 g625(.A(KEYINPUT117), .B(new_n826), .C1(new_n648), .C2(new_n652), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n822), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n826), .B1(new_n648), .B2(new_n652), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(KEYINPUT117), .ZN(new_n831));
  AND4_X1   g630(.A1(new_n593), .A2(new_n828), .A3(new_n592), .A4(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(new_n618), .ZN(new_n833));
  OAI21_X1  g632(.A(KEYINPUT55), .B1(new_n814), .B2(new_n817), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n820), .A2(new_n819), .A3(new_n813), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n836), .B1(new_n728), .B2(new_n729), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n625), .A2(new_n829), .ZN(new_n838));
  AOI22_X1  g637(.A1(new_n837), .A2(new_n838), .B1(new_n592), .B2(new_n593), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n532), .B1(new_n832), .B2(new_n839), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n531), .A2(new_n594), .A3(new_n626), .A4(new_n730), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n811), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n493), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(G113gat), .B1(new_n846), .B2(new_n664), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n301), .A2(new_n445), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n842), .A2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(new_n245), .A3(new_n739), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n847), .A2(new_n851), .ZN(G1340gat));
  OAI21_X1  g651(.A(G120gat), .B1(new_n846), .B2(new_n626), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n850), .A2(new_n243), .A3(new_n625), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(G1341gat));
  NAND2_X1  g654(.A1(new_n850), .A2(new_n531), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n254), .A2(new_n255), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n532), .A2(new_n857), .ZN(new_n858));
  AOI22_X1  g657(.A1(new_n856), .A2(new_n857), .B1(new_n845), .B2(new_n858), .ZN(G1342gat));
  AOI21_X1  g658(.A(new_n250), .B1(new_n845), .B2(new_n595), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(KEYINPUT118), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n860), .A2(KEYINPUT118), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n849), .B1(new_n252), .B2(new_n251), .ZN(new_n864));
  AOI21_X1  g663(.A(KEYINPUT56), .B1(new_n864), .B2(new_n595), .ZN(new_n865));
  AND3_X1   g664(.A1(new_n864), .A2(KEYINPUT56), .A3(new_n595), .ZN(new_n866));
  OAI22_X1  g665(.A1(new_n862), .A2(new_n863), .B1(new_n865), .B2(new_n866), .ZN(G1343gat));
  INV_X1    g666(.A(KEYINPUT58), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n662), .A2(new_n663), .A3(new_n836), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n838), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n594), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n828), .A2(new_n592), .A3(new_n593), .A4(new_n831), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n531), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n841), .ZN(new_n874));
  OAI211_X1 g673(.A(KEYINPUT57), .B(new_n691), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n445), .B1(new_n840), .B2(new_n841), .ZN(new_n876));
  XNOR2_X1  g675(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n683), .A2(new_n811), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n878), .A2(new_n739), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(G141gat), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n842), .A2(new_n691), .A3(new_n698), .A4(new_n686), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n882), .A2(G141gat), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n868), .B1(new_n881), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n868), .B1(new_n882), .B2(G141gat), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n878), .A2(new_n698), .A3(new_n879), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n886), .B1(G141gat), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(KEYINPUT120), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n887), .A2(G141gat), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n890), .A2(new_n868), .A3(new_n884), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT120), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n883), .B1(new_n880), .B2(G141gat), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n891), .B(new_n892), .C1(new_n868), .C2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n889), .A2(new_n894), .ZN(G1344gat));
  NOR3_X1   g694(.A1(new_n843), .A2(new_n445), .A3(new_n687), .ZN(new_n896));
  INV_X1    g695(.A(G148gat), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n896), .A2(new_n897), .A3(new_n625), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT59), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n697), .A2(new_n664), .ZN(new_n900));
  INV_X1    g699(.A(new_n873), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n691), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT57), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n876), .A2(new_n877), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n626), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n879), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n899), .B1(new_n908), .B2(G148gat), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n878), .A2(new_n879), .ZN(new_n910));
  AOI211_X1 g709(.A(KEYINPUT59), .B(new_n897), .C1(new_n910), .C2(new_n625), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n898), .B1(new_n909), .B2(new_n911), .ZN(G1345gat));
  AOI21_X1  g711(.A(G155gat), .B1(new_n896), .B2(new_n531), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n531), .A2(G155gat), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n913), .B1(new_n910), .B2(new_n914), .ZN(G1346gat));
  AOI21_X1  g714(.A(G162gat), .B1(new_n896), .B2(new_n595), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n595), .A2(G162gat), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n916), .B1(new_n910), .B2(new_n917), .ZN(G1347gat));
  NAND2_X1  g717(.A1(new_n487), .A2(new_n666), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT111), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n660), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n653), .A2(new_n659), .A3(KEYINPUT111), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n822), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n830), .B1(new_n623), .B2(new_n624), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n594), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n531), .B1(new_n926), .B2(new_n872), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n493), .B(new_n920), .C1(new_n927), .C2(new_n874), .ZN(new_n928));
  OAI21_X1  g727(.A(G169gat), .B1(new_n928), .B2(new_n664), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n919), .B1(new_n840), .B2(new_n841), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(new_n848), .ZN(new_n931));
  OR2_X1    g730(.A1(new_n730), .A2(G169gat), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(G1348gat));
  NOR3_X1   g732(.A1(new_n928), .A2(new_n614), .A3(new_n626), .ZN(new_n934));
  INV_X1    g733(.A(new_n931), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(new_n625), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n934), .B1(new_n936), .B2(new_n614), .ZN(G1349gat));
  OAI21_X1  g736(.A(KEYINPUT121), .B1(new_n928), .B2(new_n532), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT121), .ZN(new_n939));
  NAND4_X1  g738(.A1(new_n930), .A2(new_n939), .A3(new_n531), .A4(new_n493), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n938), .A2(new_n940), .A3(G183gat), .ZN(new_n941));
  OR2_X1    g740(.A1(new_n203), .A2(new_n204), .ZN(new_n942));
  NAND4_X1  g741(.A1(new_n930), .A2(new_n531), .A3(new_n942), .A4(new_n848), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(KEYINPUT122), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT122), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n941), .A2(new_n946), .A3(new_n943), .ZN(new_n947));
  NAND4_X1  g746(.A1(new_n945), .A2(KEYINPUT123), .A3(KEYINPUT60), .A4(new_n947), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n941), .A2(new_n946), .A3(new_n943), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n946), .B1(new_n941), .B2(new_n943), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT60), .ZN(new_n951));
  NOR3_X1   g750(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n941), .A2(new_n951), .A3(new_n943), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n953), .A2(KEYINPUT123), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n948), .B1(new_n952), .B2(new_n954), .ZN(G1350gat));
  OAI21_X1  g754(.A(G190gat), .B1(new_n928), .B2(new_n594), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n956), .B(KEYINPUT61), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n935), .A2(new_n202), .A3(new_n595), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(G1351gat));
  NOR3_X1   g758(.A1(new_n684), .A2(new_n685), .A3(new_n919), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n876), .A2(new_n960), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n962), .A2(new_n371), .A3(new_n739), .ZN(new_n963));
  AOI21_X1  g762(.A(KEYINPUT57), .B1(new_n902), .B2(new_n691), .ZN(new_n964));
  INV_X1    g763(.A(new_n906), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g765(.A(new_n960), .ZN(new_n967));
  NOR3_X1   g766(.A1(new_n966), .A2(new_n664), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n963), .B1(new_n968), .B2(new_n371), .ZN(G1352gat));
  AOI21_X1  g768(.A(new_n376), .B1(new_n907), .B2(new_n960), .ZN(new_n970));
  NAND4_X1  g769(.A1(new_n876), .A2(new_n376), .A3(new_n625), .A4(new_n960), .ZN(new_n971));
  XNOR2_X1  g770(.A(new_n971), .B(KEYINPUT62), .ZN(new_n972));
  OAI21_X1  g771(.A(KEYINPUT124), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT124), .ZN(new_n974));
  INV_X1    g773(.A(new_n972), .ZN(new_n975));
  NOR3_X1   g774(.A1(new_n966), .A2(new_n626), .A3(new_n967), .ZN(new_n976));
  OAI211_X1 g775(.A(new_n974), .B(new_n975), .C1(new_n976), .C2(new_n376), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n973), .A2(new_n977), .ZN(G1353gat));
  NAND3_X1  g777(.A1(new_n962), .A2(new_n389), .A3(new_n531), .ZN(new_n979));
  OAI211_X1 g778(.A(new_n531), .B(new_n960), .C1(new_n964), .C2(new_n965), .ZN(new_n980));
  AND3_X1   g779(.A1(new_n980), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n981));
  AOI21_X1  g780(.A(KEYINPUT63), .B1(new_n980), .B2(G211gat), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n979), .B1(new_n981), .B2(new_n982), .ZN(G1354gat));
  INV_X1    g782(.A(KEYINPUT126), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n984), .B1(new_n966), .B2(new_n967), .ZN(new_n985));
  AND2_X1   g784(.A1(new_n595), .A2(new_n369), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n986), .A2(KEYINPUT127), .ZN(new_n987));
  OAI211_X1 g786(.A(KEYINPUT126), .B(new_n960), .C1(new_n964), .C2(new_n965), .ZN(new_n988));
  OR2_X1    g787(.A1(new_n986), .A2(KEYINPUT127), .ZN(new_n989));
  NAND4_X1  g788(.A1(new_n985), .A2(new_n987), .A3(new_n988), .A4(new_n989), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n382), .B1(new_n961), .B2(new_n594), .ZN(new_n991));
  XOR2_X1   g790(.A(new_n991), .B(KEYINPUT125), .Z(new_n992));
  AND2_X1   g791(.A1(new_n990), .A2(new_n992), .ZN(G1355gat));
endmodule


