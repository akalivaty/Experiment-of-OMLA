

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X2 U552 ( .A(KEYINPUT64), .B(n540), .ZN(n582) );
  NAND2_X1 U553 ( .A1(n722), .A2(n612), .ZN(n670) );
  NOR2_X1 U554 ( .A1(G543), .A2(G651), .ZN(n807) );
  XNOR2_X1 U555 ( .A(n775), .B(KEYINPUT40), .ZN(n776) );
  XNOR2_X1 U556 ( .A(n777), .B(n776), .ZN(G329) );
  NOR2_X1 U557 ( .A1(n532), .A2(n531), .ZN(G160) );
  INV_X1 U558 ( .A(KEYINPUT67), .ZN(n520) );
  NAND2_X1 U559 ( .A1(G2105), .A2(G2104), .ZN(n518) );
  XOR2_X1 U560 ( .A(KEYINPUT66), .B(n518), .Z(n729) );
  NAND2_X1 U561 ( .A1(G113), .A2(n729), .ZN(n519) );
  XNOR2_X1 U562 ( .A(n520), .B(n519), .ZN(n523) );
  NOR2_X1 U563 ( .A1(G2105), .A2(G2104), .ZN(n521) );
  XOR2_X2 U564 ( .A(KEYINPUT17), .B(n521), .Z(n895) );
  NAND2_X1 U565 ( .A1(n895), .A2(G137), .ZN(n522) );
  NAND2_X1 U566 ( .A1(n523), .A2(n522), .ZN(n525) );
  INV_X1 U567 ( .A(KEYINPUT68), .ZN(n524) );
  XNOR2_X1 U568 ( .A(n525), .B(n524), .ZN(n528) );
  INV_X1 U569 ( .A(G2104), .ZN(n529) );
  NAND2_X1 U570 ( .A1(n529), .A2(G2105), .ZN(n526) );
  XNOR2_X1 U571 ( .A(n526), .B(KEYINPUT65), .ZN(n890) );
  NAND2_X1 U572 ( .A1(n890), .A2(G125), .ZN(n527) );
  NAND2_X1 U573 ( .A1(n528), .A2(n527), .ZN(n532) );
  NOR2_X1 U574 ( .A1(G2105), .A2(n529), .ZN(n894) );
  NAND2_X1 U575 ( .A1(G101), .A2(n894), .ZN(n530) );
  XNOR2_X1 U576 ( .A(KEYINPUT23), .B(n530), .ZN(n531) );
  NAND2_X1 U577 ( .A1(G102), .A2(n894), .ZN(n534) );
  NAND2_X1 U578 ( .A1(G138), .A2(n895), .ZN(n533) );
  NAND2_X1 U579 ( .A1(n534), .A2(n533), .ZN(n538) );
  NAND2_X1 U580 ( .A1(G126), .A2(n890), .ZN(n536) );
  NAND2_X1 U581 ( .A1(G114), .A2(n729), .ZN(n535) );
  NAND2_X1 U582 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U583 ( .A1(n538), .A2(n537), .ZN(G164) );
  INV_X1 U584 ( .A(G651), .ZN(n543) );
  NOR2_X1 U585 ( .A1(G543), .A2(n543), .ZN(n539) );
  XOR2_X1 U586 ( .A(KEYINPUT1), .B(n539), .Z(n804) );
  NAND2_X1 U587 ( .A1(n804), .A2(G65), .ZN(n542) );
  XOR2_X1 U588 ( .A(KEYINPUT0), .B(G543), .Z(n586) );
  NOR2_X1 U589 ( .A1(n586), .A2(G651), .ZN(n540) );
  NAND2_X1 U590 ( .A1(G53), .A2(n582), .ZN(n541) );
  NAND2_X1 U591 ( .A1(n542), .A2(n541), .ZN(n546) );
  NOR2_X1 U592 ( .A1(n586), .A2(n543), .ZN(n808) );
  NAND2_X1 U593 ( .A1(G78), .A2(n808), .ZN(n544) );
  XNOR2_X1 U594 ( .A(KEYINPUT71), .B(n544), .ZN(n545) );
  NOR2_X1 U595 ( .A1(n546), .A2(n545), .ZN(n548) );
  NAND2_X1 U596 ( .A1(n807), .A2(G91), .ZN(n547) );
  NAND2_X1 U597 ( .A1(n548), .A2(n547), .ZN(G299) );
  NAND2_X1 U598 ( .A1(G52), .A2(n582), .ZN(n549) );
  XNOR2_X1 U599 ( .A(KEYINPUT69), .B(n549), .ZN(n557) );
  NAND2_X1 U600 ( .A1(G90), .A2(n807), .ZN(n551) );
  NAND2_X1 U601 ( .A1(G77), .A2(n808), .ZN(n550) );
  NAND2_X1 U602 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U603 ( .A(n552), .B(KEYINPUT9), .ZN(n553) );
  XNOR2_X1 U604 ( .A(n553), .B(KEYINPUT70), .ZN(n555) );
  NAND2_X1 U605 ( .A1(n804), .A2(G64), .ZN(n554) );
  NAND2_X1 U606 ( .A1(n555), .A2(n554), .ZN(n556) );
  NOR2_X1 U607 ( .A1(n557), .A2(n556), .ZN(G171) );
  INV_X1 U608 ( .A(G171), .ZN(G301) );
  NAND2_X1 U609 ( .A1(G51), .A2(n582), .ZN(n558) );
  XOR2_X1 U610 ( .A(KEYINPUT77), .B(n558), .Z(n560) );
  NAND2_X1 U611 ( .A1(n804), .A2(G63), .ZN(n559) );
  NAND2_X1 U612 ( .A1(n560), .A2(n559), .ZN(n562) );
  XOR2_X1 U613 ( .A(KEYINPUT6), .B(KEYINPUT78), .Z(n561) );
  XOR2_X1 U614 ( .A(n562), .B(n561), .Z(n570) );
  NAND2_X1 U615 ( .A1(n808), .A2(G76), .ZN(n563) );
  XOR2_X1 U616 ( .A(KEYINPUT76), .B(n563), .Z(n567) );
  NAND2_X1 U617 ( .A1(G89), .A2(n807), .ZN(n564) );
  XNOR2_X1 U618 ( .A(n564), .B(KEYINPUT75), .ZN(n565) );
  XNOR2_X1 U619 ( .A(n565), .B(KEYINPUT4), .ZN(n566) );
  NOR2_X1 U620 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U621 ( .A(KEYINPUT5), .B(n568), .ZN(n569) );
  NOR2_X1 U622 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U623 ( .A(n571), .B(KEYINPUT7), .ZN(n572) );
  XNOR2_X1 U624 ( .A(n572), .B(KEYINPUT79), .ZN(G168) );
  NAND2_X1 U625 ( .A1(G88), .A2(n807), .ZN(n574) );
  NAND2_X1 U626 ( .A1(G75), .A2(n808), .ZN(n573) );
  NAND2_X1 U627 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U628 ( .A(KEYINPUT88), .B(n575), .ZN(n580) );
  NAND2_X1 U629 ( .A1(n804), .A2(G62), .ZN(n577) );
  NAND2_X1 U630 ( .A1(G50), .A2(n582), .ZN(n576) );
  NAND2_X1 U631 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U632 ( .A(KEYINPUT87), .B(n578), .Z(n579) );
  NOR2_X1 U633 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U634 ( .A(KEYINPUT89), .B(n581), .ZN(G303) );
  XOR2_X1 U635 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U636 ( .A(G303), .ZN(G166) );
  NAND2_X1 U637 ( .A1(G651), .A2(G74), .ZN(n584) );
  NAND2_X1 U638 ( .A1(G49), .A2(n582), .ZN(n583) );
  NAND2_X1 U639 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U640 ( .A(KEYINPUT84), .B(n585), .Z(n588) );
  NAND2_X1 U641 ( .A1(n586), .A2(G87), .ZN(n587) );
  NAND2_X1 U642 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U643 ( .A1(n589), .A2(n804), .ZN(n590) );
  XNOR2_X1 U644 ( .A(n590), .B(KEYINPUT85), .ZN(G288) );
  XOR2_X1 U645 ( .A(KEYINPUT86), .B(KEYINPUT2), .Z(n592) );
  NAND2_X1 U646 ( .A1(G73), .A2(n808), .ZN(n591) );
  XNOR2_X1 U647 ( .A(n592), .B(n591), .ZN(n596) );
  NAND2_X1 U648 ( .A1(n804), .A2(G61), .ZN(n594) );
  NAND2_X1 U649 ( .A1(G48), .A2(n582), .ZN(n593) );
  NAND2_X1 U650 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U651 ( .A1(n596), .A2(n595), .ZN(n598) );
  NAND2_X1 U652 ( .A1(n807), .A2(G86), .ZN(n597) );
  NAND2_X1 U653 ( .A1(n598), .A2(n597), .ZN(G305) );
  AND2_X1 U654 ( .A1(n804), .A2(G60), .ZN(n602) );
  NAND2_X1 U655 ( .A1(n807), .A2(G85), .ZN(n600) );
  NAND2_X1 U656 ( .A1(G47), .A2(n582), .ZN(n599) );
  NAND2_X1 U657 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U658 ( .A1(n602), .A2(n601), .ZN(n604) );
  NAND2_X1 U659 ( .A1(n808), .A2(G72), .ZN(n603) );
  NAND2_X1 U660 ( .A1(n604), .A2(n603), .ZN(G290) );
  NAND2_X1 U661 ( .A1(G92), .A2(n807), .ZN(n606) );
  NAND2_X1 U662 ( .A1(G79), .A2(n808), .ZN(n605) );
  NAND2_X1 U663 ( .A1(n606), .A2(n605), .ZN(n610) );
  NAND2_X1 U664 ( .A1(n804), .A2(G66), .ZN(n608) );
  NAND2_X1 U665 ( .A1(G54), .A2(n582), .ZN(n607) );
  NAND2_X1 U666 ( .A1(n608), .A2(n607), .ZN(n609) );
  NOR2_X1 U667 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U668 ( .A(n611), .B(KEYINPUT15), .ZN(n928) );
  NOR2_X1 U669 ( .A1(G164), .A2(G1384), .ZN(n722) );
  NAND2_X1 U670 ( .A1(G160), .A2(G40), .ZN(n721) );
  INV_X1 U671 ( .A(n721), .ZN(n612) );
  NAND2_X1 U672 ( .A1(G1348), .A2(n670), .ZN(n614) );
  INV_X1 U673 ( .A(n670), .ZN(n649) );
  NAND2_X1 U674 ( .A1(G2067), .A2(n649), .ZN(n613) );
  NAND2_X1 U675 ( .A1(n614), .A2(n613), .ZN(n632) );
  NOR2_X1 U676 ( .A1(n928), .A2(n632), .ZN(n631) );
  NAND2_X1 U677 ( .A1(n582), .A2(G43), .ZN(n624) );
  NAND2_X1 U678 ( .A1(n804), .A2(G56), .ZN(n615) );
  XNOR2_X1 U679 ( .A(KEYINPUT14), .B(n615), .ZN(n621) );
  NAND2_X1 U680 ( .A1(n807), .A2(G81), .ZN(n616) );
  XNOR2_X1 U681 ( .A(n616), .B(KEYINPUT12), .ZN(n618) );
  NAND2_X1 U682 ( .A1(G68), .A2(n808), .ZN(n617) );
  NAND2_X1 U683 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U684 ( .A(KEYINPUT13), .B(n619), .ZN(n620) );
  NAND2_X1 U685 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U686 ( .A(KEYINPUT73), .B(n622), .ZN(n623) );
  NAND2_X1 U687 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U688 ( .A(n625), .B(KEYINPUT74), .ZN(n939) );
  NAND2_X1 U689 ( .A1(n649), .A2(G1996), .ZN(n626) );
  XNOR2_X1 U690 ( .A(n626), .B(KEYINPUT26), .ZN(n628) );
  NAND2_X1 U691 ( .A1(n670), .A2(G1341), .ZN(n627) );
  NAND2_X1 U692 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U693 ( .A1(n939), .A2(n629), .ZN(n630) );
  NOR2_X1 U694 ( .A1(n631), .A2(n630), .ZN(n634) );
  AND2_X1 U695 ( .A1(n928), .A2(n632), .ZN(n633) );
  NOR2_X1 U696 ( .A1(n634), .A2(n633), .ZN(n641) );
  INV_X1 U697 ( .A(n670), .ZN(n635) );
  NAND2_X1 U698 ( .A1(n635), .A2(G2072), .ZN(n636) );
  XOR2_X1 U699 ( .A(n636), .B(KEYINPUT27), .Z(n638) );
  NAND2_X1 U700 ( .A1(G1956), .A2(n670), .ZN(n637) );
  NAND2_X1 U701 ( .A1(n638), .A2(n637), .ZN(n642) );
  NOR2_X1 U702 ( .A1(G299), .A2(n642), .ZN(n639) );
  XOR2_X1 U703 ( .A(KEYINPUT99), .B(n639), .Z(n640) );
  NOR2_X1 U704 ( .A1(n641), .A2(n640), .ZN(n645) );
  NAND2_X1 U705 ( .A1(G299), .A2(n642), .ZN(n643) );
  XOR2_X1 U706 ( .A(KEYINPUT28), .B(n643), .Z(n644) );
  NOR2_X1 U707 ( .A1(n645), .A2(n644), .ZN(n648) );
  XNOR2_X1 U708 ( .A(KEYINPUT100), .B(KEYINPUT101), .ZN(n646) );
  XNOR2_X1 U709 ( .A(n646), .B(KEYINPUT29), .ZN(n647) );
  XNOR2_X1 U710 ( .A(n648), .B(n647), .ZN(n678) );
  XOR2_X1 U711 ( .A(KEYINPUT25), .B(G2078), .Z(n988) );
  NOR2_X1 U712 ( .A1(n988), .A2(n670), .ZN(n651) );
  NOR2_X1 U713 ( .A1(n649), .A2(G1961), .ZN(n650) );
  NOR2_X1 U714 ( .A1(n651), .A2(n650), .ZN(n657) );
  NOR2_X1 U715 ( .A1(G301), .A2(n657), .ZN(n676) );
  INV_X1 U716 ( .A(G8), .ZN(n652) );
  NOR2_X1 U717 ( .A1(n652), .A2(G1966), .ZN(n653) );
  AND2_X1 U718 ( .A1(n670), .A2(n653), .ZN(n659) );
  NOR2_X1 U719 ( .A1(G2084), .A2(n670), .ZN(n658) );
  AND2_X1 U720 ( .A1(G8), .A2(n658), .ZN(n654) );
  OR2_X1 U721 ( .A1(n659), .A2(n654), .ZN(n656) );
  OR2_X1 U722 ( .A1(n676), .A2(n656), .ZN(n655) );
  NOR2_X1 U723 ( .A1(n678), .A2(n655), .ZN(n668) );
  INV_X1 U724 ( .A(n656), .ZN(n666) );
  AND2_X1 U725 ( .A1(G301), .A2(n657), .ZN(n664) );
  NOR2_X1 U726 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U727 ( .A1(G8), .A2(n660), .ZN(n661) );
  XNOR2_X1 U728 ( .A(KEYINPUT30), .B(n661), .ZN(n662) );
  NOR2_X1 U729 ( .A1(G168), .A2(n662), .ZN(n663) );
  NOR2_X1 U730 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U731 ( .A(n665), .B(KEYINPUT31), .ZN(n681) );
  AND2_X1 U732 ( .A1(n666), .A2(n681), .ZN(n667) );
  NOR2_X1 U733 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U734 ( .A(n669), .B(KEYINPUT102), .ZN(n700) );
  NAND2_X1 U735 ( .A1(G8), .A2(n670), .ZN(n714) );
  NOR2_X1 U736 ( .A1(G1971), .A2(n714), .ZN(n672) );
  NOR2_X1 U737 ( .A1(G2090), .A2(n670), .ZN(n671) );
  NOR2_X1 U738 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U739 ( .A1(n673), .A2(G303), .ZN(n674) );
  NOR2_X1 U740 ( .A1(n652), .A2(n674), .ZN(n680) );
  AND2_X1 U741 ( .A1(G286), .A2(G8), .ZN(n675) );
  NOR2_X1 U742 ( .A1(n680), .A2(n675), .ZN(n679) );
  OR2_X1 U743 ( .A1(n676), .A2(n679), .ZN(n677) );
  NOR2_X1 U744 ( .A1(n678), .A2(n677), .ZN(n685) );
  INV_X1 U745 ( .A(n679), .ZN(n683) );
  OR2_X1 U746 ( .A1(n681), .A2(n680), .ZN(n682) );
  AND2_X1 U747 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U748 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U749 ( .A(n686), .B(KEYINPUT32), .ZN(n697) );
  NAND2_X1 U750 ( .A1(n700), .A2(n697), .ZN(n689) );
  NAND2_X1 U751 ( .A1(G166), .A2(G8), .ZN(n687) );
  OR2_X1 U752 ( .A1(G2090), .A2(n687), .ZN(n688) );
  NAND2_X1 U753 ( .A1(n689), .A2(n688), .ZN(n691) );
  INV_X1 U754 ( .A(KEYINPUT105), .ZN(n690) );
  XNOR2_X1 U755 ( .A(n691), .B(n690), .ZN(n692) );
  NAND2_X1 U756 ( .A1(n692), .A2(n714), .ZN(n720) );
  NAND2_X1 U757 ( .A1(G1976), .A2(G288), .ZN(n937) );
  INV_X1 U758 ( .A(KEYINPUT33), .ZN(n704) );
  NOR2_X1 U759 ( .A1(G1976), .A2(G288), .ZN(n693) );
  XNOR2_X1 U760 ( .A(KEYINPUT103), .B(n693), .ZN(n948) );
  OR2_X1 U761 ( .A1(n714), .A2(n948), .ZN(n694) );
  NOR2_X1 U762 ( .A1(n704), .A2(n694), .ZN(n695) );
  XOR2_X1 U763 ( .A(n695), .B(KEYINPUT104), .Z(n703) );
  NAND2_X1 U764 ( .A1(n937), .A2(n703), .ZN(n696) );
  OR2_X1 U765 ( .A1(n696), .A2(n714), .ZN(n708) );
  INV_X1 U766 ( .A(n708), .ZN(n698) );
  AND2_X1 U767 ( .A1(n698), .A2(n697), .ZN(n702) );
  XNOR2_X1 U768 ( .A(G1981), .B(G305), .ZN(n941) );
  INV_X1 U769 ( .A(n941), .ZN(n699) );
  AND2_X1 U770 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U771 ( .A1(n702), .A2(n701), .ZN(n718) );
  INV_X1 U772 ( .A(n703), .ZN(n705) );
  OR2_X1 U773 ( .A1(n705), .A2(n704), .ZN(n710) );
  OR2_X1 U774 ( .A1(G1971), .A2(G303), .ZN(n706) );
  AND2_X1 U775 ( .A1(n948), .A2(n706), .ZN(n707) );
  OR2_X1 U776 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U777 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U778 ( .A1(n941), .A2(n711), .ZN(n716) );
  NOR2_X1 U779 ( .A1(G1981), .A2(G305), .ZN(n712) );
  XOR2_X1 U780 ( .A(n712), .B(KEYINPUT24), .Z(n713) );
  NOR2_X1 U781 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U782 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U783 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U784 ( .A1(n720), .A2(n719), .ZN(n737) );
  NOR2_X1 U785 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U786 ( .A(KEYINPUT93), .B(n723), .ZN(n772) );
  XOR2_X1 U787 ( .A(G2067), .B(KEYINPUT37), .Z(n760) );
  NAND2_X1 U788 ( .A1(n895), .A2(G140), .ZN(n724) );
  XNOR2_X1 U789 ( .A(n724), .B(KEYINPUT94), .ZN(n726) );
  NAND2_X1 U790 ( .A1(G104), .A2(n894), .ZN(n725) );
  NAND2_X1 U791 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U792 ( .A(KEYINPUT34), .B(n727), .ZN(n734) );
  NAND2_X1 U793 ( .A1(n890), .A2(G128), .ZN(n728) );
  XOR2_X1 U794 ( .A(KEYINPUT95), .B(n728), .Z(n731) );
  BUF_X1 U795 ( .A(n729), .Z(n891) );
  NAND2_X1 U796 ( .A1(G116), .A2(n891), .ZN(n730) );
  NAND2_X1 U797 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U798 ( .A(KEYINPUT35), .B(n732), .Z(n733) );
  NOR2_X1 U799 ( .A1(n734), .A2(n733), .ZN(n735) );
  XOR2_X1 U800 ( .A(KEYINPUT36), .B(n735), .Z(n887) );
  NAND2_X1 U801 ( .A1(n760), .A2(n887), .ZN(n955) );
  NOR2_X1 U802 ( .A1(n772), .A2(n955), .ZN(n768) );
  INV_X1 U803 ( .A(n768), .ZN(n736) );
  NAND2_X1 U804 ( .A1(n737), .A2(n736), .ZN(n758) );
  XNOR2_X1 U805 ( .A(G1986), .B(G290), .ZN(n932) );
  XOR2_X1 U806 ( .A(KEYINPUT38), .B(KEYINPUT98), .Z(n739) );
  NAND2_X1 U807 ( .A1(G105), .A2(n894), .ZN(n738) );
  XNOR2_X1 U808 ( .A(n739), .B(n738), .ZN(n744) );
  NAND2_X1 U809 ( .A1(G129), .A2(n890), .ZN(n741) );
  NAND2_X1 U810 ( .A1(G117), .A2(n891), .ZN(n740) );
  NAND2_X1 U811 ( .A1(n741), .A2(n740), .ZN(n742) );
  XOR2_X1 U812 ( .A(KEYINPUT97), .B(n742), .Z(n743) );
  NOR2_X1 U813 ( .A1(n744), .A2(n743), .ZN(n746) );
  NAND2_X1 U814 ( .A1(n895), .A2(G141), .ZN(n745) );
  NAND2_X1 U815 ( .A1(n746), .A2(n745), .ZN(n881) );
  NAND2_X1 U816 ( .A1(G1996), .A2(n881), .ZN(n755) );
  NAND2_X1 U817 ( .A1(G95), .A2(n894), .ZN(n748) );
  NAND2_X1 U818 ( .A1(G119), .A2(n890), .ZN(n747) );
  NAND2_X1 U819 ( .A1(n748), .A2(n747), .ZN(n751) );
  NAND2_X1 U820 ( .A1(n895), .A2(G131), .ZN(n749) );
  XOR2_X1 U821 ( .A(KEYINPUT96), .B(n749), .Z(n750) );
  NOR2_X1 U822 ( .A1(n751), .A2(n750), .ZN(n753) );
  NAND2_X1 U823 ( .A1(G107), .A2(n891), .ZN(n752) );
  NAND2_X1 U824 ( .A1(n753), .A2(n752), .ZN(n901) );
  NAND2_X1 U825 ( .A1(G1991), .A2(n901), .ZN(n754) );
  NAND2_X1 U826 ( .A1(n755), .A2(n754), .ZN(n956) );
  NOR2_X1 U827 ( .A1(n932), .A2(n956), .ZN(n756) );
  NOR2_X1 U828 ( .A1(n772), .A2(n756), .ZN(n757) );
  NOR2_X1 U829 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U830 ( .A(n759), .B(KEYINPUT106), .ZN(n774) );
  NOR2_X1 U831 ( .A1(n760), .A2(n887), .ZN(n761) );
  XOR2_X1 U832 ( .A(KEYINPUT109), .B(n761), .Z(n966) );
  NOR2_X1 U833 ( .A1(G1996), .A2(n881), .ZN(n762) );
  XOR2_X1 U834 ( .A(KEYINPUT107), .B(n762), .Z(n953) );
  NOR2_X1 U835 ( .A1(G1986), .A2(G290), .ZN(n763) );
  NOR2_X1 U836 ( .A1(G1991), .A2(n901), .ZN(n961) );
  NOR2_X1 U837 ( .A1(n763), .A2(n961), .ZN(n764) );
  NOR2_X1 U838 ( .A1(n956), .A2(n764), .ZN(n765) );
  NOR2_X1 U839 ( .A1(n953), .A2(n765), .ZN(n766) );
  XOR2_X1 U840 ( .A(KEYINPUT39), .B(n766), .Z(n767) );
  NOR2_X1 U841 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U842 ( .A(n769), .B(KEYINPUT108), .ZN(n770) );
  NOR2_X1 U843 ( .A1(n966), .A2(n770), .ZN(n771) );
  NOR2_X1 U844 ( .A1(n772), .A2(n771), .ZN(n773) );
  NOR2_X1 U845 ( .A1(n774), .A2(n773), .ZN(n777) );
  INV_X1 U846 ( .A(KEYINPUT110), .ZN(n775) );
  AND2_X1 U847 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U848 ( .A(G57), .ZN(G237) );
  INV_X1 U849 ( .A(G132), .ZN(G219) );
  NAND2_X1 U850 ( .A1(G7), .A2(G661), .ZN(n778) );
  XNOR2_X1 U851 ( .A(n778), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U852 ( .A(G223), .ZN(n839) );
  NAND2_X1 U853 ( .A1(n839), .A2(G567), .ZN(n779) );
  XOR2_X1 U854 ( .A(KEYINPUT11), .B(n779), .Z(G234) );
  INV_X1 U855 ( .A(G860), .ZN(n785) );
  OR2_X1 U856 ( .A1(n785), .A2(n939), .ZN(G153) );
  NAND2_X1 U857 ( .A1(G868), .A2(G301), .ZN(n781) );
  INV_X1 U858 ( .A(G868), .ZN(n782) );
  NAND2_X1 U859 ( .A1(n928), .A2(n782), .ZN(n780) );
  NAND2_X1 U860 ( .A1(n781), .A2(n780), .ZN(G284) );
  NOR2_X1 U861 ( .A1(G286), .A2(n782), .ZN(n784) );
  NOR2_X1 U862 ( .A1(G868), .A2(G299), .ZN(n783) );
  NOR2_X1 U863 ( .A1(n784), .A2(n783), .ZN(G297) );
  NAND2_X1 U864 ( .A1(n785), .A2(G559), .ZN(n786) );
  INV_X1 U865 ( .A(n928), .ZN(n907) );
  NAND2_X1 U866 ( .A1(n786), .A2(n907), .ZN(n787) );
  XNOR2_X1 U867 ( .A(n787), .B(KEYINPUT16), .ZN(n788) );
  XNOR2_X1 U868 ( .A(KEYINPUT80), .B(n788), .ZN(G148) );
  NOR2_X1 U869 ( .A1(n939), .A2(G868), .ZN(n791) );
  NAND2_X1 U870 ( .A1(n907), .A2(G868), .ZN(n789) );
  NOR2_X1 U871 ( .A1(G559), .A2(n789), .ZN(n790) );
  NOR2_X1 U872 ( .A1(n791), .A2(n790), .ZN(G282) );
  XNOR2_X1 U873 ( .A(G2096), .B(KEYINPUT82), .ZN(n800) );
  NAND2_X1 U874 ( .A1(G123), .A2(n890), .ZN(n792) );
  XNOR2_X1 U875 ( .A(n792), .B(KEYINPUT18), .ZN(n799) );
  NAND2_X1 U876 ( .A1(G99), .A2(n894), .ZN(n794) );
  NAND2_X1 U877 ( .A1(G111), .A2(n891), .ZN(n793) );
  NAND2_X1 U878 ( .A1(n794), .A2(n793), .ZN(n797) );
  NAND2_X1 U879 ( .A1(G135), .A2(n895), .ZN(n795) );
  XNOR2_X1 U880 ( .A(KEYINPUT81), .B(n795), .ZN(n796) );
  NOR2_X1 U881 ( .A1(n797), .A2(n796), .ZN(n798) );
  NAND2_X1 U882 ( .A1(n799), .A2(n798), .ZN(n958) );
  XNOR2_X1 U883 ( .A(n800), .B(n958), .ZN(n801) );
  NOR2_X1 U884 ( .A1(G2100), .A2(n801), .ZN(n802) );
  XNOR2_X1 U885 ( .A(KEYINPUT83), .B(n802), .ZN(G156) );
  NAND2_X1 U886 ( .A1(G559), .A2(n907), .ZN(n803) );
  XNOR2_X1 U887 ( .A(n803), .B(n939), .ZN(n822) );
  NOR2_X1 U888 ( .A1(G860), .A2(n822), .ZN(n813) );
  NAND2_X1 U889 ( .A1(n804), .A2(G67), .ZN(n806) );
  NAND2_X1 U890 ( .A1(G55), .A2(n582), .ZN(n805) );
  NAND2_X1 U891 ( .A1(n806), .A2(n805), .ZN(n812) );
  NAND2_X1 U892 ( .A1(G93), .A2(n807), .ZN(n810) );
  NAND2_X1 U893 ( .A1(G80), .A2(n808), .ZN(n809) );
  NAND2_X1 U894 ( .A1(n810), .A2(n809), .ZN(n811) );
  NOR2_X1 U895 ( .A1(n812), .A2(n811), .ZN(n819) );
  XNOR2_X1 U896 ( .A(n813), .B(n819), .ZN(G145) );
  NOR2_X1 U897 ( .A1(G868), .A2(n819), .ZN(n814) );
  XNOR2_X1 U898 ( .A(n814), .B(KEYINPUT91), .ZN(n825) );
  XOR2_X1 U899 ( .A(KEYINPUT19), .B(KEYINPUT90), .Z(n815) );
  XNOR2_X1 U900 ( .A(G299), .B(n815), .ZN(n816) );
  XNOR2_X1 U901 ( .A(n816), .B(G290), .ZN(n817) );
  XNOR2_X1 U902 ( .A(n817), .B(G288), .ZN(n818) );
  XNOR2_X1 U903 ( .A(n819), .B(n818), .ZN(n820) );
  XNOR2_X1 U904 ( .A(n820), .B(G305), .ZN(n821) );
  XNOR2_X1 U905 ( .A(G166), .B(n821), .ZN(n910) );
  XNOR2_X1 U906 ( .A(n910), .B(n822), .ZN(n823) );
  NAND2_X1 U907 ( .A1(G868), .A2(n823), .ZN(n824) );
  NAND2_X1 U908 ( .A1(n825), .A2(n824), .ZN(G295) );
  NAND2_X1 U909 ( .A1(G2078), .A2(G2084), .ZN(n826) );
  XOR2_X1 U910 ( .A(KEYINPUT20), .B(n826), .Z(n827) );
  NAND2_X1 U911 ( .A1(G2090), .A2(n827), .ZN(n828) );
  XNOR2_X1 U912 ( .A(KEYINPUT21), .B(n828), .ZN(n829) );
  NAND2_X1 U913 ( .A1(n829), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U914 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U915 ( .A(KEYINPUT72), .B(G82), .Z(G220) );
  NAND2_X1 U916 ( .A1(G483), .A2(G661), .ZN(n837) );
  NOR2_X1 U917 ( .A1(G220), .A2(G219), .ZN(n830) );
  XOR2_X1 U918 ( .A(KEYINPUT22), .B(n830), .Z(n831) );
  NOR2_X1 U919 ( .A1(G218), .A2(n831), .ZN(n832) );
  NAND2_X1 U920 ( .A1(G96), .A2(n832), .ZN(n845) );
  NAND2_X1 U921 ( .A1(n845), .A2(G2106), .ZN(n836) );
  NAND2_X1 U922 ( .A1(G120), .A2(G69), .ZN(n833) );
  NOR2_X1 U923 ( .A1(G237), .A2(n833), .ZN(n834) );
  NAND2_X1 U924 ( .A1(G108), .A2(n834), .ZN(n846) );
  NAND2_X1 U925 ( .A1(n846), .A2(G567), .ZN(n835) );
  NAND2_X1 U926 ( .A1(n836), .A2(n835), .ZN(n847) );
  NOR2_X1 U927 ( .A1(n837), .A2(n847), .ZN(n838) );
  XNOR2_X1 U928 ( .A(n838), .B(KEYINPUT92), .ZN(n844) );
  NAND2_X1 U929 ( .A1(G36), .A2(n844), .ZN(G176) );
  NAND2_X1 U930 ( .A1(G2106), .A2(n839), .ZN(G217) );
  NAND2_X1 U931 ( .A1(G15), .A2(G2), .ZN(n841) );
  INV_X1 U932 ( .A(G661), .ZN(n840) );
  NOR2_X1 U933 ( .A1(n841), .A2(n840), .ZN(n842) );
  XNOR2_X1 U934 ( .A(n842), .B(KEYINPUT111), .ZN(G259) );
  NAND2_X1 U935 ( .A1(G3), .A2(G1), .ZN(n843) );
  NAND2_X1 U936 ( .A1(n844), .A2(n843), .ZN(G188) );
  XOR2_X1 U937 ( .A(G69), .B(KEYINPUT112), .Z(G235) );
  INV_X1 U939 ( .A(G120), .ZN(G236) );
  INV_X1 U940 ( .A(G96), .ZN(G221) );
  NOR2_X1 U941 ( .A1(n846), .A2(n845), .ZN(G325) );
  INV_X1 U942 ( .A(G325), .ZN(G261) );
  INV_X1 U943 ( .A(n847), .ZN(G319) );
  XOR2_X1 U944 ( .A(G2100), .B(G2096), .Z(n849) );
  XNOR2_X1 U945 ( .A(KEYINPUT42), .B(G2678), .ZN(n848) );
  XNOR2_X1 U946 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U947 ( .A(KEYINPUT43), .B(G2072), .Z(n851) );
  XNOR2_X1 U948 ( .A(G2067), .B(G2090), .ZN(n850) );
  XNOR2_X1 U949 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U950 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U951 ( .A(G2078), .B(G2084), .ZN(n854) );
  XNOR2_X1 U952 ( .A(n855), .B(n854), .ZN(G227) );
  XOR2_X1 U953 ( .A(G2474), .B(G1986), .Z(n857) );
  XNOR2_X1 U954 ( .A(G1996), .B(G1991), .ZN(n856) );
  XNOR2_X1 U955 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U956 ( .A(n858), .B(KEYINPUT113), .Z(n860) );
  XNOR2_X1 U957 ( .A(G1966), .B(G1981), .ZN(n859) );
  XNOR2_X1 U958 ( .A(n860), .B(n859), .ZN(n864) );
  XOR2_X1 U959 ( .A(G1976), .B(G1956), .Z(n862) );
  XNOR2_X1 U960 ( .A(G1971), .B(G1961), .ZN(n861) );
  XNOR2_X1 U961 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U962 ( .A(n864), .B(n863), .Z(n866) );
  XNOR2_X1 U963 ( .A(KEYINPUT41), .B(KEYINPUT114), .ZN(n865) );
  XNOR2_X1 U964 ( .A(n866), .B(n865), .ZN(G229) );
  NAND2_X1 U965 ( .A1(G100), .A2(n894), .ZN(n868) );
  NAND2_X1 U966 ( .A1(G136), .A2(n895), .ZN(n867) );
  NAND2_X1 U967 ( .A1(n868), .A2(n867), .ZN(n873) );
  NAND2_X1 U968 ( .A1(n890), .A2(G124), .ZN(n869) );
  XNOR2_X1 U969 ( .A(n869), .B(KEYINPUT44), .ZN(n871) );
  NAND2_X1 U970 ( .A1(G112), .A2(n891), .ZN(n870) );
  NAND2_X1 U971 ( .A1(n871), .A2(n870), .ZN(n872) );
  NOR2_X1 U972 ( .A1(n873), .A2(n872), .ZN(G162) );
  NAND2_X1 U973 ( .A1(G103), .A2(n894), .ZN(n875) );
  NAND2_X1 U974 ( .A1(G139), .A2(n895), .ZN(n874) );
  NAND2_X1 U975 ( .A1(n875), .A2(n874), .ZN(n880) );
  NAND2_X1 U976 ( .A1(G127), .A2(n890), .ZN(n877) );
  NAND2_X1 U977 ( .A1(G115), .A2(n891), .ZN(n876) );
  NAND2_X1 U978 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U979 ( .A(KEYINPUT47), .B(n878), .Z(n879) );
  NOR2_X1 U980 ( .A1(n880), .A2(n879), .ZN(n970) );
  XNOR2_X1 U981 ( .A(n970), .B(n881), .ZN(n882) );
  XNOR2_X1 U982 ( .A(n882), .B(n958), .ZN(n886) );
  XOR2_X1 U983 ( .A(KEYINPUT48), .B(KEYINPUT115), .Z(n884) );
  XNOR2_X1 U984 ( .A(G164), .B(KEYINPUT46), .ZN(n883) );
  XNOR2_X1 U985 ( .A(n884), .B(n883), .ZN(n885) );
  XOR2_X1 U986 ( .A(n886), .B(n885), .Z(n889) );
  XNOR2_X1 U987 ( .A(G160), .B(n887), .ZN(n888) );
  XNOR2_X1 U988 ( .A(n889), .B(n888), .ZN(n905) );
  NAND2_X1 U989 ( .A1(G130), .A2(n890), .ZN(n893) );
  NAND2_X1 U990 ( .A1(G118), .A2(n891), .ZN(n892) );
  NAND2_X1 U991 ( .A1(n893), .A2(n892), .ZN(n900) );
  NAND2_X1 U992 ( .A1(G106), .A2(n894), .ZN(n897) );
  NAND2_X1 U993 ( .A1(G142), .A2(n895), .ZN(n896) );
  NAND2_X1 U994 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U995 ( .A(n898), .B(KEYINPUT45), .Z(n899) );
  NOR2_X1 U996 ( .A1(n900), .A2(n899), .ZN(n902) );
  XNOR2_X1 U997 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U998 ( .A(G162), .B(n903), .Z(n904) );
  XNOR2_X1 U999 ( .A(n905), .B(n904), .ZN(n906) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n906), .ZN(G395) );
  XOR2_X1 U1001 ( .A(n907), .B(n939), .Z(n909) );
  XNOR2_X1 U1002 ( .A(G286), .B(G171), .ZN(n908) );
  XNOR2_X1 U1003 ( .A(n909), .B(n908), .ZN(n911) );
  XNOR2_X1 U1004 ( .A(n911), .B(n910), .ZN(n912) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n912), .ZN(G397) );
  XOR2_X1 U1006 ( .A(G2451), .B(G2430), .Z(n914) );
  XNOR2_X1 U1007 ( .A(G2438), .B(G2443), .ZN(n913) );
  XNOR2_X1 U1008 ( .A(n914), .B(n913), .ZN(n920) );
  XOR2_X1 U1009 ( .A(G2435), .B(G2454), .Z(n916) );
  XNOR2_X1 U1010 ( .A(G1341), .B(G1348), .ZN(n915) );
  XNOR2_X1 U1011 ( .A(n916), .B(n915), .ZN(n918) );
  XOR2_X1 U1012 ( .A(G2446), .B(G2427), .Z(n917) );
  XNOR2_X1 U1013 ( .A(n918), .B(n917), .ZN(n919) );
  XOR2_X1 U1014 ( .A(n920), .B(n919), .Z(n921) );
  NAND2_X1 U1015 ( .A1(G14), .A2(n921), .ZN(n927) );
  NAND2_X1 U1016 ( .A1(G319), .A2(n927), .ZN(n924) );
  NOR2_X1 U1017 ( .A1(G227), .A2(G229), .ZN(n922) );
  XNOR2_X1 U1018 ( .A(KEYINPUT49), .B(n922), .ZN(n923) );
  NOR2_X1 U1019 ( .A1(n924), .A2(n923), .ZN(n926) );
  NOR2_X1 U1020 ( .A1(G395), .A2(G397), .ZN(n925) );
  NAND2_X1 U1021 ( .A1(n926), .A2(n925), .ZN(G225) );
  INV_X1 U1022 ( .A(G225), .ZN(G308) );
  INV_X1 U1023 ( .A(G108), .ZN(G238) );
  INV_X1 U1024 ( .A(n927), .ZN(G401) );
  XNOR2_X1 U1025 ( .A(G16), .B(KEYINPUT56), .ZN(n951) );
  XNOR2_X1 U1026 ( .A(G301), .B(G1961), .ZN(n930) );
  XNOR2_X1 U1027 ( .A(n928), .B(G1348), .ZN(n929) );
  NOR2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n934) );
  XNOR2_X1 U1029 ( .A(G1956), .B(G299), .ZN(n931) );
  NOR2_X1 U1030 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n936) );
  XNOR2_X1 U1032 ( .A(G1971), .B(G303), .ZN(n935) );
  NOR2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(n938) );
  NAND2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(n947) );
  XOR2_X1 U1035 ( .A(n939), .B(G1341), .Z(n945) );
  XOR2_X1 U1036 ( .A(G1966), .B(G168), .Z(n940) );
  NOR2_X1 U1037 ( .A1(n941), .A2(n940), .ZN(n942) );
  XOR2_X1 U1038 ( .A(KEYINPUT122), .B(n942), .Z(n943) );
  XNOR2_X1 U1039 ( .A(KEYINPUT57), .B(n943), .ZN(n944) );
  NAND2_X1 U1040 ( .A1(n945), .A2(n944), .ZN(n946) );
  NOR2_X1 U1041 ( .A1(n947), .A2(n946), .ZN(n949) );
  NAND2_X1 U1042 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1043 ( .A1(n951), .A2(n950), .ZN(n1034) );
  INV_X1 U1044 ( .A(KEYINPUT55), .ZN(n980) );
  XNOR2_X1 U1045 ( .A(KEYINPUT52), .B(KEYINPUT119), .ZN(n978) );
  XOR2_X1 U1046 ( .A(G2090), .B(G162), .Z(n952) );
  NOR2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n954) );
  XOR2_X1 U1048 ( .A(KEYINPUT51), .B(n954), .Z(n968) );
  INV_X1 U1049 ( .A(n955), .ZN(n957) );
  NOR2_X1 U1050 ( .A1(n957), .A2(n956), .ZN(n964) );
  XNOR2_X1 U1051 ( .A(G160), .B(G2084), .ZN(n959) );
  NAND2_X1 U1052 ( .A1(n959), .A2(n958), .ZN(n960) );
  NOR2_X1 U1053 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1054 ( .A(n962), .B(KEYINPUT116), .ZN(n963) );
  NAND2_X1 U1055 ( .A1(n964), .A2(n963), .ZN(n965) );
  NOR2_X1 U1056 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1057 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1058 ( .A(KEYINPUT117), .B(n969), .ZN(n976) );
  XOR2_X1 U1059 ( .A(G2072), .B(n970), .Z(n972) );
  XOR2_X1 U1060 ( .A(G164), .B(G2078), .Z(n971) );
  NOR2_X1 U1061 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1062 ( .A(n973), .B(KEYINPUT50), .ZN(n974) );
  XNOR2_X1 U1063 ( .A(n974), .B(KEYINPUT118), .ZN(n975) );
  NAND2_X1 U1064 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1065 ( .A(n978), .B(n977), .ZN(n979) );
  NAND2_X1 U1066 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1067 ( .A1(n981), .A2(G29), .ZN(n1005) );
  XOR2_X1 U1068 ( .A(G2090), .B(G35), .Z(n984) );
  XOR2_X1 U1069 ( .A(KEYINPUT54), .B(G34), .Z(n982) );
  XNOR2_X1 U1070 ( .A(n982), .B(G2084), .ZN(n983) );
  NAND2_X1 U1071 ( .A1(n984), .A2(n983), .ZN(n998) );
  XOR2_X1 U1072 ( .A(G1991), .B(G25), .Z(n985) );
  NAND2_X1 U1073 ( .A1(n985), .A2(G28), .ZN(n994) );
  XNOR2_X1 U1074 ( .A(G1996), .B(G32), .ZN(n987) );
  XNOR2_X1 U1075 ( .A(G33), .B(G2072), .ZN(n986) );
  NOR2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n992) );
  XNOR2_X1 U1077 ( .A(G2067), .B(G26), .ZN(n990) );
  XNOR2_X1 U1078 ( .A(G27), .B(n988), .ZN(n989) );
  NOR2_X1 U1079 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1080 ( .A1(n992), .A2(n991), .ZN(n993) );
  NOR2_X1 U1081 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1082 ( .A(KEYINPUT120), .B(n995), .ZN(n996) );
  XNOR2_X1 U1083 ( .A(KEYINPUT53), .B(n996), .ZN(n997) );
  NOR2_X1 U1084 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1085 ( .A(KEYINPUT55), .B(n999), .ZN(n1001) );
  INV_X1 U1086 ( .A(G29), .ZN(n1000) );
  NAND2_X1 U1087 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1088 ( .A1(n1002), .A2(G11), .ZN(n1003) );
  XNOR2_X1 U1089 ( .A(KEYINPUT121), .B(n1003), .ZN(n1004) );
  NAND2_X1 U1090 ( .A1(n1005), .A2(n1004), .ZN(n1032) );
  XNOR2_X1 U1091 ( .A(G1348), .B(KEYINPUT59), .ZN(n1006) );
  XNOR2_X1 U1092 ( .A(n1006), .B(G4), .ZN(n1010) );
  XNOR2_X1 U1093 ( .A(G1341), .B(G19), .ZN(n1008) );
  XNOR2_X1 U1094 ( .A(G1981), .B(G6), .ZN(n1007) );
  NOR2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1096 ( .A1(n1010), .A2(n1009), .ZN(n1013) );
  XOR2_X1 U1097 ( .A(KEYINPUT123), .B(G1956), .Z(n1011) );
  XNOR2_X1 U1098 ( .A(G20), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1099 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1100 ( .A(KEYINPUT60), .B(n1014), .ZN(n1018) );
  XNOR2_X1 U1101 ( .A(G1961), .B(G5), .ZN(n1016) );
  XNOR2_X1 U1102 ( .A(G1966), .B(G21), .ZN(n1015) );
  NOR2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1026) );
  XNOR2_X1 U1105 ( .A(G1986), .B(G24), .ZN(n1020) );
  XNOR2_X1 U1106 ( .A(G23), .B(G1976), .ZN(n1019) );
  NOR2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1023) );
  XOR2_X1 U1108 ( .A(G1971), .B(KEYINPUT124), .Z(n1021) );
  XNOR2_X1 U1109 ( .A(G22), .B(n1021), .ZN(n1022) );
  NAND2_X1 U1110 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1111 ( .A(KEYINPUT58), .B(n1024), .ZN(n1025) );
  NOR2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1113 ( .A(n1027), .B(KEYINPUT61), .ZN(n1028) );
  XNOR2_X1 U1114 ( .A(KEYINPUT125), .B(n1028), .ZN(n1029) );
  NOR2_X1 U1115 ( .A1(G16), .A2(n1029), .ZN(n1030) );
  XNOR2_X1 U1116 ( .A(n1030), .B(KEYINPUT126), .ZN(n1031) );
  NOR2_X1 U1117 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NAND2_X1 U1118 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XOR2_X1 U1119 ( .A(KEYINPUT62), .B(n1035), .Z(G311) );
  INV_X1 U1120 ( .A(G311), .ZN(G150) );
endmodule

